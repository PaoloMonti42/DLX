
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_dlx is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
subtype bus32 is std_logic_vector (31 downto 0);
type aluOp is (NOP, ADDOP, SUBOP, MULOP, ANDOP, OROP, XOROP, SLLOP, SRLOP, 
   SRAOP, GTOP, GETOP, LTOP, LETOP, EQOP, NEQOP, GTUOP, GETUOP, LTUOP, LETUOP, 
   LHIOP);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_dlx;

package body CONV_PACK_dlx is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return ADDOP;
         when "00010" => return SUBOP;
         when "00011" => return MULOP;
         when "00100" => return ANDOP;
         when "00101" => return OROP;
         when "00110" => return XOROP;
         when "00111" => return SLLOP;
         when "01000" => return SRLOP;
         when "01001" => return SRAOP;
         when "01010" => return GTOP;
         when "01011" => return GETOP;
         when "01100" => return LTOP;
         when "01101" => return LETOP;
         when "01110" => return EQOP;
         when "01111" => return NEQOP;
         when "10000" => return GTUOP;
         when "10001" => return GETUOP;
         when "10010" => return LTUOP;
         when "10011" => return LETUOP;
         when "10100" => return LHIOP;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when ADDOP => return "00001";
         when SUBOP => return "00010";
         when MULOP => return "00011";
         when ANDOP => return "00100";
         when OROP => return "00101";
         when XOROP => return "00110";
         when SLLOP => return "00111";
         when SRLOP => return "01000";
         when SRAOP => return "01001";
         when GTOP => return "01010";
         when GETOP => return "01011";
         when LTOP => return "01100";
         when LETOP => return "01101";
         when EQOP => return "01110";
         when NEQOP => return "01111";
         when GTUOP => return "10000";
         when GETUOP => return "10001";
         when LTUOP => return "10010";
         when LETUOP => return "10011";
         when LHIOP => return "10100";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_dlx;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_217 is

   port( A : in std_logic;  Y : out std_logic);

end IV_217;

architecture SYN_BEHAVIORAL of IV_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_216 is

   port( A : in std_logic;  Y : out std_logic);

end IV_216;

architecture SYN_BEHAVIORAL of IV_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_215 is

   port( A : in std_logic;  Y : out std_logic);

end IV_215;

architecture SYN_BEHAVIORAL of IV_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_214 is

   port( A : in std_logic;  Y : out std_logic);

end IV_214;

architecture SYN_BEHAVIORAL of IV_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_213 is

   port( A : in std_logic;  Y : out std_logic);

end IV_213;

architecture SYN_BEHAVIORAL of IV_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_212 is

   port( A : in std_logic;  Y : out std_logic);

end IV_212;

architecture SYN_BEHAVIORAL of IV_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_211 is

   port( A : in std_logic;  Y : out std_logic);

end IV_211;

architecture SYN_BEHAVIORAL of IV_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_210 is

   port( A : in std_logic;  Y : out std_logic);

end IV_210;

architecture SYN_BEHAVIORAL of IV_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_209 is

   port( A : in std_logic;  Y : out std_logic);

end IV_209;

architecture SYN_BEHAVIORAL of IV_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_208 is

   port( A : in std_logic;  Y : out std_logic);

end IV_208;

architecture SYN_BEHAVIORAL of IV_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_207 is

   port( A : in std_logic;  Y : out std_logic);

end IV_207;

architecture SYN_BEHAVIORAL of IV_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_206 is

   port( A : in std_logic;  Y : out std_logic);

end IV_206;

architecture SYN_BEHAVIORAL of IV_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_205 is

   port( A : in std_logic;  Y : out std_logic);

end IV_205;

architecture SYN_BEHAVIORAL of IV_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_204 is

   port( A : in std_logic;  Y : out std_logic);

end IV_204;

architecture SYN_BEHAVIORAL of IV_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_203 is

   port( A : in std_logic;  Y : out std_logic);

end IV_203;

architecture SYN_BEHAVIORAL of IV_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_202 is

   port( A : in std_logic;  Y : out std_logic);

end IV_202;

architecture SYN_BEHAVIORAL of IV_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_201 is

   port( A : in std_logic;  Y : out std_logic);

end IV_201;

architecture SYN_BEHAVIORAL of IV_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_200 is

   port( A : in std_logic;  Y : out std_logic);

end IV_200;

architecture SYN_BEHAVIORAL of IV_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_199 is

   port( A : in std_logic;  Y : out std_logic);

end IV_199;

architecture SYN_BEHAVIORAL of IV_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_198 is

   port( A : in std_logic;  Y : out std_logic);

end IV_198;

architecture SYN_BEHAVIORAL of IV_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_197 is

   port( A : in std_logic;  Y : out std_logic);

end IV_197;

architecture SYN_BEHAVIORAL of IV_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_196 is

   port( A : in std_logic;  Y : out std_logic);

end IV_196;

architecture SYN_BEHAVIORAL of IV_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_195 is

   port( A : in std_logic;  Y : out std_logic);

end IV_195;

architecture SYN_BEHAVIORAL of IV_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_194 is

   port( A : in std_logic;  Y : out std_logic);

end IV_194;

architecture SYN_BEHAVIORAL of IV_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_193 is

   port( A : in std_logic;  Y : out std_logic);

end IV_193;

architecture SYN_BEHAVIORAL of IV_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_192 is

   port( A : in std_logic;  Y : out std_logic);

end IV_192;

architecture SYN_BEHAVIORAL of IV_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_191 is

   port( A : in std_logic;  Y : out std_logic);

end IV_191;

architecture SYN_BEHAVIORAL of IV_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_190 is

   port( A : in std_logic;  Y : out std_logic);

end IV_190;

architecture SYN_BEHAVIORAL of IV_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_189 is

   port( A : in std_logic;  Y : out std_logic);

end IV_189;

architecture SYN_BEHAVIORAL of IV_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_188 is

   port( A : in std_logic;  Y : out std_logic);

end IV_188;

architecture SYN_BEHAVIORAL of IV_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_187 is

   port( A : in std_logic;  Y : out std_logic);

end IV_187;

architecture SYN_BEHAVIORAL of IV_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_186 is

   port( A : in std_logic;  Y : out std_logic);

end IV_186;

architecture SYN_BEHAVIORAL of IV_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_185 is

   port( A : in std_logic;  Y : out std_logic);

end IV_185;

architecture SYN_BEHAVIORAL of IV_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_184 is

   port( A : in std_logic;  Y : out std_logic);

end IV_184;

architecture SYN_BEHAVIORAL of IV_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_183 is

   port( A : in std_logic;  Y : out std_logic);

end IV_183;

architecture SYN_BEHAVIORAL of IV_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_182 is

   port( A : in std_logic;  Y : out std_logic);

end IV_182;

architecture SYN_BEHAVIORAL of IV_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_181 is

   port( A : in std_logic;  Y : out std_logic);

end IV_181;

architecture SYN_BEHAVIORAL of IV_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_180 is

   port( A : in std_logic;  Y : out std_logic);

end IV_180;

architecture SYN_BEHAVIORAL of IV_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_179 is

   port( A : in std_logic;  Y : out std_logic);

end IV_179;

architecture SYN_BEHAVIORAL of IV_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_178 is

   port( A : in std_logic;  Y : out std_logic);

end IV_178;

architecture SYN_BEHAVIORAL of IV_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_177 is

   port( A : in std_logic;  Y : out std_logic);

end IV_177;

architecture SYN_BEHAVIORAL of IV_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_176 is

   port( A : in std_logic;  Y : out std_logic);

end IV_176;

architecture SYN_BEHAVIORAL of IV_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_175 is

   port( A : in std_logic;  Y : out std_logic);

end IV_175;

architecture SYN_BEHAVIORAL of IV_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_174 is

   port( A : in std_logic;  Y : out std_logic);

end IV_174;

architecture SYN_BEHAVIORAL of IV_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_173 is

   port( A : in std_logic;  Y : out std_logic);

end IV_173;

architecture SYN_BEHAVIORAL of IV_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_172 is

   port( A : in std_logic;  Y : out std_logic);

end IV_172;

architecture SYN_BEHAVIORAL of IV_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_171 is

   port( A : in std_logic;  Y : out std_logic);

end IV_171;

architecture SYN_BEHAVIORAL of IV_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_170 is

   port( A : in std_logic;  Y : out std_logic);

end IV_170;

architecture SYN_BEHAVIORAL of IV_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_169 is

   port( A : in std_logic;  Y : out std_logic);

end IV_169;

architecture SYN_BEHAVIORAL of IV_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_168 is

   port( A : in std_logic;  Y : out std_logic);

end IV_168;

architecture SYN_BEHAVIORAL of IV_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_167 is

   port( A : in std_logic;  Y : out std_logic);

end IV_167;

architecture SYN_BEHAVIORAL of IV_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_166 is

   port( A : in std_logic;  Y : out std_logic);

end IV_166;

architecture SYN_BEHAVIORAL of IV_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_165 is

   port( A : in std_logic;  Y : out std_logic);

end IV_165;

architecture SYN_BEHAVIORAL of IV_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_164 is

   port( A : in std_logic;  Y : out std_logic);

end IV_164;

architecture SYN_BEHAVIORAL of IV_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_163 is

   port( A : in std_logic;  Y : out std_logic);

end IV_163;

architecture SYN_BEHAVIORAL of IV_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_162 is

   port( A : in std_logic;  Y : out std_logic);

end IV_162;

architecture SYN_BEHAVIORAL of IV_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_161 is

   port( A : in std_logic;  Y : out std_logic);

end IV_161;

architecture SYN_BEHAVIORAL of IV_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_160 is

   port( A : in std_logic;  Y : out std_logic);

end IV_160;

architecture SYN_BEHAVIORAL of IV_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_159 is

   port( A : in std_logic;  Y : out std_logic);

end IV_159;

architecture SYN_BEHAVIORAL of IV_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_158 is

   port( A : in std_logic;  Y : out std_logic);

end IV_158;

architecture SYN_BEHAVIORAL of IV_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_157 is

   port( A : in std_logic;  Y : out std_logic);

end IV_157;

architecture SYN_BEHAVIORAL of IV_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_156 is

   port( A : in std_logic;  Y : out std_logic);

end IV_156;

architecture SYN_BEHAVIORAL of IV_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_155 is

   port( A : in std_logic;  Y : out std_logic);

end IV_155;

architecture SYN_BEHAVIORAL of IV_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_154 is

   port( A : in std_logic;  Y : out std_logic);

end IV_154;

architecture SYN_BEHAVIORAL of IV_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_153 is

   port( A : in std_logic;  Y : out std_logic);

end IV_153;

architecture SYN_BEHAVIORAL of IV_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_152 is

   port( A : in std_logic;  Y : out std_logic);

end IV_152;

architecture SYN_BEHAVIORAL of IV_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_151 is

   port( A : in std_logic;  Y : out std_logic);

end IV_151;

architecture SYN_BEHAVIORAL of IV_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_150 is

   port( A : in std_logic;  Y : out std_logic);

end IV_150;

architecture SYN_BEHAVIORAL of IV_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_149 is

   port( A : in std_logic;  Y : out std_logic);

end IV_149;

architecture SYN_BEHAVIORAL of IV_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_148 is

   port( A : in std_logic;  Y : out std_logic);

end IV_148;

architecture SYN_BEHAVIORAL of IV_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_147 is

   port( A : in std_logic;  Y : out std_logic);

end IV_147;

architecture SYN_BEHAVIORAL of IV_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_146 is

   port( A : in std_logic;  Y : out std_logic);

end IV_146;

architecture SYN_BEHAVIORAL of IV_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_145 is

   port( A : in std_logic;  Y : out std_logic);

end IV_145;

architecture SYN_BEHAVIORAL of IV_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_144 is

   port( A : in std_logic;  Y : out std_logic);

end IV_144;

architecture SYN_BEHAVIORAL of IV_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_143 is

   port( A : in std_logic;  Y : out std_logic);

end IV_143;

architecture SYN_BEHAVIORAL of IV_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_142 is

   port( A : in std_logic;  Y : out std_logic);

end IV_142;

architecture SYN_BEHAVIORAL of IV_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_141 is

   port( A : in std_logic;  Y : out std_logic);

end IV_141;

architecture SYN_BEHAVIORAL of IV_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_140 is

   port( A : in std_logic;  Y : out std_logic);

end IV_140;

architecture SYN_BEHAVIORAL of IV_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_139 is

   port( A : in std_logic;  Y : out std_logic);

end IV_139;

architecture SYN_BEHAVIORAL of IV_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_138 is

   port( A : in std_logic;  Y : out std_logic);

end IV_138;

architecture SYN_BEHAVIORAL of IV_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_137 is

   port( A : in std_logic;  Y : out std_logic);

end IV_137;

architecture SYN_BEHAVIORAL of IV_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_136 is

   port( A : in std_logic;  Y : out std_logic);

end IV_136;

architecture SYN_BEHAVIORAL of IV_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_135 is

   port( A : in std_logic;  Y : out std_logic);

end IV_135;

architecture SYN_BEHAVIORAL of IV_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_134 is

   port( A : in std_logic;  Y : out std_logic);

end IV_134;

architecture SYN_BEHAVIORAL of IV_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_133 is

   port( A : in std_logic;  Y : out std_logic);

end IV_133;

architecture SYN_BEHAVIORAL of IV_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_132 is

   port( A : in std_logic;  Y : out std_logic);

end IV_132;

architecture SYN_BEHAVIORAL of IV_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_131 is

   port( A : in std_logic;  Y : out std_logic);

end IV_131;

architecture SYN_BEHAVIORAL of IV_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_130 is

   port( A : in std_logic;  Y : out std_logic);

end IV_130;

architecture SYN_BEHAVIORAL of IV_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_129 is

   port( A : in std_logic;  Y : out std_logic);

end IV_129;

architecture SYN_BEHAVIORAL of IV_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_128 is

   port( A : in std_logic;  Y : out std_logic);

end IV_128;

architecture SYN_BEHAVIORAL of IV_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_665 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_665;

architecture SYN_ARCH1 of ND2_665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_664 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_664;

architecture SYN_ARCH1 of ND2_664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_663 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_663;

architecture SYN_ARCH1 of ND2_663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_662 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_662;

architecture SYN_ARCH1 of ND2_662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_661 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_661;

architecture SYN_ARCH1 of ND2_661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_660 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_660;

architecture SYN_ARCH1 of ND2_660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_659 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_659;

architecture SYN_ARCH1 of ND2_659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_658 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_658;

architecture SYN_ARCH1 of ND2_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_657 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_657;

architecture SYN_ARCH1 of ND2_657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_656 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_656;

architecture SYN_ARCH1 of ND2_656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_655 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_655;

architecture SYN_ARCH1 of ND2_655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_654 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_654;

architecture SYN_ARCH1 of ND2_654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_653 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_653;

architecture SYN_ARCH1 of ND2_653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_652 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_652;

architecture SYN_ARCH1 of ND2_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_651 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_651;

architecture SYN_ARCH1 of ND2_651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_650 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_650;

architecture SYN_ARCH1 of ND2_650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_649 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_649;

architecture SYN_ARCH1 of ND2_649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_648 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_648;

architecture SYN_ARCH1 of ND2_648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_647 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_647;

architecture SYN_ARCH1 of ND2_647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_646 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_646;

architecture SYN_ARCH1 of ND2_646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_645 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_645;

architecture SYN_ARCH1 of ND2_645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_644 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_644;

architecture SYN_ARCH1 of ND2_644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_643 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_643;

architecture SYN_ARCH1 of ND2_643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_642 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_642;

architecture SYN_ARCH1 of ND2_642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_641 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_641;

architecture SYN_ARCH1 of ND2_641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_640 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_640;

architecture SYN_ARCH1 of ND2_640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_639 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_639;

architecture SYN_ARCH1 of ND2_639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_638 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_638;

architecture SYN_ARCH1 of ND2_638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_637 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_637;

architecture SYN_ARCH1 of ND2_637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_636 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_636;

architecture SYN_ARCH1 of ND2_636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_635 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_635;

architecture SYN_ARCH1 of ND2_635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_634 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_634;

architecture SYN_ARCH1 of ND2_634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_633 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_633;

architecture SYN_ARCH1 of ND2_633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_632 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_632;

architecture SYN_ARCH1 of ND2_632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_631 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_631;

architecture SYN_ARCH1 of ND2_631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_630 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_630;

architecture SYN_ARCH1 of ND2_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_629 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_629;

architecture SYN_ARCH1 of ND2_629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_628 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_628;

architecture SYN_ARCH1 of ND2_628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_627 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_627;

architecture SYN_ARCH1 of ND2_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_626 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_626;

architecture SYN_ARCH1 of ND2_626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_625 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_625;

architecture SYN_ARCH1 of ND2_625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_624 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_624;

architecture SYN_ARCH1 of ND2_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_623 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_623;

architecture SYN_ARCH1 of ND2_623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_622 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_622;

architecture SYN_ARCH1 of ND2_622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_621 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_621;

architecture SYN_ARCH1 of ND2_621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_620 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_620;

architecture SYN_ARCH1 of ND2_620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_619 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_619;

architecture SYN_ARCH1 of ND2_619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_618 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_618;

architecture SYN_ARCH1 of ND2_618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_617 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_617;

architecture SYN_ARCH1 of ND2_617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_616 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_616;

architecture SYN_ARCH1 of ND2_616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_615 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_615;

architecture SYN_ARCH1 of ND2_615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_614 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_614;

architecture SYN_ARCH1 of ND2_614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_613 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_613;

architecture SYN_ARCH1 of ND2_613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_612 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_612;

architecture SYN_ARCH1 of ND2_612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_611 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_611;

architecture SYN_ARCH1 of ND2_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_610 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_610;

architecture SYN_ARCH1 of ND2_610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_609 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_609;

architecture SYN_ARCH1 of ND2_609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_608 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_608;

architecture SYN_ARCH1 of ND2_608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_607 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_607;

architecture SYN_ARCH1 of ND2_607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_606 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_606;

architecture SYN_ARCH1 of ND2_606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_605 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_605;

architecture SYN_ARCH1 of ND2_605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_604 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_604;

architecture SYN_ARCH1 of ND2_604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_603 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_603;

architecture SYN_ARCH1 of ND2_603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_602 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_602;

architecture SYN_ARCH1 of ND2_602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_601 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_601;

architecture SYN_ARCH1 of ND2_601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_600 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_600;

architecture SYN_ARCH1 of ND2_600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_599 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_599;

architecture SYN_ARCH1 of ND2_599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_598 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_598;

architecture SYN_ARCH1 of ND2_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_597 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_597;

architecture SYN_ARCH1 of ND2_597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_596 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_596;

architecture SYN_ARCH1 of ND2_596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_595 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_595;

architecture SYN_ARCH1 of ND2_595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_594 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_594;

architecture SYN_ARCH1 of ND2_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_593 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_593;

architecture SYN_ARCH1 of ND2_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_592 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_592;

architecture SYN_ARCH1 of ND2_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_591 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_591;

architecture SYN_ARCH1 of ND2_591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_590 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_590;

architecture SYN_ARCH1 of ND2_590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_589 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_589;

architecture SYN_ARCH1 of ND2_589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_588 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_588;

architecture SYN_ARCH1 of ND2_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_587 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_587;

architecture SYN_ARCH1 of ND2_587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_586 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_586;

architecture SYN_ARCH1 of ND2_586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_585 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_585;

architecture SYN_ARCH1 of ND2_585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_584 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_584;

architecture SYN_ARCH1 of ND2_584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_583 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_583;

architecture SYN_ARCH1 of ND2_583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_582 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_582;

architecture SYN_ARCH1 of ND2_582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_581 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_581;

architecture SYN_ARCH1 of ND2_581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_580 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_580;

architecture SYN_ARCH1 of ND2_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_579 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_579;

architecture SYN_ARCH1 of ND2_579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_578 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_578;

architecture SYN_ARCH1 of ND2_578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_577 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_577;

architecture SYN_ARCH1 of ND2_577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_576 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_576;

architecture SYN_ARCH1 of ND2_576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_575 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_575;

architecture SYN_ARCH1 of ND2_575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_574 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_574;

architecture SYN_ARCH1 of ND2_574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_573 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_573;

architecture SYN_ARCH1 of ND2_573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_572 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_572;

architecture SYN_ARCH1 of ND2_572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_571 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_571;

architecture SYN_ARCH1 of ND2_571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_570 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_570;

architecture SYN_ARCH1 of ND2_570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_569 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_569;

architecture SYN_ARCH1 of ND2_569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_568 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_568;

architecture SYN_ARCH1 of ND2_568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_567 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_567;

architecture SYN_ARCH1 of ND2_567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_566 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_566;

architecture SYN_ARCH1 of ND2_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_565 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_565;

architecture SYN_ARCH1 of ND2_565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_564 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_564;

architecture SYN_ARCH1 of ND2_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_563 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_563;

architecture SYN_ARCH1 of ND2_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_562 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_562;

architecture SYN_ARCH1 of ND2_562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_561 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_561;

architecture SYN_ARCH1 of ND2_561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_560 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_560;

architecture SYN_ARCH1 of ND2_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_559 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_559;

architecture SYN_ARCH1 of ND2_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_558 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_558;

architecture SYN_ARCH1 of ND2_558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_557 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_557;

architecture SYN_ARCH1 of ND2_557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_556 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_556;

architecture SYN_ARCH1 of ND2_556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_555 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_555;

architecture SYN_ARCH1 of ND2_555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_554 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_554;

architecture SYN_ARCH1 of ND2_554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_553 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_553;

architecture SYN_ARCH1 of ND2_553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_552 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_552;

architecture SYN_ARCH1 of ND2_552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_551 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_551;

architecture SYN_ARCH1 of ND2_551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_550 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_550;

architecture SYN_ARCH1 of ND2_550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_549 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_549;

architecture SYN_ARCH1 of ND2_549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_548 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_548;

architecture SYN_ARCH1 of ND2_548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_547 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_547;

architecture SYN_ARCH1 of ND2_547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_546 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_546;

architecture SYN_ARCH1 of ND2_546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_545 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_545;

architecture SYN_ARCH1 of ND2_545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_544 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_544;

architecture SYN_ARCH1 of ND2_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_543 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_543;

architecture SYN_ARCH1 of ND2_543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_542 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_542;

architecture SYN_ARCH1 of ND2_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_541 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_541;

architecture SYN_ARCH1 of ND2_541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_540 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_540;

architecture SYN_ARCH1 of ND2_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_539 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_539;

architecture SYN_ARCH1 of ND2_539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_538 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_538;

architecture SYN_ARCH1 of ND2_538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_537 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_537;

architecture SYN_ARCH1 of ND2_537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_536 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_536;

architecture SYN_ARCH1 of ND2_536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_535 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_535;

architecture SYN_ARCH1 of ND2_535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_534 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_534;

architecture SYN_ARCH1 of ND2_534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_533 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_533;

architecture SYN_ARCH1 of ND2_533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_532 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_532;

architecture SYN_ARCH1 of ND2_532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_531 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_531;

architecture SYN_ARCH1 of ND2_531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_530 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_530;

architecture SYN_ARCH1 of ND2_530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_529 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_529;

architecture SYN_ARCH1 of ND2_529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_528 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_528;

architecture SYN_ARCH1 of ND2_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_527 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_527;

architecture SYN_ARCH1 of ND2_527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_526 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_526;

architecture SYN_ARCH1 of ND2_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_525 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_525;

architecture SYN_ARCH1 of ND2_525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_524 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_524;

architecture SYN_ARCH1 of ND2_524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_523 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_523;

architecture SYN_ARCH1 of ND2_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_522 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_522;

architecture SYN_ARCH1 of ND2_522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_521 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_521;

architecture SYN_ARCH1 of ND2_521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_520 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_520;

architecture SYN_ARCH1 of ND2_520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_519 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_519;

architecture SYN_ARCH1 of ND2_519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_518 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_518;

architecture SYN_ARCH1 of ND2_518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_517 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_517;

architecture SYN_ARCH1 of ND2_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_516 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_516;

architecture SYN_ARCH1 of ND2_516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_515 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_515;

architecture SYN_ARCH1 of ND2_515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_514 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_514;

architecture SYN_ARCH1 of ND2_514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_513 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_513;

architecture SYN_ARCH1 of ND2_513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_512 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_512;

architecture SYN_ARCH1 of ND2_512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_511 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_511;

architecture SYN_ARCH1 of ND2_511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_510 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_510;

architecture SYN_ARCH1 of ND2_510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_509 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_509;

architecture SYN_ARCH1 of ND2_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_508 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_508;

architecture SYN_ARCH1 of ND2_508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_507 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_507;

architecture SYN_ARCH1 of ND2_507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_506 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_506;

architecture SYN_ARCH1 of ND2_506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_505 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_505;

architecture SYN_ARCH1 of ND2_505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_504 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_504;

architecture SYN_ARCH1 of ND2_504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_503 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_503;

architecture SYN_ARCH1 of ND2_503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_502 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_502;

architecture SYN_ARCH1 of ND2_502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_501 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_501;

architecture SYN_ARCH1 of ND2_501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_500 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_500;

architecture SYN_ARCH1 of ND2_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_499 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_499;

architecture SYN_ARCH1 of ND2_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_498 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_498;

architecture SYN_ARCH1 of ND2_498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_497 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_497;

architecture SYN_ARCH1 of ND2_497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_496 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_496;

architecture SYN_ARCH1 of ND2_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_495 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_495;

architecture SYN_ARCH1 of ND2_495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_494 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_494;

architecture SYN_ARCH1 of ND2_494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_493 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_493;

architecture SYN_ARCH1 of ND2_493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_492 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_492;

architecture SYN_ARCH1 of ND2_492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_491 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_491;

architecture SYN_ARCH1 of ND2_491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_490 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_490;

architecture SYN_ARCH1 of ND2_490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_489 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_489;

architecture SYN_ARCH1 of ND2_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_488 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_488;

architecture SYN_ARCH1 of ND2_488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_487 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_487;

architecture SYN_ARCH1 of ND2_487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_486 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_486;

architecture SYN_ARCH1 of ND2_486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_485 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_485;

architecture SYN_ARCH1 of ND2_485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_484 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_484;

architecture SYN_ARCH1 of ND2_484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_483 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_483;

architecture SYN_ARCH1 of ND2_483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_482 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_482;

architecture SYN_ARCH1 of ND2_482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_481 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_481;

architecture SYN_ARCH1 of ND2_481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_480 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_480;

architecture SYN_ARCH1 of ND2_480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_479 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_479;

architecture SYN_ARCH1 of ND2_479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_478 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_478;

architecture SYN_ARCH1 of ND2_478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_477 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_477;

architecture SYN_ARCH1 of ND2_477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_476 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_476;

architecture SYN_ARCH1 of ND2_476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_475 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_475;

architecture SYN_ARCH1 of ND2_475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_474 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_474;

architecture SYN_ARCH1 of ND2_474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_473 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_473;

architecture SYN_ARCH1 of ND2_473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_472 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_472;

architecture SYN_ARCH1 of ND2_472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_471 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_471;

architecture SYN_ARCH1 of ND2_471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_470 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_470;

architecture SYN_ARCH1 of ND2_470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_469 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_469;

architecture SYN_ARCH1 of ND2_469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_468 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_468;

architecture SYN_ARCH1 of ND2_468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_467 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_467;

architecture SYN_ARCH1 of ND2_467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_466 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_466;

architecture SYN_ARCH1 of ND2_466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_465 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_465;

architecture SYN_ARCH1 of ND2_465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_464 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_464;

architecture SYN_ARCH1 of ND2_464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_463 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_463;

architecture SYN_ARCH1 of ND2_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_462 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_462;

architecture SYN_ARCH1 of ND2_462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_461 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_461;

architecture SYN_ARCH1 of ND2_461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_460 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_460;

architecture SYN_ARCH1 of ND2_460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_459 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_459;

architecture SYN_ARCH1 of ND2_459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_458 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_458;

architecture SYN_ARCH1 of ND2_458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_457 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_457;

architecture SYN_ARCH1 of ND2_457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_456 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_456;

architecture SYN_ARCH1 of ND2_456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_455 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_455;

architecture SYN_ARCH1 of ND2_455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_454 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_454;

architecture SYN_ARCH1 of ND2_454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_453 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_453;

architecture SYN_ARCH1 of ND2_453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_452 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_452;

architecture SYN_ARCH1 of ND2_452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_451 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_451;

architecture SYN_ARCH1 of ND2_451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_450 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_450;

architecture SYN_ARCH1 of ND2_450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_449 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_449;

architecture SYN_ARCH1 of ND2_449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_448 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_448;

architecture SYN_ARCH1 of ND2_448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_447 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_447;

architecture SYN_ARCH1 of ND2_447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_446 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_446;

architecture SYN_ARCH1 of ND2_446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_445 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_445;

architecture SYN_ARCH1 of ND2_445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_444 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_444;

architecture SYN_ARCH1 of ND2_444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_443 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_443;

architecture SYN_ARCH1 of ND2_443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_442 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_442;

architecture SYN_ARCH1 of ND2_442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_441 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_441;

architecture SYN_ARCH1 of ND2_441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_440 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_440;

architecture SYN_ARCH1 of ND2_440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_439 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_439;

architecture SYN_ARCH1 of ND2_439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_438 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_438;

architecture SYN_ARCH1 of ND2_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_437 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_437;

architecture SYN_ARCH1 of ND2_437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_436 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_436;

architecture SYN_ARCH1 of ND2_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_435 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_435;

architecture SYN_ARCH1 of ND2_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_434 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_434;

architecture SYN_ARCH1 of ND2_434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_433 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_433;

architecture SYN_ARCH1 of ND2_433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_432 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_432;

architecture SYN_ARCH1 of ND2_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_431 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_431;

architecture SYN_ARCH1 of ND2_431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_430 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_430;

architecture SYN_ARCH1 of ND2_430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_429 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_429;

architecture SYN_ARCH1 of ND2_429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_428 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_428;

architecture SYN_ARCH1 of ND2_428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_427 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_427;

architecture SYN_ARCH1 of ND2_427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_426 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_426;

architecture SYN_ARCH1 of ND2_426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_425 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_425;

architecture SYN_ARCH1 of ND2_425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_424 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_424;

architecture SYN_ARCH1 of ND2_424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_423 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_423;

architecture SYN_ARCH1 of ND2_423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_422 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_422;

architecture SYN_ARCH1 of ND2_422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_421 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_421;

architecture SYN_ARCH1 of ND2_421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_420 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_420;

architecture SYN_ARCH1 of ND2_420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_419 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_419;

architecture SYN_ARCH1 of ND2_419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_418 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_418;

architecture SYN_ARCH1 of ND2_418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_417 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_417;

architecture SYN_ARCH1 of ND2_417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_416 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_416;

architecture SYN_ARCH1 of ND2_416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_415 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_415;

architecture SYN_ARCH1 of ND2_415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_414 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_414;

architecture SYN_ARCH1 of ND2_414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_413 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_413;

architecture SYN_ARCH1 of ND2_413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_412 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_412;

architecture SYN_ARCH1 of ND2_412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_411 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_411;

architecture SYN_ARCH1 of ND2_411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_410 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_410;

architecture SYN_ARCH1 of ND2_410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_409 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_409;

architecture SYN_ARCH1 of ND2_409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_408 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_408;

architecture SYN_ARCH1 of ND2_408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_407 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_407;

architecture SYN_ARCH1 of ND2_407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_406 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_406;

architecture SYN_ARCH1 of ND2_406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_405 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_405;

architecture SYN_ARCH1 of ND2_405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_404 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_404;

architecture SYN_ARCH1 of ND2_404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_403 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_403;

architecture SYN_ARCH1 of ND2_403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_402 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_402;

architecture SYN_ARCH1 of ND2_402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_401 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_401;

architecture SYN_ARCH1 of ND2_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_400 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_400;

architecture SYN_ARCH1 of ND2_400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_399 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_399;

architecture SYN_ARCH1 of ND2_399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_398 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_398;

architecture SYN_ARCH1 of ND2_398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_397 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_397;

architecture SYN_ARCH1 of ND2_397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_396 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_396;

architecture SYN_ARCH1 of ND2_396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_395 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_395;

architecture SYN_ARCH1 of ND2_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_394 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_394;

architecture SYN_ARCH1 of ND2_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_393 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_393;

architecture SYN_ARCH1 of ND2_393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_392 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_392;

architecture SYN_ARCH1 of ND2_392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_391 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_391;

architecture SYN_ARCH1 of ND2_391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_390 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_390;

architecture SYN_ARCH1 of ND2_390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_389 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_389;

architecture SYN_ARCH1 of ND2_389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_388 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_388;

architecture SYN_ARCH1 of ND2_388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_387 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_387;

architecture SYN_ARCH1 of ND2_387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_386 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_386;

architecture SYN_ARCH1 of ND2_386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_385 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_385;

architecture SYN_ARCH1 of ND2_385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_384 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_384;

architecture SYN_ARCH1 of ND2_384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_383 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_383;

architecture SYN_ARCH1 of ND2_383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_382 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_382;

architecture SYN_ARCH1 of ND2_382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_381 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_381;

architecture SYN_ARCH1 of ND2_381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_380 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_380;

architecture SYN_ARCH1 of ND2_380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_379 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_379;

architecture SYN_ARCH1 of ND2_379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_378 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_378;

architecture SYN_ARCH1 of ND2_378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_377 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_377;

architecture SYN_ARCH1 of ND2_377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_376 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_376;

architecture SYN_ARCH1 of ND2_376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_375 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_375;

architecture SYN_ARCH1 of ND2_375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_374 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_374;

architecture SYN_ARCH1 of ND2_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_373 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_373;

architecture SYN_ARCH1 of ND2_373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_372 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_372;

architecture SYN_ARCH1 of ND2_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_371 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_371;

architecture SYN_ARCH1 of ND2_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_370 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_370;

architecture SYN_ARCH1 of ND2_370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_369 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_369;

architecture SYN_ARCH1 of ND2_369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_368 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_368;

architecture SYN_ARCH1 of ND2_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_367 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_367;

architecture SYN_ARCH1 of ND2_367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_366 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_366;

architecture SYN_ARCH1 of ND2_366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_365 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_365;

architecture SYN_ARCH1 of ND2_365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_364 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_364;

architecture SYN_ARCH1 of ND2_364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_363 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_363;

architecture SYN_ARCH1 of ND2_363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_362 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_362;

architecture SYN_ARCH1 of ND2_362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_361 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_361;

architecture SYN_ARCH1 of ND2_361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_360 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_360;

architecture SYN_ARCH1 of ND2_360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_359 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_359;

architecture SYN_ARCH1 of ND2_359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_358 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_358;

architecture SYN_ARCH1 of ND2_358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_357 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_357;

architecture SYN_ARCH1 of ND2_357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_356 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_356;

architecture SYN_ARCH1 of ND2_356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_355 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_355;

architecture SYN_ARCH1 of ND2_355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_354 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_354;

architecture SYN_ARCH1 of ND2_354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_353 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_353;

architecture SYN_ARCH1 of ND2_353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_352 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_352;

architecture SYN_ARCH1 of ND2_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_351 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_351;

architecture SYN_ARCH1 of ND2_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_350 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_350;

architecture SYN_ARCH1 of ND2_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_349 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_349;

architecture SYN_ARCH1 of ND2_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_348 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_348;

architecture SYN_ARCH1 of ND2_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_347 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_347;

architecture SYN_ARCH1 of ND2_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_346 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_346;

architecture SYN_ARCH1 of ND2_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_345 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_345;

architecture SYN_ARCH1 of ND2_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_344 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_344;

architecture SYN_ARCH1 of ND2_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_343 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_343;

architecture SYN_ARCH1 of ND2_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_342 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_342;

architecture SYN_ARCH1 of ND2_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_341 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_341;

architecture SYN_ARCH1 of ND2_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_340 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_340;

architecture SYN_ARCH1 of ND2_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_339 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_339;

architecture SYN_ARCH1 of ND2_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_338 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_338;

architecture SYN_ARCH1 of ND2_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_337 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_337;

architecture SYN_ARCH1 of ND2_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_336 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_336;

architecture SYN_ARCH1 of ND2_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_335 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_335;

architecture SYN_ARCH1 of ND2_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_334 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_334;

architecture SYN_ARCH1 of ND2_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_333 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_333;

architecture SYN_ARCH1 of ND2_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_332 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_332;

architecture SYN_ARCH1 of ND2_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_331 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_331;

architecture SYN_ARCH1 of ND2_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_330 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_330;

architecture SYN_ARCH1 of ND2_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_329 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_329;

architecture SYN_ARCH1 of ND2_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_328 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_328;

architecture SYN_ARCH1 of ND2_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_327 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_327;

architecture SYN_ARCH1 of ND2_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_326 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_326;

architecture SYN_ARCH1 of ND2_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_325 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_325;

architecture SYN_ARCH1 of ND2_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_324 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_324;

architecture SYN_ARCH1 of ND2_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_323 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_323;

architecture SYN_ARCH1 of ND2_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_322 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_322;

architecture SYN_ARCH1 of ND2_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_321 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_321;

architecture SYN_ARCH1 of ND2_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_320 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_320;

architecture SYN_ARCH1 of ND2_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_319 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_319;

architecture SYN_ARCH1 of ND2_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_318 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_318;

architecture SYN_ARCH1 of ND2_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_317 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_317;

architecture SYN_ARCH1 of ND2_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_316 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_316;

architecture SYN_ARCH1 of ND2_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_315 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_315;

architecture SYN_ARCH1 of ND2_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_314 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_314;

architecture SYN_ARCH1 of ND2_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_313 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_313;

architecture SYN_ARCH1 of ND2_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_312 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_312;

architecture SYN_ARCH1 of ND2_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_311 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_311;

architecture SYN_ARCH1 of ND2_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_310 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_310;

architecture SYN_ARCH1 of ND2_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_309 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_309;

architecture SYN_ARCH1 of ND2_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_308 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_308;

architecture SYN_ARCH1 of ND2_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_307 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_307;

architecture SYN_ARCH1 of ND2_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_306 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_306;

architecture SYN_ARCH1 of ND2_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_305 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_305;

architecture SYN_ARCH1 of ND2_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_304 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_304;

architecture SYN_ARCH1 of ND2_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_303 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_303;

architecture SYN_ARCH1 of ND2_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_302 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_302;

architecture SYN_ARCH1 of ND2_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_301 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_301;

architecture SYN_ARCH1 of ND2_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_300 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_300;

architecture SYN_ARCH1 of ND2_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_299 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_299;

architecture SYN_ARCH1 of ND2_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_298 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_298;

architecture SYN_ARCH1 of ND2_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_297 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_297;

architecture SYN_ARCH1 of ND2_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_296 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_296;

architecture SYN_ARCH1 of ND2_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_295 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_295;

architecture SYN_ARCH1 of ND2_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_294 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_294;

architecture SYN_ARCH1 of ND2_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_293 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_293;

architecture SYN_ARCH1 of ND2_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_292 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_292;

architecture SYN_ARCH1 of ND2_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_291 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_291;

architecture SYN_ARCH1 of ND2_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_290 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_290;

architecture SYN_ARCH1 of ND2_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_289 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_289;

architecture SYN_ARCH1 of ND2_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_288 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_288;

architecture SYN_ARCH1 of ND2_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_287 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_287;

architecture SYN_ARCH1 of ND2_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_286 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_286;

architecture SYN_ARCH1 of ND2_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_285 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_285;

architecture SYN_ARCH1 of ND2_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_284 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_284;

architecture SYN_ARCH1 of ND2_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_283 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_283;

architecture SYN_ARCH1 of ND2_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_282 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_282;

architecture SYN_ARCH1 of ND2_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_281 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_281;

architecture SYN_ARCH1 of ND2_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_280 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_280;

architecture SYN_ARCH1 of ND2_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_279 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_279;

architecture SYN_ARCH1 of ND2_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_278 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_278;

architecture SYN_ARCH1 of ND2_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_277 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_277;

architecture SYN_ARCH1 of ND2_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_276 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_276;

architecture SYN_ARCH1 of ND2_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_275 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_275;

architecture SYN_ARCH1 of ND2_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_274 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_274;

architecture SYN_ARCH1 of ND2_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_273 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_273;

architecture SYN_ARCH1 of ND2_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_272 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_272;

architecture SYN_ARCH1 of ND2_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_271 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_271;

architecture SYN_ARCH1 of ND2_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_270 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_270;

architecture SYN_ARCH1 of ND2_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_269 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_269;

architecture SYN_ARCH1 of ND2_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_268 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_268;

architecture SYN_ARCH1 of ND2_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_267 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_267;

architecture SYN_ARCH1 of ND2_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_266 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_266;

architecture SYN_ARCH1 of ND2_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_265 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_265;

architecture SYN_ARCH1 of ND2_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_264 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_264;

architecture SYN_ARCH1 of ND2_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_263 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_263;

architecture SYN_ARCH1 of ND2_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_262 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_262;

architecture SYN_ARCH1 of ND2_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_261 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_261;

architecture SYN_ARCH1 of ND2_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_260 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_260;

architecture SYN_ARCH1 of ND2_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_259 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_259;

architecture SYN_ARCH1 of ND2_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_258 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_258;

architecture SYN_ARCH1 of ND2_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_257 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_257;

architecture SYN_ARCH1 of ND2_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_256 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_256;

architecture SYN_ARCH1 of ND2_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_255 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_255;

architecture SYN_ARCH1 of ND2_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_254 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_254;

architecture SYN_ARCH1 of ND2_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_253 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_253;

architecture SYN_ARCH1 of ND2_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_252 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_252;

architecture SYN_ARCH1 of ND2_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_251 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_251;

architecture SYN_ARCH1 of ND2_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_250 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_250;

architecture SYN_ARCH1 of ND2_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_249 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_249;

architecture SYN_ARCH1 of ND2_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_248 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_248;

architecture SYN_ARCH1 of ND2_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_247 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_247;

architecture SYN_ARCH1 of ND2_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_246 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_246;

architecture SYN_ARCH1 of ND2_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_245 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_245;

architecture SYN_ARCH1 of ND2_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_244 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_244;

architecture SYN_ARCH1 of ND2_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_243 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_243;

architecture SYN_ARCH1 of ND2_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_242 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_242;

architecture SYN_ARCH1 of ND2_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_241 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_241;

architecture SYN_ARCH1 of ND2_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_240 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_240;

architecture SYN_ARCH1 of ND2_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_239 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_239;

architecture SYN_ARCH1 of ND2_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_238 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_238;

architecture SYN_ARCH1 of ND2_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_237 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_237;

architecture SYN_ARCH1 of ND2_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_236 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_236;

architecture SYN_ARCH1 of ND2_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_235 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_235;

architecture SYN_ARCH1 of ND2_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_234 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_234;

architecture SYN_ARCH1 of ND2_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_233 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_233;

architecture SYN_ARCH1 of ND2_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_232 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_232;

architecture SYN_ARCH1 of ND2_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_231 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_231;

architecture SYN_ARCH1 of ND2_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_230 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_230;

architecture SYN_ARCH1 of ND2_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_229 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_229;

architecture SYN_ARCH1 of ND2_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_228;

architecture SYN_ARCH1 of ND2_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_227;

architecture SYN_ARCH1 of ND2_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_226;

architecture SYN_ARCH1 of ND2_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_225;

architecture SYN_ARCH1 of ND2_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_224;

architecture SYN_ARCH1 of ND2_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_223;

architecture SYN_ARCH1 of ND2_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_222;

architecture SYN_ARCH1 of ND2_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_221;

architecture SYN_ARCH1 of ND2_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_220;

architecture SYN_ARCH1 of ND2_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_219;

architecture SYN_ARCH1 of ND2_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_218;

architecture SYN_ARCH1 of ND2_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_217;

architecture SYN_ARCH1 of ND2_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_216;

architecture SYN_ARCH1 of ND2_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_215;

architecture SYN_ARCH1 of ND2_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_214;

architecture SYN_ARCH1 of ND2_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_213;

architecture SYN_ARCH1 of ND2_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_212;

architecture SYN_ARCH1 of ND2_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_211;

architecture SYN_ARCH1 of ND2_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_210;

architecture SYN_ARCH1 of ND2_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_209;

architecture SYN_ARCH1 of ND2_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_208;

architecture SYN_ARCH1 of ND2_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_207;

architecture SYN_ARCH1 of ND2_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_206;

architecture SYN_ARCH1 of ND2_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_205;

architecture SYN_ARCH1 of ND2_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_204;

architecture SYN_ARCH1 of ND2_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_203;

architecture SYN_ARCH1 of ND2_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_202;

architecture SYN_ARCH1 of ND2_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_201;

architecture SYN_ARCH1 of ND2_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_200;

architecture SYN_ARCH1 of ND2_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_199;

architecture SYN_ARCH1 of ND2_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_198;

architecture SYN_ARCH1 of ND2_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_197;

architecture SYN_ARCH1 of ND2_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_196;

architecture SYN_ARCH1 of ND2_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_195;

architecture SYN_ARCH1 of ND2_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_194;

architecture SYN_ARCH1 of ND2_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_193;

architecture SYN_ARCH1 of ND2_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_192;

architecture SYN_ARCH1 of ND2_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH1 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH1 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH1 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH1 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH1 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_STRUCTURAL of MUX21_217 is

   component ND2_661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_217 port map( A => S, Y => SB);
   UND1 : ND2_663 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_662 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_661 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_STRUCTURAL of MUX21_216 is

   component ND2_658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_216 port map( A => S, Y => SB);
   UND1 : ND2_660 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_659 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_658 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_STRUCTURAL of MUX21_215 is

   component ND2_655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_215 port map( A => S, Y => SB);
   UND1 : ND2_657 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_656 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_655 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_STRUCTURAL of MUX21_214 is

   component ND2_652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_214 port map( A => S, Y => SB);
   UND1 : ND2_654 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_653 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_652 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_STRUCTURAL of MUX21_213 is

   component ND2_649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_213 port map( A => S, Y => SB);
   UND1 : ND2_651 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_650 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_649 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_STRUCTURAL of MUX21_212 is

   component ND2_646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_212 port map( A => S, Y => SB);
   UND1 : ND2_648 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_647 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_646 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_STRUCTURAL of MUX21_211 is

   component ND2_643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_211 port map( A => S, Y => SB);
   UND1 : ND2_645 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_644 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_643 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_STRUCTURAL of MUX21_210 is

   component ND2_640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_210 port map( A => S, Y => SB);
   UND1 : ND2_642 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_641 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_640 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_STRUCTURAL of MUX21_209 is

   component ND2_637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_209 port map( A => S, Y => SB);
   UND1 : ND2_639 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_638 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_637 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_STRUCTURAL of MUX21_208 is

   component ND2_634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_208 port map( A => S, Y => SB);
   UND1 : ND2_636 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_635 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_634 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_STRUCTURAL of MUX21_207 is

   component ND2_631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_207 port map( A => S, Y => SB);
   UND1 : ND2_633 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_632 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_631 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_STRUCTURAL of MUX21_206 is

   component ND2_628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_206 port map( A => S, Y => SB);
   UND1 : ND2_630 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_629 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_628 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_STRUCTURAL of MUX21_205 is

   component ND2_625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_205 port map( A => S, Y => SB);
   UND1 : ND2_627 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_626 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_625 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_STRUCTURAL of MUX21_204 is

   component ND2_622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_204 port map( A => S, Y => SB);
   UND1 : ND2_624 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_623 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_622 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_STRUCTURAL of MUX21_203 is

   component ND2_619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_203 port map( A => S, Y => SB);
   UND1 : ND2_621 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_620 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_619 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_STRUCTURAL of MUX21_202 is

   component ND2_616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_202 port map( A => S, Y => SB);
   UND1 : ND2_618 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_617 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_616 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_STRUCTURAL of MUX21_201 is

   component ND2_613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_201 port map( A => S, Y => SB);
   UND1 : ND2_615 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_614 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_613 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_STRUCTURAL of MUX21_200 is

   component ND2_610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_200 port map( A => S, Y => SB);
   UND1 : ND2_612 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_611 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_610 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_STRUCTURAL of MUX21_199 is

   component ND2_607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_199 port map( A => S, Y => SB);
   UND1 : ND2_609 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_608 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_607 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_STRUCTURAL of MUX21_198 is

   component ND2_604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_198 port map( A => S, Y => SB);
   UND1 : ND2_606 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_605 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_604 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_STRUCTURAL of MUX21_197 is

   component ND2_601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_197 port map( A => S, Y => SB);
   UND1 : ND2_603 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_602 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_601 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_STRUCTURAL of MUX21_196 is

   component ND2_598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_196 port map( A => S, Y => SB);
   UND1 : ND2_600 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_599 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_598 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_STRUCTURAL of MUX21_195 is

   component ND2_595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_195 port map( A => S, Y => SB);
   UND1 : ND2_597 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_596 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_595 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_STRUCTURAL of MUX21_194 is

   component ND2_592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_194 port map( A => S, Y => SB);
   UND1 : ND2_594 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_593 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_592 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_STRUCTURAL of MUX21_193 is

   component ND2_589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_193 port map( A => S, Y => SB);
   UND1 : ND2_591 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_590 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_589 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_STRUCTURAL of MUX21_192 is

   component ND2_586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_192 port map( A => S, Y => SB);
   UND1 : ND2_588 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_587 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_586 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_STRUCTURAL of MUX21_191 is

   component ND2_583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_191 port map( A => S, Y => SB);
   UND1 : ND2_585 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_584 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_583 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_STRUCTURAL of MUX21_190 is

   component ND2_580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_190 port map( A => S, Y => SB);
   UND1 : ND2_582 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_581 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_580 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_STRUCTURAL of MUX21_189 is

   component ND2_577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_189 port map( A => S, Y => SB);
   UND1 : ND2_579 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_578 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_577 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_STRUCTURAL of MUX21_188 is

   component ND2_574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_188 port map( A => S, Y => SB);
   UND1 : ND2_576 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_575 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_574 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_STRUCTURAL of MUX21_187 is

   component ND2_571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_187 port map( A => S, Y => SB);
   UND1 : ND2_573 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_572 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_571 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_STRUCTURAL of MUX21_186 is

   component ND2_568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_186 port map( A => S, Y => SB);
   UND1 : ND2_570 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_569 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_568 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_STRUCTURAL of MUX21_185 is

   component ND2_565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_185 port map( A => S, Y => SB);
   UND1 : ND2_567 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_566 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_565 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_STRUCTURAL of MUX21_184 is

   component ND2_562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_184 port map( A => S, Y => SB);
   UND1 : ND2_564 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_563 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_562 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_STRUCTURAL of MUX21_183 is

   component ND2_559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_183 port map( A => S, Y => SB);
   UND1 : ND2_561 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_560 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_559 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_STRUCTURAL of MUX21_182 is

   component ND2_556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_182 port map( A => S, Y => SB);
   UND1 : ND2_558 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_557 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_556 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_STRUCTURAL of MUX21_181 is

   component ND2_553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_181 port map( A => S, Y => SB);
   UND1 : ND2_555 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_554 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_553 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_STRUCTURAL of MUX21_180 is

   component ND2_550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_180 port map( A => S, Y => SB);
   UND1 : ND2_552 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_551 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_550 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_STRUCTURAL of MUX21_179 is

   component ND2_547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_179 port map( A => S, Y => SB);
   UND1 : ND2_549 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_548 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_547 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_STRUCTURAL of MUX21_178 is

   component ND2_544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_178 port map( A => S, Y => SB);
   UND1 : ND2_546 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_545 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_544 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_STRUCTURAL of MUX21_177 is

   component ND2_541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_177 port map( A => S, Y => SB);
   UND1 : ND2_543 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_542 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_541 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_STRUCTURAL of MUX21_176 is

   component ND2_538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_176 port map( A => S, Y => SB);
   UND1 : ND2_540 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_539 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_538 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_STRUCTURAL of MUX21_175 is

   component ND2_535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_175 port map( A => S, Y => SB);
   UND1 : ND2_537 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_536 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_535 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_STRUCTURAL of MUX21_174 is

   component ND2_532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_174 port map( A => S, Y => SB);
   UND1 : ND2_534 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_533 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_532 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_STRUCTURAL of MUX21_173 is

   component ND2_529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_173 port map( A => S, Y => SB);
   UND1 : ND2_531 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_530 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_529 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_STRUCTURAL of MUX21_172 is

   component ND2_526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_172 port map( A => S, Y => SB);
   UND1 : ND2_528 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_527 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_526 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_STRUCTURAL of MUX21_171 is

   component ND2_523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_171 port map( A => S, Y => SB);
   UND1 : ND2_525 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_524 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_523 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_STRUCTURAL of MUX21_170 is

   component ND2_520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_170 port map( A => S, Y => SB);
   UND1 : ND2_522 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_521 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_520 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_STRUCTURAL of MUX21_169 is

   component ND2_517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_169 port map( A => S, Y => SB);
   UND1 : ND2_519 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_518 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_517 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_STRUCTURAL of MUX21_168 is

   component ND2_514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_168 port map( A => S, Y => SB);
   UND1 : ND2_516 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_515 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_514 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_STRUCTURAL of MUX21_167 is

   component ND2_511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_167 port map( A => S, Y => SB);
   UND1 : ND2_513 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_512 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_511 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_STRUCTURAL of MUX21_166 is

   component ND2_508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_166 port map( A => S, Y => SB);
   UND1 : ND2_510 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_509 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_508 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_STRUCTURAL of MUX21_165 is

   component ND2_505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_165 port map( A => S, Y => SB);
   UND1 : ND2_507 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_506 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_505 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_STRUCTURAL of MUX21_164 is

   component ND2_502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_164 port map( A => S, Y => SB);
   UND1 : ND2_504 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_503 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_502 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_STRUCTURAL of MUX21_163 is

   component ND2_499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_163 port map( A => S, Y => SB);
   UND1 : ND2_501 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_500 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_499 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_STRUCTURAL of MUX21_162 is

   component ND2_496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_162 port map( A => S, Y => SB);
   UND1 : ND2_498 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_497 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_496 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_STRUCTURAL of MUX21_161 is

   component ND2_493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_161 port map( A => S, Y => SB);
   UND1 : ND2_495 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_494 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_493 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_STRUCTURAL of MUX21_160 is

   component ND2_490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_160 port map( A => S, Y => SB);
   UND1 : ND2_492 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_491 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_490 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_STRUCTURAL of MUX21_159 is

   component ND2_487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_159 port map( A => S, Y => SB);
   UND1 : ND2_489 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_488 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_487 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_STRUCTURAL of MUX21_158 is

   component ND2_484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_158 port map( A => S, Y => SB);
   UND1 : ND2_486 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_485 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_484 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_STRUCTURAL of MUX21_157 is

   component ND2_481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_157 port map( A => S, Y => SB);
   UND1 : ND2_483 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_482 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_481 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_STRUCTURAL of MUX21_156 is

   component ND2_478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_156 port map( A => S, Y => SB);
   UND1 : ND2_480 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_479 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_478 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_STRUCTURAL of MUX21_155 is

   component ND2_475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_155 port map( A => S, Y => SB);
   UND1 : ND2_477 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_476 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_475 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_STRUCTURAL of MUX21_154 is

   component ND2_472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_154 port map( A => S, Y => SB);
   UND1 : ND2_474 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_473 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_472 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_STRUCTURAL of MUX21_153 is

   component ND2_469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_153 port map( A => S, Y => SB);
   UND1 : ND2_471 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_470 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_469 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_STRUCTURAL of MUX21_152 is

   component ND2_466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_152 port map( A => S, Y => SB);
   UND1 : ND2_468 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_467 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_466 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_STRUCTURAL of MUX21_151 is

   component ND2_463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_151 port map( A => S, Y => SB);
   UND1 : ND2_465 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_464 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_463 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_STRUCTURAL of MUX21_150 is

   component ND2_460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_150 port map( A => S, Y => SB);
   UND1 : ND2_462 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_461 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_460 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_STRUCTURAL of MUX21_149 is

   component ND2_457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_149 port map( A => S, Y => SB);
   UND1 : ND2_459 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_458 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_457 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_STRUCTURAL of MUX21_148 is

   component ND2_454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_148 port map( A => S, Y => SB);
   UND1 : ND2_456 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_455 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_454 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_STRUCTURAL of MUX21_147 is

   component ND2_451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_147 port map( A => S, Y => SB);
   UND1 : ND2_453 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_452 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_451 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_STRUCTURAL of MUX21_146 is

   component ND2_448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_146 port map( A => S, Y => SB);
   UND1 : ND2_450 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_449 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_448 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_STRUCTURAL of MUX21_145 is

   component ND2_445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_145 port map( A => S, Y => SB);
   UND1 : ND2_447 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_446 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_445 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_STRUCTURAL of MUX21_144 is

   component ND2_442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_144 port map( A => S, Y => SB);
   UND1 : ND2_444 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_443 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_442 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_STRUCTURAL of MUX21_143 is

   component ND2_439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_143 port map( A => S, Y => SB);
   UND1 : ND2_441 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_440 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_439 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_STRUCTURAL of MUX21_142 is

   component ND2_436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_142 port map( A => S, Y => SB);
   UND1 : ND2_438 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_437 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_436 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_STRUCTURAL of MUX21_141 is

   component ND2_433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_141 port map( A => S, Y => SB);
   UND1 : ND2_435 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_434 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_433 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_STRUCTURAL of MUX21_140 is

   component ND2_430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_140 port map( A => S, Y => SB);
   UND1 : ND2_432 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_431 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_430 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_STRUCTURAL of MUX21_139 is

   component ND2_427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_139 port map( A => S, Y => SB);
   UND1 : ND2_429 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_428 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_427 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_STRUCTURAL of MUX21_138 is

   component ND2_424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_138 port map( A => S, Y => SB);
   UND1 : ND2_426 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_425 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_424 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_STRUCTURAL of MUX21_137 is

   component ND2_421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_137 port map( A => S, Y => SB);
   UND1 : ND2_423 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_422 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_421 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_STRUCTURAL of MUX21_136 is

   component ND2_418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_136 port map( A => S, Y => SB);
   UND1 : ND2_420 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_419 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_418 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_STRUCTURAL of MUX21_135 is

   component ND2_415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_135 port map( A => S, Y => SB);
   UND1 : ND2_417 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_416 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_415 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_STRUCTURAL of MUX21_134 is

   component ND2_412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_134 port map( A => S, Y => SB);
   UND1 : ND2_414 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_413 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_412 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_STRUCTURAL of MUX21_133 is

   component ND2_409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_133 port map( A => S, Y => SB);
   UND1 : ND2_411 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_410 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_409 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_STRUCTURAL of MUX21_132 is

   component ND2_406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_132 port map( A => S, Y => SB);
   UND1 : ND2_408 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_407 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_406 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_STRUCTURAL of MUX21_131 is

   component ND2_403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_131 port map( A => S, Y => SB);
   UND1 : ND2_405 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_404 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_403 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_STRUCTURAL of MUX21_130 is

   component ND2_400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_130 port map( A => S, Y => SB);
   UND1 : ND2_402 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_401 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_400 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_STRUCTURAL of MUX21_129 is

   component ND2_397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_129 port map( A => S, Y => SB);
   UND1 : ND2_399 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_398 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_397 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_STRUCTURAL of MUX21_128 is

   component ND2_394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_128 port map( A => S, Y => SB);
   UND1 : ND2_396 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_395 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_394 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_STRUCTURAL of MUX21_127 is

   component ND2_391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_127 port map( A => S, Y => SB);
   UND1 : ND2_393 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_392 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_391 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_STRUCTURAL of MUX21_126 is

   component ND2_388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_126 port map( A => S, Y => SB);
   UND1 : ND2_390 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_389 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_388 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_STRUCTURAL of MUX21_125 is

   component ND2_385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_125 port map( A => S, Y => SB);
   UND1 : ND2_387 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_386 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_385 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_STRUCTURAL of MUX21_124 is

   component ND2_382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_124 port map( A => S, Y => SB);
   UND1 : ND2_384 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_383 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_382 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_STRUCTURAL of MUX21_123 is

   component ND2_379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_123 port map( A => S, Y => SB);
   UND1 : ND2_381 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_380 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_379 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_STRUCTURAL of MUX21_122 is

   component ND2_376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_122 port map( A => S, Y => SB);
   UND1 : ND2_378 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_377 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_376 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_STRUCTURAL of MUX21_121 is

   component ND2_373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_121 port map( A => S, Y => SB);
   UND1 : ND2_375 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_374 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_373 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_STRUCTURAL of MUX21_120 is

   component ND2_370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_120 port map( A => S, Y => SB);
   UND1 : ND2_372 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_371 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_370 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_STRUCTURAL of MUX21_119 is

   component ND2_367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_119 port map( A => S, Y => SB);
   UND1 : ND2_369 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_368 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_367 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_STRUCTURAL of MUX21_118 is

   component ND2_364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_118 port map( A => S, Y => SB);
   UND1 : ND2_366 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_365 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_364 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_STRUCTURAL of MUX21_117 is

   component ND2_361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_117 port map( A => S, Y => SB);
   UND1 : ND2_363 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_362 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_361 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_STRUCTURAL of MUX21_116 is

   component ND2_358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_116 port map( A => S, Y => SB);
   UND1 : ND2_360 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_359 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_358 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_STRUCTURAL of MUX21_115 is

   component ND2_355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_115 port map( A => S, Y => SB);
   UND1 : ND2_357 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_356 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_355 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_STRUCTURAL of MUX21_114 is

   component ND2_352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_114 port map( A => S, Y => SB);
   UND1 : ND2_354 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_353 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_352 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_STRUCTURAL of MUX21_113 is

   component ND2_349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_113 port map( A => S, Y => SB);
   UND1 : ND2_351 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_350 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_349 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_STRUCTURAL of MUX21_112 is

   component ND2_346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_112 port map( A => S, Y => SB);
   UND1 : ND2_348 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_347 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_346 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_STRUCTURAL of MUX21_111 is

   component ND2_343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_111 port map( A => S, Y => SB);
   UND1 : ND2_345 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_344 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_343 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_STRUCTURAL of MUX21_110 is

   component ND2_340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_110 port map( A => S, Y => SB);
   UND1 : ND2_342 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_341 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_340 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_STRUCTURAL of MUX21_109 is

   component ND2_337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_109 port map( A => S, Y => SB);
   UND1 : ND2_339 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_338 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_337 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_STRUCTURAL of MUX21_108 is

   component ND2_334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_108 port map( A => S, Y => SB);
   UND1 : ND2_336 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_335 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_334 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_STRUCTURAL of MUX21_107 is

   component ND2_331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_107 port map( A => S, Y => SB);
   UND1 : ND2_333 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_332 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_331 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_STRUCTURAL of MUX21_106 is

   component ND2_328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_106 port map( A => S, Y => SB);
   UND1 : ND2_330 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_329 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_328 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_STRUCTURAL of MUX21_105 is

   component ND2_325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_105 port map( A => S, Y => SB);
   UND1 : ND2_327 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_326 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_325 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_STRUCTURAL of MUX21_104 is

   component ND2_322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_104 port map( A => S, Y => SB);
   UND1 : ND2_324 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_323 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_322 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_STRUCTURAL of MUX21_103 is

   component ND2_319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_103 port map( A => S, Y => SB);
   UND1 : ND2_321 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_320 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_319 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_STRUCTURAL of MUX21_102 is

   component ND2_316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_102 port map( A => S, Y => SB);
   UND1 : ND2_318 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_317 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_316 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_STRUCTURAL of MUX21_101 is

   component ND2_313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_101 port map( A => S, Y => SB);
   UND1 : ND2_315 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_314 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_313 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_STRUCTURAL of MUX21_100 is

   component ND2_310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_100 port map( A => S, Y => SB);
   UND1 : ND2_312 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_311 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_310 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_STRUCTURAL of MUX21_99 is

   component ND2_307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_99 port map( A => S, Y => SB);
   UND1 : ND2_309 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_308 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_307 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_STRUCTURAL of MUX21_98 is

   component ND2_304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_98 port map( A => S, Y => SB);
   UND1 : ND2_306 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_305 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_304 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_STRUCTURAL of MUX21_97 is

   component ND2_301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_97 port map( A => S, Y => SB);
   UND1 : ND2_303 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_302 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_301 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_STRUCTURAL of MUX21_96 is

   component ND2_298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_96 port map( A => S, Y => SB);
   UND1 : ND2_300 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_299 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_298 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_STRUCTURAL of MUX21_95 is

   component ND2_295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_95 port map( A => S, Y => SB);
   UND1 : ND2_297 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_296 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_295 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_STRUCTURAL of MUX21_94 is

   component ND2_292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_94 port map( A => S, Y => SB);
   UND1 : ND2_294 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_293 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_292 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_STRUCTURAL of MUX21_93 is

   component ND2_289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_93 port map( A => S, Y => SB);
   UND1 : ND2_291 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_290 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_289 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_STRUCTURAL of MUX21_92 is

   component ND2_286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_92 port map( A => S, Y => SB);
   UND1 : ND2_288 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_287 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_286 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_STRUCTURAL of MUX21_91 is

   component ND2_283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_91 port map( A => S, Y => SB);
   UND1 : ND2_285 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_284 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_283 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_STRUCTURAL of MUX21_90 is

   component ND2_280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_90 port map( A => S, Y => SB);
   UND1 : ND2_282 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_281 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_280 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_STRUCTURAL of MUX21_89 is

   component ND2_277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_89 port map( A => S, Y => SB);
   UND1 : ND2_279 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_278 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_277 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_STRUCTURAL of MUX21_88 is

   component ND2_274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_88 port map( A => S, Y => SB);
   UND1 : ND2_276 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_275 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_274 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_STRUCTURAL of MUX21_87 is

   component ND2_271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_87 port map( A => S, Y => SB);
   UND1 : ND2_273 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_272 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_271 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_STRUCTURAL of MUX21_86 is

   component ND2_268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_86 port map( A => S, Y => SB);
   UND1 : ND2_270 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_269 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_268 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_STRUCTURAL of MUX21_85 is

   component ND2_265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_85 port map( A => S, Y => SB);
   UND1 : ND2_267 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_266 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_265 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_STRUCTURAL of MUX21_84 is

   component ND2_262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_84 port map( A => S, Y => SB);
   UND1 : ND2_264 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_263 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_262 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_STRUCTURAL of MUX21_83 is

   component ND2_259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_83 port map( A => S, Y => SB);
   UND1 : ND2_261 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_260 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_259 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_STRUCTURAL of MUX21_82 is

   component ND2_256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_82 port map( A => S, Y => SB);
   UND1 : ND2_258 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_257 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_256 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_STRUCTURAL of MUX21_81 is

   component ND2_253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_81 port map( A => S, Y => SB);
   UND1 : ND2_255 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_254 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_253 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_STRUCTURAL of MUX21_80 is

   component ND2_250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_80 port map( A => S, Y => SB);
   UND1 : ND2_252 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_251 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_250 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_STRUCTURAL of MUX21_79 is

   component ND2_247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_79 port map( A => S, Y => SB);
   UND1 : ND2_249 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_248 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_247 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_STRUCTURAL of MUX21_78 is

   component ND2_244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_78 port map( A => S, Y => SB);
   UND1 : ND2_246 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_245 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_244 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_STRUCTURAL of MUX21_77 is

   component ND2_241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_77 port map( A => S, Y => SB);
   UND1 : ND2_243 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_242 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_241 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_STRUCTURAL of MUX21_76 is

   component ND2_238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_76 port map( A => S, Y => SB);
   UND1 : ND2_240 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_239 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_238 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_STRUCTURAL of MUX21_75 is

   component ND2_235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_75 port map( A => S, Y => SB);
   UND1 : ND2_237 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_236 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_235 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_STRUCTURAL of MUX21_74 is

   component ND2_232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_74 port map( A => S, Y => SB);
   UND1 : ND2_234 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_233 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_232 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_STRUCTURAL of MUX21_73 is

   component ND2_229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_73 port map( A => S, Y => SB);
   UND1 : ND2_231 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_230 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_229 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_STRUCTURAL of MUX21_72 is

   component ND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_72 port map( A => S, Y => SB);
   UND1 : ND2_228 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_227 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_226 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_STRUCTURAL of MUX21_71 is

   component ND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_71 port map( A => S, Y => SB);
   UND1 : ND2_225 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_224 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_223 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_STRUCTURAL of MUX21_70 is

   component ND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_70 port map( A => S, Y => SB);
   UND1 : ND2_222 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_221 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_220 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_STRUCTURAL of MUX21_69 is

   component ND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_69 port map( A => S, Y => SB);
   UND1 : ND2_219 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_218 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_217 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_STRUCTURAL of MUX21_68 is

   component ND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_68 port map( A => S, Y => SB);
   UND1 : ND2_216 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_215 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_214 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_STRUCTURAL of MUX21_67 is

   component ND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_67 port map( A => S, Y => SB);
   UND1 : ND2_213 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_212 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_211 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_STRUCTURAL of MUX21_66 is

   component ND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_66 port map( A => S, Y => SB);
   UND1 : ND2_210 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_209 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_208 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_STRUCTURAL of MUX21_65 is

   component ND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_65 port map( A => S, Y => SB);
   UND1 : ND2_207 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_206 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_205 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_STRUCTURAL of MUX21_64 is

   component ND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_64 port map( A => S, Y => SB);
   UND1 : ND2_204 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_203 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_202 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_STRUCTURAL of MUX21_63 is

   component ND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_63 port map( A => S, Y => SB);
   UND1 : ND2_201 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_200 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_199 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_STRUCTURAL of MUX21_62 is

   component ND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_62 port map( A => S, Y => SB);
   UND1 : ND2_198 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_197 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_196 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_STRUCTURAL of MUX21_61 is

   component ND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_61 port map( A => S, Y => SB);
   UND1 : ND2_195 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_194 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_193 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_192 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_191 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_190 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_189 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N2_1 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (1 downto 0);  
         d_out : out std_logic_vector (1 downto 0));

end reg_N2_1;

architecture SYN_behav of reg_N2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, n1, n3_port : std_logic;

begin
   
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n1);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n3_port);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in(1), ZN => N3);
   U4 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_31 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_31;

architecture SYN_behav of ff_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_30 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_30;

architecture SYN_behav of ff_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_29 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_29;

architecture SYN_behav of ff_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_28 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_28;

architecture SYN_behav of ff_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_27 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_27;

architecture SYN_behav of ff_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_26 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_26;

architecture SYN_behav of ff_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_25 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_25;

architecture SYN_behav of ff_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_24 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_24;

architecture SYN_behav of ff_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_23 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_23;

architecture SYN_behav of ff_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_22 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_22;

architecture SYN_behav of ff_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_21 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_21;

architecture SYN_behav of ff_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_20 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_20;

architecture SYN_behav of ff_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_19 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_19;

architecture SYN_behav of ff_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_18 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_18;

architecture SYN_behav of ff_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_17 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_17;

architecture SYN_behav of ff_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_16 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_16;

architecture SYN_behav of ff_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_15 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_15;

architecture SYN_behav of ff_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_14 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_14;

architecture SYN_behav of ff_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_13 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_13;

architecture SYN_behav of ff_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_12 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_12;

architecture SYN_behav of ff_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_11 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_11;

architecture SYN_behav of ff_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_10 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_10;

architecture SYN_behav of ff_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_9 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_9;

architecture SYN_behav of ff_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_8 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_8;

architecture SYN_behav of ff_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_7 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_7;

architecture SYN_behav of ff_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_6 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_6;

architecture SYN_behav of ff_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_5 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_5;

architecture SYN_behav of ff_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_4 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_4;

architecture SYN_behav of ff_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_3 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_3;

architecture SYN_behav of ff_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_2 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_2;

architecture SYN_behav of ff_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_1 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_1;

architecture SYN_behav of ff_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_4;

architecture SYN_struct of MUX21_GENERIC_N32_4 is

   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_186 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_185 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_184 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_183 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   M_4 : MUX21_182 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   M_5 : MUX21_181 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   M_6 : MUX21_180 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   M_7 : MUX21_179 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   M_8 : MUX21_178 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   M_9 : MUX21_177 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   M_10 : MUX21_176 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   M_11 : MUX21_175 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   M_12 : MUX21_174 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   M_13 : MUX21_173 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   M_14 : MUX21_172 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   M_15 : MUX21_171 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   M_16 : MUX21_170 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   M_17 : MUX21_169 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   M_18 : MUX21_168 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   M_19 : MUX21_167 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   M_20 : MUX21_166 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   M_21 : MUX21_165 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   M_22 : MUX21_164 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   M_23 : MUX21_163 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   M_24 : MUX21_162 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   M_25 : MUX21_161 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   M_26 : MUX21_160 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   M_27 : MUX21_159 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   M_28 : MUX21_158 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   M_29 : MUX21_157 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   M_30 : MUX21_156 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   M_31 : MUX21_155 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_3;

architecture SYN_struct of MUX21_GENERIC_N32_3 is

   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_154 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_153 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_152 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_151 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   M_4 : MUX21_150 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   M_5 : MUX21_149 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   M_6 : MUX21_148 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   M_7 : MUX21_147 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   M_8 : MUX21_146 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   M_9 : MUX21_145 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   M_10 : MUX21_144 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   M_11 : MUX21_143 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   M_12 : MUX21_142 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   M_13 : MUX21_141 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   M_14 : MUX21_140 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   M_15 : MUX21_139 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   M_16 : MUX21_138 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   M_17 : MUX21_137 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   M_18 : MUX21_136 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   M_19 : MUX21_135 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   M_20 : MUX21_134 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   M_21 : MUX21_133 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   M_22 : MUX21_132 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   M_23 : MUX21_131 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   M_24 : MUX21_130 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   M_25 : MUX21_129 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   M_26 : MUX21_128 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   M_27 : MUX21_127 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   M_28 : MUX21_126 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   M_29 : MUX21_125 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   M_30 : MUX21_124 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   M_31 : MUX21_123 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_2;

architecture SYN_struct of MUX21_GENERIC_N32_2 is

   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_122 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_121 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_120 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_119 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   M_4 : MUX21_118 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   M_5 : MUX21_117 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   M_6 : MUX21_116 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   M_7 : MUX21_115 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   M_8 : MUX21_114 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   M_9 : MUX21_113 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   M_10 : MUX21_112 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   M_11 : MUX21_111 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   M_12 : MUX21_110 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   M_13 : MUX21_109 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   M_14 : MUX21_108 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   M_15 : MUX21_107 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   M_16 : MUX21_106 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   M_17 : MUX21_105 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   M_18 : MUX21_104 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   M_19 : MUX21_103 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   M_20 : MUX21_102 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   M_21 : MUX21_101 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   M_22 : MUX21_100 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   M_23 : MUX21_99 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   M_24 : MUX21_98 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   M_25 : MUX21_97 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   M_26 : MUX21_96 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   M_27 : MUX21_95 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   M_28 : MUX21_94 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   M_29 : MUX21_93 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   M_30 : MUX21_92 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   M_31 : MUX21_91 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_7 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_7;

architecture SYN_behav of reg_N32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U9 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U10 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U11 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U12 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U13 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U14 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U15 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U16 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U17 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U18 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U19 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U20 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U21 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U22 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U23 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U24 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U25 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U26 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U27 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U28 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U29 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U30 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U31 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U32 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U33 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U34 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U35 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U36 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U37 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_2 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_2;

architecture SYN_behav of reg_N32_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U9 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U10 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U11 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U12 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U13 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U14 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U15 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U16 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U17 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U18 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U19 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U20 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U21 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U22 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U23 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U24 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U25 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U26 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U27 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U28 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U29 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U30 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U31 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U32 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U33 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U34 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U35 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U36 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U37 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_12 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_12;

architecture SYN_behav of reg_N32_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_11 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_11;

architecture SYN_behav of reg_N32_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_9 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_9;

architecture SYN_behav of reg_N32_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_8 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_8;

architecture SYN_behav of reg_N32_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_3 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_3;

architecture SYN_behav of reg_N32_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_1 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_1;

architecture SYN_behav of reg_N32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH1 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH1 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH1 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH1 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH1 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH1 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH1 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH1 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH1 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH1 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH1 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH1 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH1 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH1 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH1 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH1 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH1 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH1 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH1 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH1 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH1 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH1 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH1 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH1 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH1 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH1 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH1 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH1 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH1 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH1 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH1 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH1 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH1 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH1 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH1 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH1 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH1 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH1 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH1 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH1 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH1 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH1 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH1 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH1 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH1 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH1 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH1 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH1 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH1 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH1 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH1 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH1 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH1 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH1 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH1 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH1 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH1 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH1 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH1 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH1 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH1 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH1 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH1 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH1 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH1 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH1 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH1 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH1 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH1 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH1 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH1 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH1 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH1 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH1 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH1 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH1 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH1 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH1 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH1 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH1 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH1 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH1 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH1 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH1 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH1 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH1 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH1 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH1 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH1 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH1 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_30_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30_1;

architecture SYN_BEHAVIORAL of IV_30_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH1 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH1 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH1 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_31_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31_1;

architecture SYN_BEHAVIORAL of IV_31_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_94_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94_1;

architecture SYN_ARCH1 of ND2_94_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_95_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95_1;

architecture SYN_ARCH1 of ND2_95_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_0_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0_1;

architecture SYN_ARCH1 of ND2_0_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_0_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0_1;

architecture SYN_BEHAVIORAL of IV_0_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH1 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH1 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH1 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH1 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH1 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH1 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH1 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH1 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH1 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH1 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH1 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH1 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH1 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH1 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH1 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH1 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH1 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH1 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH1 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH1 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH1 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH1 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH1 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH1 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH1 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH1 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH1 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH1 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH1 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH1 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH1 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH1 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH1 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH1 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH1 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH1 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH1 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH1 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH1 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH1 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH1 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH1 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH1 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH1 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH1 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH1 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH1 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH1 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH1 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH1 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH1 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH1 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH1 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH1 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH1 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH1 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH1 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH1 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH1 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH1 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH1 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH1 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH1 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH1 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH1 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH1 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH1 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH1 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH1 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH1 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH1 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH1 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH1 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH1 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH1 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH1 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH1 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH1 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH1 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH1 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH1 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH1 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH1 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH1 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH1 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH1 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH1 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH1 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH1 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH1 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_30_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30_0;

architecture SYN_BEHAVIORAL of IV_30_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH1 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH1 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH1 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_31_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31_0;

architecture SYN_BEHAVIORAL of IV_31_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_94_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94_0;

architecture SYN_ARCH1 of ND2_94_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_95_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95_0;

architecture SYN_ARCH1 of ND2_95_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_0_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0_0;

architecture SYN_ARCH1 of ND2_0_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_0_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0_0;

architecture SYN_BEHAVIORAL of IV_0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n17, n18 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n18, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n18);
   U1 : INV_X1 port map( A => n17, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n18, B2 => Ci, ZN => n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_30_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30_1;

architecture SYN_STRUCTURAL of MUX21_30_1 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30_1 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_31_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31_1;

architecture SYN_STRUCTURAL of MUX21_31_1 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31_1 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_0_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0_1;

architecture SYN_STRUCTURAL of MUX21_0_1 is

   component ND2_94_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0_1 port map( A => S, Y => SB);
   UND1 : ND2_0_1 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95_1 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_62_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62_1;

architecture SYN_BEHAVIORAL of FA_62_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_63_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63_1;

architecture SYN_BEHAVIORAL of FA_63_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_0_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_1;

architecture SYN_BEHAVIORAL of FA_0_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n7, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_98 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_97 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_96 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_101 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_100 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_99 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_104 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_103 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_102 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_107 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_106 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_105 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_110 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_109 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_108 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_113 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_112 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_111 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_116 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_115 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_114 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_119 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_118 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_117 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_122 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_121 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_120 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_125 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_124 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_123 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_128 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_127 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_126 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_131 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_130 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_129 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_134 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_133 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_132 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_137 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_136 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_135 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_140 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_139 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_138 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_143 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_142 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_141 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_146 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_145 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_144 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_149 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_148 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_147 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_152 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_151 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_150 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_155 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_154 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_153 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_158 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_157 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_156 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_161 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_160 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_159 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_164 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_163 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_162 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_167 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_166 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_165 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_170 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_169 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_168 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_173 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_172 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_171 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_176 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_175 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_174 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_179 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_178 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_177 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_182 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_181 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_180 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_30_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30_0;

architecture SYN_STRUCTURAL of MUX21_30_0 is

   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30_0 port map( A => S, Y => SB);
   UND1 : ND2_185 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_184 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_183 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_31_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31_0;

architecture SYN_STRUCTURAL of MUX21_31_0 is

   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31_0 port map( A => S, Y => SB);
   UND1 : ND2_188 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_187 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_186 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_0_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0_0;

architecture SYN_STRUCTURAL of MUX21_0_0 is

   component ND2_94_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0_0 port map( A => S, Y => SB);
   UND1 : ND2_0_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95_0 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94_0 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_62_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62_0;

architecture SYN_BEHAVIORAL of FA_62_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_63_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63_0;

architecture SYN_BEHAVIORAL of FA_63_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_0_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_0;

architecture SYN_BEHAVIORAL of FA_0_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2;

architecture SYN_ARCH1 of ND2 is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0 : std_logic;

begin
   
   I_0 : GTECH_NOT port map( A => N0, Z => Y);
   C7 : GTECH_AND2 port map( A => A, B => B, Z => N0);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV is

   port( A : in std_logic;  Y : out std_logic);

end IV;

architecture SYN_BEHAVIORAL of IV is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;

begin
   
   I_0 : GTECH_NOT port map( A => A, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_1;

architecture SYN_struct of MUX21_GENERIC_N4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_1;

architecture SYN_STRUCTURAL of rca_generic_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_2;

architecture SYN_STRUCTURAL of rca_generic_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_2;

architecture SYN_struct of MUX21_GENERIC_N4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_3;

architecture SYN_STRUCTURAL of rca_generic_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_4;

architecture SYN_STRUCTURAL of rca_generic_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_3;

architecture SYN_struct of MUX21_GENERIC_N4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_5;

architecture SYN_STRUCTURAL of rca_generic_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_6;

architecture SYN_STRUCTURAL of rca_generic_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_4;

architecture SYN_struct of MUX21_GENERIC_N4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_7;

architecture SYN_STRUCTURAL of rca_generic_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_8;

architecture SYN_STRUCTURAL of rca_generic_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_5;

architecture SYN_struct of MUX21_GENERIC_N4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_9;

architecture SYN_STRUCTURAL of rca_generic_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_10;

architecture SYN_STRUCTURAL of rca_generic_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_6_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6_1;

architecture SYN_struct of MUX21_GENERIC_N4_6_1 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_11;

architecture SYN_STRUCTURAL of rca_generic_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_12;

architecture SYN_STRUCTURAL of rca_generic_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_7_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7_1;

architecture SYN_struct of MUX21_GENERIC_N4_7_1 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_13;

architecture SYN_STRUCTURAL of rca_generic_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_14_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_14_1;

architecture SYN_STRUCTURAL of rca_generic_N4_14_1 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0_1;

architecture SYN_struct of MUX21_GENERIC_N4_0_1 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_0_1 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_31_1 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_30_1 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_15_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_15_1;

architecture SYN_STRUCTURAL of rca_generic_N4_15_1 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_0_1;

architecture SYN_STRUCTURAL of rca_generic_N4_0_1 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0_1 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63_1 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_62_1 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_8;

architecture SYN_struct of MUX21_GENERIC_N4_8 is

   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_35 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_34 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_33 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_32 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_16;

architecture SYN_STRUCTURAL of rca_generic_N4_16 is

   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_259 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_258 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_257 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_256 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_17;

architecture SYN_STRUCTURAL of rca_generic_N4_17 is

   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_263 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_262 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_261 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_260 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_9;

architecture SYN_struct of MUX21_GENERIC_N4_9 is

   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_39 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_38 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_37 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_36 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_18;

architecture SYN_STRUCTURAL of rca_generic_N4_18 is

   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_267 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_266 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_265 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_264 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_19;

architecture SYN_STRUCTURAL of rca_generic_N4_19 is

   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_271 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_270 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_269 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_268 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_10;

architecture SYN_struct of MUX21_GENERIC_N4_10 is

   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_43 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_42 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_41 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_40 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_20;

architecture SYN_STRUCTURAL of rca_generic_N4_20 is

   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_275 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_274 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_273 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_272 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_21;

architecture SYN_STRUCTURAL of rca_generic_N4_21 is

   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_279 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_278 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_277 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_276 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_11;

architecture SYN_struct of MUX21_GENERIC_N4_11 is

   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_47 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_46 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_45 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_44 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_22;

architecture SYN_STRUCTURAL of rca_generic_N4_22 is

   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_283 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_282 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_281 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_280 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_23;

architecture SYN_STRUCTURAL of rca_generic_N4_23 is

   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_287 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_286 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_285 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_284 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_12;

architecture SYN_struct of MUX21_GENERIC_N4_12 is

   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_51 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_50 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_49 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_48 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_24;

architecture SYN_STRUCTURAL of rca_generic_N4_24 is

   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_291 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_290 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_289 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_288 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_25;

architecture SYN_STRUCTURAL of rca_generic_N4_25 is

   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_295 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_294 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_293 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_292 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_6_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6_0;

architecture SYN_struct of MUX21_GENERIC_N4_6_0 is

   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_55 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_54 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_53 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_52 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_26;

architecture SYN_STRUCTURAL of rca_generic_N4_26 is

   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_299 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_298 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_297 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_296 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_27;

architecture SYN_STRUCTURAL of rca_generic_N4_27 is

   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_303 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_302 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_301 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_300 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_7_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7_0;

architecture SYN_struct of MUX21_GENERIC_N4_7_0 is

   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_59 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_58 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_57 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_56 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_28;

architecture SYN_STRUCTURAL of rca_generic_N4_28 is

   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_307 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_306 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_305 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_304 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_14_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_14_0;

architecture SYN_STRUCTURAL of rca_generic_N4_14_0 is

   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_311 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_310 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_309 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_308 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0_0;

architecture SYN_struct of MUX21_GENERIC_N4_0_0 is

   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_0_0 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_31_0 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_30_0 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_60 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_15_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_15_0;

architecture SYN_STRUCTURAL of rca_generic_N4_15_0 is

   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_315 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_314 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_313 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_312 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_0_0;

architecture SYN_STRUCTURAL of rca_generic_N4_0_0 is

   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63_0 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_62_0 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_316 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_STRUCTURAL of MUX21 is

   component ND2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV port map( A => S, Y => SB);
   UND1 : ND2 port map( A => A, B => S, Y => Y1);
   UND2 : ND2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA;

architecture SYN_BEHAVIORAL of FA is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_XOR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0, N1, N2, N3, N4 : std_logic;

begin
   
   C7 : GTECH_XOR2 port map( A => N0, B => Ci, Z => S);
   C8 : GTECH_XOR2 port map( A => A, B => B, Z => N0);
   C9 : GTECH_OR2 port map( A => N3, B => N4, Z => Co);
   C10 : GTECH_OR2 port map( A => N1, B => N2, Z => N3);
   C11 : GTECH_AND2 port map( A => A, B => B, Z => N1);
   C12 : GTECH_AND2 port map( A => B, B => Ci, Z => N2);
   C13 : GTECH_AND2 port map( A => A, B => Ci, Z => N4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_1;

architecture SYN_STRUCTURAL of carry_select_N4_1 is

   component MUX21_GENERIC_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_2;

architecture SYN_STRUCTURAL of carry_select_N4_2 is

   component MUX21_GENERIC_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_2 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_3;

architecture SYN_STRUCTURAL of carry_select_N4_3 is

   component MUX21_GENERIC_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_3 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_4;

architecture SYN_STRUCTURAL of carry_select_N4_4 is

   component MUX21_GENERIC_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_4 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_5;

architecture SYN_STRUCTURAL of carry_select_N4_5 is

   component MUX21_GENERIC_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_5 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_6_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_6_1;

architecture SYN_STRUCTURAL of carry_select_N4_6_1 is

   component MUX21_GENERIC_N4_6_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_6_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_7_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_7_1;

architecture SYN_STRUCTURAL of carry_select_N4_7_1 is

   component MUX21_GENERIC_N4_7_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_14_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_14_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_7_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_0_1;

architecture SYN_STRUCTURAL of carry_select_N4_0_1 is

   component MUX21_GENERIC_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_15_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_15_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_0_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_3 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_3;

architecture SYN_STRUCTURAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_4 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_4;

architecture SYN_STRUCTURAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_7 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_7;

architecture SYN_STRUCTURAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_9 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_9;

architecture SYN_STRUCTURAL of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_2 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_2;

architecture SYN_STRUCTURAL of PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_1;

architecture SYN_STRUCTURAL of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_5_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_5_1;

architecture SYN_STRUCTURAL of G_5_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_6_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_6_1;

architecture SYN_STRUCTURAL of G_6_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n6);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_3 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_3;

architecture SYN_STRUCTURAL of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_4_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_4_1;

architecture SYN_STRUCTURAL of PG_4_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n6);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_13 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_13;

architecture SYN_STRUCTURAL of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_1;

architecture SYN_STRUCTURAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n11 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n11);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_5 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_5;

architecture SYN_STRUCTURAL of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_6 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_6;

architecture SYN_STRUCTURAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_14 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_14;

architecture SYN_STRUCTURAL of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_15 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_15;

architecture SYN_STRUCTURAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_16 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_16;

architecture SYN_STRUCTURAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_17 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_17;

architecture SYN_STRUCTURAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_19 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_19;

architecture SYN_STRUCTURAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U2 : INV_X1 port map( A => n8, ZN => gout);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_8_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_8_1;

architecture SYN_STRUCTURAL of G_8_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n6);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_7 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_7;

architecture SYN_STRUCTURAL of PG_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_8 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_8;

architecture SYN_STRUCTURAL of PG_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_9 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_9;

architecture SYN_STRUCTURAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_10 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_10;

architecture SYN_STRUCTURAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_20 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_20;

architecture SYN_STRUCTURAL of PG_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n9, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_18_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_18_1;

architecture SYN_STRUCTURAL of PG_18_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n8, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_11 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_11;

architecture SYN_STRUCTURAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_23 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_23;

architecture SYN_STRUCTURAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_21_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_21_1;

architecture SYN_STRUCTURAL of PG_21_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_22_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_22_1;

architecture SYN_STRUCTURAL of PG_22_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_12 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_12;

architecture SYN_STRUCTURAL of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_24_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_24_1;

architecture SYN_STRUCTURAL of PG_24_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n6);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_25_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_25_1;

architecture SYN_STRUCTURAL of PG_25_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_26_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_26_1;

architecture SYN_STRUCTURAL of PG_26_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_0_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_0_1;

architecture SYN_STRUCTURAL of PG_0_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_2 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_2;

architecture SYN_STRUCTURAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_1;

architecture SYN_STRUCTURAL of PGnet_block_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_2 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_2;

architecture SYN_STRUCTURAL of PGnet_block_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_3 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_3;

architecture SYN_STRUCTURAL of PGnet_block_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_4 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_4;

architecture SYN_STRUCTURAL of PGnet_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_5 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_5;

architecture SYN_STRUCTURAL of PGnet_block_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_6 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_6;

architecture SYN_STRUCTURAL of PGnet_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_7 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_7;

architecture SYN_STRUCTURAL of PGnet_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_8 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_8;

architecture SYN_STRUCTURAL of PGnet_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_9 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_9;

architecture SYN_STRUCTURAL of PGnet_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_10 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_10;

architecture SYN_STRUCTURAL of PGnet_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_11 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_11;

architecture SYN_STRUCTURAL of PGnet_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_12 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_12;

architecture SYN_STRUCTURAL of PGnet_block_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_13 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_13;

architecture SYN_STRUCTURAL of PGnet_block_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_14 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_14;

architecture SYN_STRUCTURAL of PGnet_block_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_15 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_15;

architecture SYN_STRUCTURAL of PGnet_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_16 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_16;

architecture SYN_STRUCTURAL of PGnet_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_17 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_17;

architecture SYN_STRUCTURAL of PGnet_block_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_18 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_18;

architecture SYN_STRUCTURAL of PGnet_block_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_19 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_19;

architecture SYN_STRUCTURAL of PGnet_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_20 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_20;

architecture SYN_STRUCTURAL of PGnet_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_21 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_21;

architecture SYN_STRUCTURAL of PGnet_block_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_22 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_22;

architecture SYN_STRUCTURAL of PGnet_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_23 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_23;

architecture SYN_STRUCTURAL of PGnet_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_24 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_24;

architecture SYN_STRUCTURAL of PGnet_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_25 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_25;

architecture SYN_STRUCTURAL of PGnet_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_26 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_26;

architecture SYN_STRUCTURAL of PGnet_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_27 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_27;

architecture SYN_STRUCTURAL of PGnet_block_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_28 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_28;

architecture SYN_STRUCTURAL of PGnet_block_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_29 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_29;

architecture SYN_STRUCTURAL of PGnet_block_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_30_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_30_1;

architecture SYN_STRUCTURAL of PGnet_block_30_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_31_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_31_1;

architecture SYN_STRUCTURAL of PGnet_block_31_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_0_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_0_1;

architecture SYN_STRUCTURAL of G_0_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_0_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_0_1;

architecture SYN_STRUCTURAL of PGnet_block_0_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_8;

architecture SYN_STRUCTURAL of carry_select_N4_8 is

   component MUX21_GENERIC_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_8 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_9;

architecture SYN_STRUCTURAL of carry_select_N4_9 is

   component MUX21_GENERIC_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_9 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_10;

architecture SYN_STRUCTURAL of carry_select_N4_10 is

   component MUX21_GENERIC_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_10 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_11;

architecture SYN_STRUCTURAL of carry_select_N4_11 is

   component MUX21_GENERIC_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_11 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_12;

architecture SYN_STRUCTURAL of carry_select_N4_12 is

   component MUX21_GENERIC_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_12 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_6_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_6_0;

architecture SYN_STRUCTURAL of carry_select_N4_6_0 is

   component MUX21_GENERIC_N4_6_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_6_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_7_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_7_0;

architecture SYN_STRUCTURAL of carry_select_N4_7_0 is

   component MUX21_GENERIC_N4_7_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_14_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_14_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_7_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_0_0;

architecture SYN_STRUCTURAL of carry_select_N4_0_0 is

   component MUX21_GENERIC_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_15_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_15_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_0_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_10 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_10;

architecture SYN_STRUCTURAL of G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_11 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_11;

architecture SYN_STRUCTURAL of G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_12 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_12;

architecture SYN_STRUCTURAL of G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_13 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_13;

architecture SYN_STRUCTURAL of G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_27 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_27;

architecture SYN_STRUCTURAL of PG_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_28 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_28;

architecture SYN_STRUCTURAL of PG_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_5_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_5_0;

architecture SYN_STRUCTURAL of G_5_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_6_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_6_0;

architecture SYN_STRUCTURAL of G_6_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_29 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_29;

architecture SYN_STRUCTURAL of PG_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_4_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_4_0;

architecture SYN_STRUCTURAL of PG_4_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_30 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_30;

architecture SYN_STRUCTURAL of PG_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_14 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_14;

architecture SYN_STRUCTURAL of G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_31 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_31;

architecture SYN_STRUCTURAL of PG_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_32 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_32;

architecture SYN_STRUCTURAL of PG_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_33 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_33;

architecture SYN_STRUCTURAL of PG_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_34 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_34;

architecture SYN_STRUCTURAL of PG_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_35 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_35;

architecture SYN_STRUCTURAL of PG_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_36 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_36;

architecture SYN_STRUCTURAL of PG_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_37 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_37;

architecture SYN_STRUCTURAL of PG_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_8_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_8_0;

architecture SYN_STRUCTURAL of G_8_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_38 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_38;

architecture SYN_STRUCTURAL of PG_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_39 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_39;

architecture SYN_STRUCTURAL of PG_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_40 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_40;

architecture SYN_STRUCTURAL of PG_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_41 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_41;

architecture SYN_STRUCTURAL of PG_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_42 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_42;

architecture SYN_STRUCTURAL of PG_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_18_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_18_0;

architecture SYN_STRUCTURAL of PG_18_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_43 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_43;

architecture SYN_STRUCTURAL of PG_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_44 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_44;

architecture SYN_STRUCTURAL of PG_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_21_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_21_0;

architecture SYN_STRUCTURAL of PG_21_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_22_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_22_0;

architecture SYN_STRUCTURAL of PG_22_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_45 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_45;

architecture SYN_STRUCTURAL of PG_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_24_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_24_0;

architecture SYN_STRUCTURAL of PG_24_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_25_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_25_0;

architecture SYN_STRUCTURAL of PG_25_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_26_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_26_0;

architecture SYN_STRUCTURAL of PG_26_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG_0_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_0_0;

architecture SYN_STRUCTURAL of PG_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_15 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_15;

architecture SYN_STRUCTURAL of G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_32 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_32;

architecture SYN_STRUCTURAL of PGnet_block_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_33 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_33;

architecture SYN_STRUCTURAL of PGnet_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_34 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_34;

architecture SYN_STRUCTURAL of PGnet_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_35 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_35;

architecture SYN_STRUCTURAL of PGnet_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_36 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_36;

architecture SYN_STRUCTURAL of PGnet_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_37 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_37;

architecture SYN_STRUCTURAL of PGnet_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_38 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_38;

architecture SYN_STRUCTURAL of PGnet_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_39 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_39;

architecture SYN_STRUCTURAL of PGnet_block_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_40 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_40;

architecture SYN_STRUCTURAL of PGnet_block_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_41 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_41;

architecture SYN_STRUCTURAL of PGnet_block_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_42 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_42;

architecture SYN_STRUCTURAL of PGnet_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_43 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_43;

architecture SYN_STRUCTURAL of PGnet_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_44 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_44;

architecture SYN_STRUCTURAL of PGnet_block_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_45 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_45;

architecture SYN_STRUCTURAL of PGnet_block_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_46 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_46;

architecture SYN_STRUCTURAL of PGnet_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_47 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_47;

architecture SYN_STRUCTURAL of PGnet_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_48 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_48;

architecture SYN_STRUCTURAL of PGnet_block_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_49 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_49;

architecture SYN_STRUCTURAL of PGnet_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_50 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_50;

architecture SYN_STRUCTURAL of PGnet_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_51 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_51;

architecture SYN_STRUCTURAL of PGnet_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_52 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_52;

architecture SYN_STRUCTURAL of PGnet_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_53 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_53;

architecture SYN_STRUCTURAL of PGnet_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_54 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_54;

architecture SYN_STRUCTURAL of PGnet_block_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_55 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_55;

architecture SYN_STRUCTURAL of PGnet_block_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_56 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_56;

architecture SYN_STRUCTURAL of PGnet_block_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_57 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_57;

architecture SYN_STRUCTURAL of PGnet_block_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_58 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_58;

architecture SYN_STRUCTURAL of PGnet_block_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_59 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_59;

architecture SYN_STRUCTURAL of PGnet_block_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_60 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_60;

architecture SYN_STRUCTURAL of PGnet_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_30_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_30_0;

architecture SYN_STRUCTURAL of PGnet_block_30_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_31_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_31_0;

architecture SYN_STRUCTURAL of PGnet_block_31_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G_0_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_0_0;

architecture SYN_STRUCTURAL of G_0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block_0_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_0_0;

architecture SYN_STRUCTURAL of PGnet_block_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4;

architecture SYN_struct of MUX21_GENERIC_N4 is

   component MUX21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity rca_generic_N4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4;

architecture SYN_STRUCTURAL of rca_generic_N4 is

   component FA
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), Co 
                           => CTMP_2_port);
   FAI_3 : FA port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), Co 
                           => CTMP_3_port);
   FAI_4 : FA port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), Co 
                           => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity sum_generator_Nbits32_Nblocks8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Carry : in std_logic_vector
         (8 downto 0);  S : out std_logic_vector (31 downto 0);  Cout : out 
         std_logic);

end sum_generator_Nbits32_Nblocks8_1;

architecture SYN_STRUCTURAL of sum_generator_Nbits32_Nblocks8_1 is

   component carry_select_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(8);
   
   CS_0 : carry_select_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Carry(0), S(3) => S(3),
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4_7_1 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Carry(1), S(3) => S(7),
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4_6_1 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Carry(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Carry(3), S(3) 
                           => S(15), S(2) => S(14), S(1) => S(13), S(0) => 
                           S(12));
   CS_4 : carry_select_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Carry(4), S(3) 
                           => S(19), S(2) => S(18), S(1) => S(17), S(0) => 
                           S(16));
   CS_5 : carry_select_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Carry(5), S(3) 
                           => S(23), S(2) => S(22), S(1) => S(21), S(0) => 
                           S(20));
   CS_6 : carry_select_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Carry(6), S(3) 
                           => S(27), S(2) => S(26), S(1) => S(25), S(0) => 
                           S(24));
   CS_7 : carry_select_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Carry(7), S(3) 
                           => S(31), S(2) => S(30), S(1) => S(29), S(0) => 
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_generator_N32_Nblocks8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_Nblocks8_1;

architecture SYN_STRUCTURAL of carry_generator_N32_Nblocks8_1 is

   component G_3
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_4
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_7
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_9
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_2
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_5_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_6_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_3
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_4_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_13
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_5
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_6
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_14
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_15
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_16
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_17
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_19
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_8_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_7
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_8
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_9
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_10
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_20
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_18_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_11
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_23
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_21_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_22_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_12
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_24_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_25_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_26_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_0_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_2
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_2
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_3
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_4
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_5
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_6
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_7
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_8
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_9
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_10
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_11
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_12
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_13
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_14
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_15
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_16
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_17
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_18
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_19
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_20
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_21
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_22
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_23
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_24
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_25
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_26
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_27
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_28
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_29
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_30_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_31_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_0_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_0_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   signal Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_3_port, 
      g_cin, p_cin, Gsignal_1_31_port, Gsignal_1_30_port, Gsignal_1_29_port, 
      Gsignal_1_28_port, Gsignal_1_27_port, Gsignal_1_26_port, 
      Gsignal_1_25_port, Gsignal_1_24_port, Gsignal_1_23_port, 
      Gsignal_1_22_port, Gsignal_1_21_port, Gsignal_1_20_port, 
      Gsignal_1_19_port, Gsignal_1_18_port, Gsignal_1_17_port, 
      Gsignal_1_16_port, Gsignal_1_15_port, Gsignal_1_14_port, 
      Gsignal_1_13_port, Gsignal_1_12_port, Gsignal_1_11_port, 
      Gsignal_1_10_port, Gsignal_1_9_port, Gsignal_1_8_port, Gsignal_1_7_port, 
      Gsignal_1_6_port, Gsignal_1_5_port, Gsignal_1_4_port, Gsignal_1_3_port, 
      Gsignal_1_2_port, Gsignal_1_1_port, Gsignal_1_0_port, Gsignal_2_31_port, 
      Gsignal_2_29_port, Gsignal_2_27_port, Gsignal_2_25_port, 
      Gsignal_2_23_port, Gsignal_2_21_port, Gsignal_2_19_port, 
      Gsignal_2_17_port, Gsignal_2_15_port, Gsignal_2_13_port, 
      Gsignal_2_11_port, Gsignal_2_9_port, Gsignal_2_7_port, Gsignal_2_5_port, 
      Gsignal_2_3_port, Gsignal_2_1_port, Gsignal_3_31_port, Gsignal_3_23_port,
      Gsignal_3_15_port, Gsignal_3_7_port, Gsignal_4_31_port, Gsignal_4_15_port
      , Gsignal_5_31_port, Gsignal_5_27_port, Psignal_1_31_port, 
      Psignal_1_30_port, Psignal_1_29_port, Psignal_1_28_port, 
      Psignal_1_27_port, Psignal_1_26_port, Psignal_1_25_port, 
      Psignal_1_24_port, Psignal_1_23_port, Psignal_1_22_port, 
      Psignal_1_21_port, Psignal_1_20_port, Psignal_1_19_port, 
      Psignal_1_18_port, Psignal_1_17_port, Psignal_1_16_port, 
      Psignal_1_15_port, Psignal_1_14_port, Psignal_1_13_port, 
      Psignal_1_12_port, Psignal_1_11_port, Psignal_1_10_port, Psignal_1_9_port
      , Psignal_1_8_port, Psignal_1_7_port, Psignal_1_6_port, Psignal_1_5_port,
      Psignal_1_4_port, Psignal_1_3_port, Psignal_1_2_port, Psignal_1_1_port, 
      Psignal_2_31_port, Psignal_2_29_port, Psignal_2_27_port, 
      Psignal_2_25_port, Psignal_2_23_port, Psignal_2_21_port, 
      Psignal_2_19_port, Psignal_2_17_port, Psignal_2_15_port, 
      Psignal_2_13_port, Psignal_2_11_port, Psignal_2_9_port, Psignal_2_7_port,
      Psignal_2_5_port, Psignal_2_3_port, Psignal_3_31_port, Psignal_3_27_port,
      Psignal_3_23_port, Psignal_3_19_port, Psignal_3_15_port, Psignal_3_7_port
      , Psignal_4_31_port, Psignal_4_23_port, Psignal_4_15_port, 
      Psignal_5_31_port, Psignal_5_27_port, n8, Cout_1_port, n10, Cout_2_port, 
      n12, n13, n15, Cout_4_port : std_logic;

begin
   Cout <= ( Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, Ci );
   
   PGnet_Cin_0 : PGnet_block_0_1 port map( A => A(0), B => B(0), pout => p_cin,
                           gout => g_cin);
   GCin_0 : G_0_1 port map( gleft => g_cin, gright => Ci, pleft => p_cin, gout 
                           => Gsignal_1_0_port);
   PGnet_1 : PGnet_block_31_1 port map( A => A(1), B => B(1), pout => 
                           Psignal_1_1_port, gout => Gsignal_1_1_port);
   PGnet_2 : PGnet_block_30_1 port map( A => A(2), B => B(2), pout => 
                           Psignal_1_2_port, gout => Gsignal_1_2_port);
   PGnet_3 : PGnet_block_29 port map( A => A(3), B => B(3), pout => 
                           Psignal_1_3_port, gout => Gsignal_1_3_port);
   PGnet_4 : PGnet_block_28 port map( A => A(4), B => B(4), pout => 
                           Psignal_1_4_port, gout => Gsignal_1_4_port);
   PGnet_5 : PGnet_block_27 port map( A => A(5), B => B(5), pout => 
                           Psignal_1_5_port, gout => Gsignal_1_5_port);
   PGnet_6 : PGnet_block_26 port map( A => A(6), B => B(6), pout => 
                           Psignal_1_6_port, gout => Gsignal_1_6_port);
   PGnet_7 : PGnet_block_25 port map( A => A(7), B => B(7), pout => 
                           Psignal_1_7_port, gout => Gsignal_1_7_port);
   PGnet_8 : PGnet_block_24 port map( A => A(8), B => B(8), pout => 
                           Psignal_1_8_port, gout => Gsignal_1_8_port);
   PGnet_9 : PGnet_block_23 port map( A => A(9), B => B(9), pout => 
                           Psignal_1_9_port, gout => Gsignal_1_9_port);
   PGnet_10 : PGnet_block_22 port map( A => A(10), B => B(10), pout => 
                           Psignal_1_10_port, gout => Gsignal_1_10_port);
   PGnet_11 : PGnet_block_21 port map( A => A(11), B => B(11), pout => 
                           Psignal_1_11_port, gout => Gsignal_1_11_port);
   PGnet_12 : PGnet_block_20 port map( A => A(12), B => B(12), pout => 
                           Psignal_1_12_port, gout => Gsignal_1_12_port);
   PGnet_13 : PGnet_block_19 port map( A => A(13), B => B(13), pout => 
                           Psignal_1_13_port, gout => Gsignal_1_13_port);
   PGnet_14 : PGnet_block_18 port map( A => A(14), B => B(14), pout => 
                           Psignal_1_14_port, gout => Gsignal_1_14_port);
   PGnet_15 : PGnet_block_17 port map( A => A(15), B => B(15), pout => 
                           Psignal_1_15_port, gout => Gsignal_1_15_port);
   PGnet_16 : PGnet_block_16 port map( A => A(16), B => B(16), pout => 
                           Psignal_1_16_port, gout => Gsignal_1_16_port);
   PGnet_17 : PGnet_block_15 port map( A => A(17), B => B(17), pout => 
                           Psignal_1_17_port, gout => Gsignal_1_17_port);
   PGnet_18 : PGnet_block_14 port map( A => A(18), B => B(18), pout => 
                           Psignal_1_18_port, gout => Gsignal_1_18_port);
   PGnet_19 : PGnet_block_13 port map( A => A(19), B => B(19), pout => 
                           Psignal_1_19_port, gout => Gsignal_1_19_port);
   PGnet_20 : PGnet_block_12 port map( A => A(20), B => B(20), pout => 
                           Psignal_1_20_port, gout => Gsignal_1_20_port);
   PGnet_21 : PGnet_block_11 port map( A => A(21), B => B(21), pout => 
                           Psignal_1_21_port, gout => Gsignal_1_21_port);
   PGnet_22 : PGnet_block_10 port map( A => A(22), B => B(22), pout => 
                           Psignal_1_22_port, gout => Gsignal_1_22_port);
   PGnet_23 : PGnet_block_9 port map( A => A(23), B => B(23), pout => 
                           Psignal_1_23_port, gout => Gsignal_1_23_port);
   PGnet_24 : PGnet_block_8 port map( A => A(24), B => B(24), pout => 
                           Psignal_1_24_port, gout => Gsignal_1_24_port);
   PGnet_25 : PGnet_block_7 port map( A => A(25), B => B(25), pout => 
                           Psignal_1_25_port, gout => Gsignal_1_25_port);
   PGnet_26 : PGnet_block_6 port map( A => A(26), B => B(26), pout => 
                           Psignal_1_26_port, gout => Gsignal_1_26_port);
   PGnet_27 : PGnet_block_5 port map( A => A(27), B => B(27), pout => 
                           Psignal_1_27_port, gout => Gsignal_1_27_port);
   PGnet_28 : PGnet_block_4 port map( A => A(28), B => B(28), pout => 
                           Psignal_1_28_port, gout => Gsignal_1_28_port);
   PGnet_29 : PGnet_block_3 port map( A => A(29), B => B(29), pout => 
                           Psignal_1_29_port, gout => Gsignal_1_29_port);
   PGnet_30 : PGnet_block_2 port map( A => A(30), B => B(30), pout => 
                           Psignal_1_30_port, gout => Gsignal_1_30_port);
   PGnet_31 : PGnet_block_1 port map( A => A(31), B => B(31), pout => 
                           Psignal_1_31_port, gout => Gsignal_1_31_port);
   Gblock_1_1 : G_2 port map( gleft => Gsignal_1_1_port, gright => 
                           Gsignal_1_0_port, pleft => Psignal_1_1_port, gout =>
                           Gsignal_2_1_port);
   PGblock_1_3 : PG_0_1 port map( gleft => Gsignal_1_3_port, gright => 
                           Gsignal_1_2_port, pleft => Psignal_1_3_port, pright 
                           => Psignal_1_2_port, pout => Psignal_2_3_port, gout 
                           => Gsignal_2_3_port);
   PGblock_1_5 : PG_26_1 port map( gleft => Gsignal_1_5_port, gright => 
                           Gsignal_1_4_port, pleft => Psignal_1_5_port, pright 
                           => Psignal_1_4_port, pout => Psignal_2_5_port, gout 
                           => Gsignal_2_5_port);
   PGblock_1_7 : PG_25_1 port map( gleft => Gsignal_1_7_port, gright => 
                           Gsignal_1_6_port, pleft => Psignal_1_7_port, pright 
                           => Psignal_1_6_port, pout => Psignal_2_7_port, gout 
                           => Gsignal_2_7_port);
   PGblock_1_9 : PG_24_1 port map( gleft => Gsignal_1_9_port, gright => 
                           Gsignal_1_8_port, pleft => Psignal_1_9_port, pright 
                           => Psignal_1_8_port, pout => Psignal_2_9_port, gout 
                           => Gsignal_2_9_port);
   PGblock_1_11 : PG_12 port map( gleft => Gsignal_1_11_port, gright => 
                           Gsignal_1_10_port, pleft => Psignal_1_11_port, 
                           pright => Psignal_1_10_port, pout => 
                           Psignal_2_11_port, gout => Gsignal_2_11_port);
   PGblock_1_13 : PG_22_1 port map( gleft => Gsignal_1_13_port, gright => 
                           Gsignal_1_12_port, pleft => Psignal_1_13_port, 
                           pright => Psignal_1_12_port, pout => 
                           Psignal_2_13_port, gout => Gsignal_2_13_port);
   PGblock_1_15 : PG_21_1 port map( gleft => Gsignal_1_15_port, gright => 
                           Gsignal_1_14_port, pleft => Psignal_1_15_port, 
                           pright => Psignal_1_14_port, pout => 
                           Psignal_2_15_port, gout => Gsignal_2_15_port);
   PGblock_1_17 : PG_23 port map( gleft => Gsignal_1_17_port, gright => 
                           Gsignal_1_16_port, pleft => Psignal_1_17_port, 
                           pright => Psignal_1_16_port, pout => 
                           Psignal_2_17_port, gout => Gsignal_2_17_port);
   PGblock_1_19 : PG_11 port map( gleft => Gsignal_1_19_port, gright => 
                           Gsignal_1_18_port, pleft => Psignal_1_19_port, 
                           pright => Psignal_1_18_port, pout => 
                           Psignal_2_19_port, gout => Gsignal_2_19_port);
   PGblock_1_21 : PG_18_1 port map( gleft => Gsignal_1_21_port, gright => 
                           Gsignal_1_20_port, pleft => Psignal_1_21_port, 
                           pright => Psignal_1_20_port, pout => 
                           Psignal_2_21_port, gout => Gsignal_2_21_port);
   PGblock_1_23 : PG_20 port map( gleft => Gsignal_1_23_port, gright => 
                           Gsignal_1_22_port, pleft => Psignal_1_23_port, 
                           pright => Psignal_1_22_port, pout => 
                           Psignal_2_23_port, gout => Gsignal_2_23_port);
   PGblock_1_25 : PG_10 port map( gleft => Gsignal_1_25_port, gright => 
                           Gsignal_1_24_port, pleft => Psignal_1_25_port, 
                           pright => Psignal_1_24_port, pout => 
                           Psignal_2_25_port, gout => Gsignal_2_25_port);
   PGblock_1_27 : PG_9 port map( gleft => Gsignal_1_27_port, gright => 
                           Gsignal_1_26_port, pleft => Psignal_1_27_port, 
                           pright => Psignal_1_26_port, pout => 
                           Psignal_2_27_port, gout => Gsignal_2_27_port);
   PGblock_1_29 : PG_8 port map( gleft => Gsignal_1_29_port, gright => 
                           Gsignal_1_28_port, pleft => Psignal_1_29_port, 
                           pright => Psignal_1_28_port, pout => 
                           Psignal_2_29_port, gout => Gsignal_2_29_port);
   PGblock_1_31 : PG_7 port map( gleft => Gsignal_1_31_port, gright => 
                           Gsignal_1_30_port, pleft => Psignal_1_31_port, 
                           pright => Psignal_1_30_port, pout => 
                           Psignal_2_31_port, gout => Gsignal_2_31_port);
   Gblock_2_3 : G_8_1 port map( gleft => Gsignal_2_3_port, gright => 
                           Gsignal_2_1_port, pleft => Psignal_2_3_port, gout =>
                           Cout_1_port);
   PGblock_2_7 : PG_19 port map( gleft => Gsignal_2_7_port, gright => 
                           Gsignal_2_5_port, pleft => Psignal_2_7_port, pright 
                           => Psignal_2_5_port, pout => Psignal_3_7_port, gout 
                           => Gsignal_3_7_port);
   PGblock_2_11 : PG_17 port map( gleft => Gsignal_2_11_port, gright => 
                           Gsignal_2_9_port, pleft => Psignal_2_11_port, pright
                           => Psignal_2_9_port, pout => n8, gout => n10);
   PGblock_2_15 : PG_16 port map( gleft => Gsignal_2_15_port, gright => 
                           Gsignal_2_13_port, pleft => Psignal_2_15_port, 
                           pright => Psignal_2_13_port, pout => 
                           Psignal_3_15_port, gout => Gsignal_3_15_port);
   PGblock_2_19 : PG_15 port map( gleft => Gsignal_2_19_port, gright => 
                           Gsignal_2_17_port, pleft => Psignal_2_19_port, 
                           pright => Psignal_2_17_port, pout => 
                           Psignal_3_19_port, gout => n13);
   PGblock_2_23 : PG_14 port map( gleft => Gsignal_2_23_port, gright => 
                           Gsignal_2_21_port, pleft => Psignal_2_23_port, 
                           pright => Psignal_2_21_port, pout => 
                           Psignal_3_23_port, gout => Gsignal_3_23_port);
   PGblock_2_27 : PG_6 port map( gleft => Gsignal_2_27_port, gright => 
                           Gsignal_2_25_port, pleft => Psignal_2_27_port, 
                           pright => Psignal_2_25_port, pout => 
                           Psignal_3_27_port, gout => n12);
   PGblock_2_31 : PG_5 port map( gleft => Gsignal_2_31_port, gright => 
                           Gsignal_2_29_port, pleft => Psignal_2_31_port, 
                           pright => Psignal_2_29_port, pout => 
                           Psignal_3_31_port, gout => Gsignal_3_31_port);
   Gblock_3_7 : G_1 port map( gleft => Gsignal_3_7_port, gright => Cout_1_port,
                           pleft => Psignal_3_7_port, gout => Cout_2_port);
   PGblock_3_15 : PG_13 port map( gleft => Gsignal_3_15_port, gright => n10, 
                           pleft => Psignal_3_15_port, pright => n8, pout => 
                           Psignal_4_15_port, gout => Gsignal_4_15_port);
   PGblock_3_23 : PG_4_1 port map( gleft => Gsignal_3_23_port, gright => n13, 
                           pleft => Psignal_3_23_port, pright => 
                           Psignal_3_19_port, pout => Psignal_4_23_port, gout 
                           => n15);
   PGblock_3_31 : PG_3 port map( gleft => Gsignal_3_31_port, gright => n12, 
                           pleft => Psignal_3_31_port, pright => 
                           Psignal_3_27_port, pout => Psignal_4_31_port, gout 
                           => Gsignal_4_31_port);
   Gblock_4_11 : G_6_1 port map( gleft => n10, gright => Cout_2_port, pleft => 
                           n8, gout => Cout_3_port);
   Gblock_4_15 : G_5_1 port map( gleft => Gsignal_4_15_port, gright => 
                           Cout_2_port, pleft => Psignal_4_15_port, gout => 
                           Cout_4_port);
   PGblock_4_27 : PG_1 port map( gleft => n12, gright => n15, pleft => 
                           Psignal_3_27_port, pright => Psignal_4_23_port, pout
                           => Psignal_5_27_port, gout => Gsignal_5_27_port);
   PGblock_4_31 : PG_2 port map( gleft => Gsignal_4_31_port, gright => n15, 
                           pleft => Psignal_4_31_port, pright => 
                           Psignal_4_23_port, pout => Psignal_5_31_port, gout 
                           => Gsignal_5_31_port);
   Gblock_5_19 : G_9 port map( gleft => n13, gright => Cout_4_port, pleft => 
                           Psignal_3_19_port, gout => Cout_5_port);
   Gblock_5_23 : G_7 port map( gleft => n15, gright => Cout_4_port, pleft => 
                           Psignal_4_23_port, gout => Cout_6_port);
   Gblock_5_27 : G_4 port map( gleft => Gsignal_5_27_port, gright => 
                           Cout_4_port, pleft => Psignal_5_27_port, gout => 
                           Cout_7_port);
   Gblock_5_31 : G_3 port map( gleft => Gsignal_5_31_port, gright => 
                           Cout_4_port, pleft => Psignal_5_31_port, gout => 
                           Cout_8_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => A, A2 => B, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity sum_generator_Nbits32_Nblocks8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Carry : in std_logic_vector
         (8 downto 0);  S : out std_logic_vector (31 downto 0);  Cout : out 
         std_logic);

end sum_generator_Nbits32_Nblocks8_0;

architecture SYN_STRUCTURAL of sum_generator_Nbits32_Nblocks8_0 is

   component carry_select_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(8);
   
   CS_0 : carry_select_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Carry(0), S(3) => S(3),
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4_7_0 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Carry(1), S(3) => S(7),
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4_6_0 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Carry(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4_12 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Carry(3), S(3) 
                           => S(15), S(2) => S(14), S(1) => S(13), S(0) => 
                           S(12));
   CS_4 : carry_select_N4_11 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Carry(4), S(3) 
                           => S(19), S(2) => S(18), S(1) => S(17), S(0) => 
                           S(16));
   CS_5 : carry_select_N4_10 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Carry(5), S(3) 
                           => S(23), S(2) => S(22), S(1) => S(21), S(0) => 
                           S(20));
   CS_6 : carry_select_N4_9 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Carry(6), S(3) 
                           => S(27), S(2) => S(26), S(1) => S(25), S(0) => 
                           S(24));
   CS_7 : carry_select_N4_8 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Carry(7), S(3) 
                           => S(31), S(2) => S(30), S(1) => S(29), S(0) => 
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_generator_N32_Nblocks8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_Nblocks8_0;

architecture SYN_STRUCTURAL of carry_generator_N32_Nblocks8_0 is

   component G_10
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_11
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_12
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_13
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_27
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_28
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_5_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_6_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_29
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_4_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_30
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_14
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_31
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_32
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_33
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_34
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_35
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_36
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_37
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_8_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_38
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_39
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_40
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_41
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_42
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_18_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_43
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_44
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_21_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_22_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_45
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_24_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_25_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_26_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_0_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_15
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_32
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_33
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_34
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_35
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_36
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_37
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_38
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_39
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_40
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_41
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_42
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_43
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_44
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_45
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_46
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_47
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_48
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_49
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_50
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_51
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_52
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_53
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_54
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_55
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_56
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_57
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_58
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_59
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_60
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_30_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_31_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_0_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_0_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   signal Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_3_port, 
      g_cin, p_cin, Gsignal_1_31_port, Gsignal_1_30_port, Gsignal_1_29_port, 
      Gsignal_1_28_port, Gsignal_1_27_port, Gsignal_1_26_port, 
      Gsignal_1_25_port, Gsignal_1_24_port, Gsignal_1_23_port, 
      Gsignal_1_22_port, Gsignal_1_21_port, Gsignal_1_20_port, 
      Gsignal_1_19_port, Gsignal_1_18_port, Gsignal_1_17_port, 
      Gsignal_1_16_port, Gsignal_1_15_port, Gsignal_1_14_port, 
      Gsignal_1_13_port, Gsignal_1_12_port, Gsignal_1_11_port, 
      Gsignal_1_10_port, Gsignal_1_9_port, Gsignal_1_8_port, Gsignal_1_7_port, 
      Gsignal_1_6_port, Gsignal_1_5_port, Gsignal_1_4_port, Gsignal_1_3_port, 
      Gsignal_1_2_port, Gsignal_1_1_port, Gsignal_1_0_port, Gsignal_2_31_port, 
      Gsignal_2_29_port, Gsignal_2_27_port, Gsignal_2_25_port, 
      Gsignal_2_23_port, Gsignal_2_21_port, Gsignal_2_19_port, 
      Gsignal_2_17_port, Gsignal_2_15_port, Gsignal_2_13_port, 
      Gsignal_2_11_port, Gsignal_2_9_port, Gsignal_2_7_port, Gsignal_2_5_port, 
      Gsignal_2_3_port, Gsignal_2_1_port, Gsignal_3_31_port, Gsignal_3_23_port,
      Gsignal_3_15_port, Gsignal_3_7_port, Gsignal_4_31_port, Gsignal_4_15_port
      , Gsignal_5_31_port, Gsignal_5_27_port, Psignal_1_31_port, 
      Psignal_1_30_port, Psignal_1_29_port, Psignal_1_28_port, 
      Psignal_1_27_port, Psignal_1_26_port, Psignal_1_25_port, 
      Psignal_1_24_port, Psignal_1_23_port, Psignal_1_22_port, 
      Psignal_1_21_port, Psignal_1_20_port, Psignal_1_19_port, 
      Psignal_1_18_port, Psignal_1_17_port, Psignal_1_16_port, 
      Psignal_1_15_port, Psignal_1_14_port, Psignal_1_13_port, 
      Psignal_1_12_port, Psignal_1_11_port, Psignal_1_10_port, Psignal_1_9_port
      , Psignal_1_8_port, Psignal_1_7_port, Psignal_1_6_port, Psignal_1_5_port,
      Psignal_1_4_port, Psignal_1_3_port, Psignal_1_2_port, Psignal_1_1_port, 
      Psignal_2_31_port, Psignal_2_29_port, Psignal_2_27_port, 
      Psignal_2_25_port, Psignal_2_23_port, Psignal_2_21_port, 
      Psignal_2_19_port, Psignal_2_17_port, Psignal_2_15_port, 
      Psignal_2_13_port, Psignal_2_11_port, Psignal_2_9_port, Psignal_2_7_port,
      Psignal_2_5_port, Psignal_2_3_port, Psignal_3_31_port, Psignal_3_27_port,
      Psignal_3_23_port, Psignal_3_19_port, Psignal_3_15_port, Psignal_3_7_port
      , Psignal_4_31_port, Psignal_4_23_port, Psignal_4_15_port, 
      Psignal_5_31_port, Psignal_5_27_port, n8, Cout_1_port, n10, Cout_2_port, 
      n12, n13, n15, Cout_4_port : std_logic;

begin
   Cout <= ( Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, Ci );
   
   PGnet_Cin_0 : PGnet_block_0_0 port map( A => A(0), B => B(0), pout => p_cin,
                           gout => g_cin);
   GCin_0 : G_0_0 port map( gleft => g_cin, gright => Ci, pleft => p_cin, gout 
                           => Gsignal_1_0_port);
   PGnet_1 : PGnet_block_31_0 port map( A => A(1), B => B(1), pout => 
                           Psignal_1_1_port, gout => Gsignal_1_1_port);
   PGnet_2 : PGnet_block_30_0 port map( A => A(2), B => B(2), pout => 
                           Psignal_1_2_port, gout => Gsignal_1_2_port);
   PGnet_3 : PGnet_block_60 port map( A => A(3), B => B(3), pout => 
                           Psignal_1_3_port, gout => Gsignal_1_3_port);
   PGnet_4 : PGnet_block_59 port map( A => A(4), B => B(4), pout => 
                           Psignal_1_4_port, gout => Gsignal_1_4_port);
   PGnet_5 : PGnet_block_58 port map( A => A(5), B => B(5), pout => 
                           Psignal_1_5_port, gout => Gsignal_1_5_port);
   PGnet_6 : PGnet_block_57 port map( A => A(6), B => B(6), pout => 
                           Psignal_1_6_port, gout => Gsignal_1_6_port);
   PGnet_7 : PGnet_block_56 port map( A => A(7), B => B(7), pout => 
                           Psignal_1_7_port, gout => Gsignal_1_7_port);
   PGnet_8 : PGnet_block_55 port map( A => A(8), B => B(8), pout => 
                           Psignal_1_8_port, gout => Gsignal_1_8_port);
   PGnet_9 : PGnet_block_54 port map( A => A(9), B => B(9), pout => 
                           Psignal_1_9_port, gout => Gsignal_1_9_port);
   PGnet_10 : PGnet_block_53 port map( A => A(10), B => B(10), pout => 
                           Psignal_1_10_port, gout => Gsignal_1_10_port);
   PGnet_11 : PGnet_block_52 port map( A => A(11), B => B(11), pout => 
                           Psignal_1_11_port, gout => Gsignal_1_11_port);
   PGnet_12 : PGnet_block_51 port map( A => A(12), B => B(12), pout => 
                           Psignal_1_12_port, gout => Gsignal_1_12_port);
   PGnet_13 : PGnet_block_50 port map( A => A(13), B => B(13), pout => 
                           Psignal_1_13_port, gout => Gsignal_1_13_port);
   PGnet_14 : PGnet_block_49 port map( A => A(14), B => B(14), pout => 
                           Psignal_1_14_port, gout => Gsignal_1_14_port);
   PGnet_15 : PGnet_block_48 port map( A => A(15), B => B(15), pout => 
                           Psignal_1_15_port, gout => Gsignal_1_15_port);
   PGnet_16 : PGnet_block_47 port map( A => A(16), B => B(16), pout => 
                           Psignal_1_16_port, gout => Gsignal_1_16_port);
   PGnet_17 : PGnet_block_46 port map( A => A(17), B => B(17), pout => 
                           Psignal_1_17_port, gout => Gsignal_1_17_port);
   PGnet_18 : PGnet_block_45 port map( A => A(18), B => B(18), pout => 
                           Psignal_1_18_port, gout => Gsignal_1_18_port);
   PGnet_19 : PGnet_block_44 port map( A => A(19), B => B(19), pout => 
                           Psignal_1_19_port, gout => Gsignal_1_19_port);
   PGnet_20 : PGnet_block_43 port map( A => A(20), B => B(20), pout => 
                           Psignal_1_20_port, gout => Gsignal_1_20_port);
   PGnet_21 : PGnet_block_42 port map( A => A(21), B => B(21), pout => 
                           Psignal_1_21_port, gout => Gsignal_1_21_port);
   PGnet_22 : PGnet_block_41 port map( A => A(22), B => B(22), pout => 
                           Psignal_1_22_port, gout => Gsignal_1_22_port);
   PGnet_23 : PGnet_block_40 port map( A => A(23), B => B(23), pout => 
                           Psignal_1_23_port, gout => Gsignal_1_23_port);
   PGnet_24 : PGnet_block_39 port map( A => A(24), B => B(24), pout => 
                           Psignal_1_24_port, gout => Gsignal_1_24_port);
   PGnet_25 : PGnet_block_38 port map( A => A(25), B => B(25), pout => 
                           Psignal_1_25_port, gout => Gsignal_1_25_port);
   PGnet_26 : PGnet_block_37 port map( A => A(26), B => B(26), pout => 
                           Psignal_1_26_port, gout => Gsignal_1_26_port);
   PGnet_27 : PGnet_block_36 port map( A => A(27), B => B(27), pout => 
                           Psignal_1_27_port, gout => Gsignal_1_27_port);
   PGnet_28 : PGnet_block_35 port map( A => A(28), B => B(28), pout => 
                           Psignal_1_28_port, gout => Gsignal_1_28_port);
   PGnet_29 : PGnet_block_34 port map( A => A(29), B => B(29), pout => 
                           Psignal_1_29_port, gout => Gsignal_1_29_port);
   PGnet_30 : PGnet_block_33 port map( A => A(30), B => B(30), pout => 
                           Psignal_1_30_port, gout => Gsignal_1_30_port);
   PGnet_31 : PGnet_block_32 port map( A => A(31), B => B(31), pout => 
                           Psignal_1_31_port, gout => Gsignal_1_31_port);
   Gblock_1_1 : G_15 port map( gleft => Gsignal_1_1_port, gright => 
                           Gsignal_1_0_port, pleft => Psignal_1_1_port, gout =>
                           Gsignal_2_1_port);
   PGblock_1_3 : PG_0_0 port map( gleft => Gsignal_1_3_port, gright => 
                           Gsignal_1_2_port, pleft => Psignal_1_3_port, pright 
                           => Psignal_1_2_port, pout => Psignal_2_3_port, gout 
                           => Gsignal_2_3_port);
   PGblock_1_5 : PG_26_0 port map( gleft => Gsignal_1_5_port, gright => 
                           Gsignal_1_4_port, pleft => Psignal_1_5_port, pright 
                           => Psignal_1_4_port, pout => Psignal_2_5_port, gout 
                           => Gsignal_2_5_port);
   PGblock_1_7 : PG_25_0 port map( gleft => Gsignal_1_7_port, gright => 
                           Gsignal_1_6_port, pleft => Psignal_1_7_port, pright 
                           => Psignal_1_6_port, pout => Psignal_2_7_port, gout 
                           => Gsignal_2_7_port);
   PGblock_1_9 : PG_24_0 port map( gleft => Gsignal_1_9_port, gright => 
                           Gsignal_1_8_port, pleft => Psignal_1_9_port, pright 
                           => Psignal_1_8_port, pout => Psignal_2_9_port, gout 
                           => Gsignal_2_9_port);
   PGblock_1_11 : PG_45 port map( gleft => Gsignal_1_11_port, gright => 
                           Gsignal_1_10_port, pleft => Psignal_1_11_port, 
                           pright => Psignal_1_10_port, pout => 
                           Psignal_2_11_port, gout => Gsignal_2_11_port);
   PGblock_1_13 : PG_22_0 port map( gleft => Gsignal_1_13_port, gright => 
                           Gsignal_1_12_port, pleft => Psignal_1_13_port, 
                           pright => Psignal_1_12_port, pout => 
                           Psignal_2_13_port, gout => Gsignal_2_13_port);
   PGblock_1_15 : PG_21_0 port map( gleft => Gsignal_1_15_port, gright => 
                           Gsignal_1_14_port, pleft => Psignal_1_15_port, 
                           pright => Psignal_1_14_port, pout => 
                           Psignal_2_15_port, gout => Gsignal_2_15_port);
   PGblock_1_17 : PG_44 port map( gleft => Gsignal_1_17_port, gright => 
                           Gsignal_1_16_port, pleft => Psignal_1_17_port, 
                           pright => Psignal_1_16_port, pout => 
                           Psignal_2_17_port, gout => Gsignal_2_17_port);
   PGblock_1_19 : PG_43 port map( gleft => Gsignal_1_19_port, gright => 
                           Gsignal_1_18_port, pleft => Psignal_1_19_port, 
                           pright => Psignal_1_18_port, pout => 
                           Psignal_2_19_port, gout => Gsignal_2_19_port);
   PGblock_1_21 : PG_18_0 port map( gleft => Gsignal_1_21_port, gright => 
                           Gsignal_1_20_port, pleft => Psignal_1_21_port, 
                           pright => Psignal_1_20_port, pout => 
                           Psignal_2_21_port, gout => Gsignal_2_21_port);
   PGblock_1_23 : PG_42 port map( gleft => Gsignal_1_23_port, gright => 
                           Gsignal_1_22_port, pleft => Psignal_1_23_port, 
                           pright => Psignal_1_22_port, pout => 
                           Psignal_2_23_port, gout => Gsignal_2_23_port);
   PGblock_1_25 : PG_41 port map( gleft => Gsignal_1_25_port, gright => 
                           Gsignal_1_24_port, pleft => Psignal_1_25_port, 
                           pright => Psignal_1_24_port, pout => 
                           Psignal_2_25_port, gout => Gsignal_2_25_port);
   PGblock_1_27 : PG_40 port map( gleft => Gsignal_1_27_port, gright => 
                           Gsignal_1_26_port, pleft => Psignal_1_27_port, 
                           pright => Psignal_1_26_port, pout => 
                           Psignal_2_27_port, gout => Gsignal_2_27_port);
   PGblock_1_29 : PG_39 port map( gleft => Gsignal_1_29_port, gright => 
                           Gsignal_1_28_port, pleft => Psignal_1_29_port, 
                           pright => Psignal_1_28_port, pout => 
                           Psignal_2_29_port, gout => Gsignal_2_29_port);
   PGblock_1_31 : PG_38 port map( gleft => Gsignal_1_31_port, gright => 
                           Gsignal_1_30_port, pleft => Psignal_1_31_port, 
                           pright => Psignal_1_30_port, pout => 
                           Psignal_2_31_port, gout => Gsignal_2_31_port);
   Gblock_2_3 : G_8_0 port map( gleft => Gsignal_2_3_port, gright => 
                           Gsignal_2_1_port, pleft => Psignal_2_3_port, gout =>
                           Cout_1_port);
   PGblock_2_7 : PG_37 port map( gleft => Gsignal_2_7_port, gright => 
                           Gsignal_2_5_port, pleft => Psignal_2_7_port, pright 
                           => Psignal_2_5_port, pout => Psignal_3_7_port, gout 
                           => Gsignal_3_7_port);
   PGblock_2_11 : PG_36 port map( gleft => Gsignal_2_11_port, gright => 
                           Gsignal_2_9_port, pleft => Psignal_2_11_port, pright
                           => Psignal_2_9_port, pout => n8, gout => n10);
   PGblock_2_15 : PG_35 port map( gleft => Gsignal_2_15_port, gright => 
                           Gsignal_2_13_port, pleft => Psignal_2_15_port, 
                           pright => Psignal_2_13_port, pout => 
                           Psignal_3_15_port, gout => Gsignal_3_15_port);
   PGblock_2_19 : PG_34 port map( gleft => Gsignal_2_19_port, gright => 
                           Gsignal_2_17_port, pleft => Psignal_2_19_port, 
                           pright => Psignal_2_17_port, pout => 
                           Psignal_3_19_port, gout => n13);
   PGblock_2_23 : PG_33 port map( gleft => Gsignal_2_23_port, gright => 
                           Gsignal_2_21_port, pleft => Psignal_2_23_port, 
                           pright => Psignal_2_21_port, pout => 
                           Psignal_3_23_port, gout => Gsignal_3_23_port);
   PGblock_2_27 : PG_32 port map( gleft => Gsignal_2_27_port, gright => 
                           Gsignal_2_25_port, pleft => Psignal_2_27_port, 
                           pright => Psignal_2_25_port, pout => 
                           Psignal_3_27_port, gout => n12);
   PGblock_2_31 : PG_31 port map( gleft => Gsignal_2_31_port, gright => 
                           Gsignal_2_29_port, pleft => Psignal_2_31_port, 
                           pright => Psignal_2_29_port, pout => 
                           Psignal_3_31_port, gout => Gsignal_3_31_port);
   Gblock_3_7 : G_14 port map( gleft => Gsignal_3_7_port, gright => Cout_1_port
                           , pleft => Psignal_3_7_port, gout => Cout_2_port);
   PGblock_3_15 : PG_30 port map( gleft => Gsignal_3_15_port, gright => n10, 
                           pleft => Psignal_3_15_port, pright => n8, pout => 
                           Psignal_4_15_port, gout => Gsignal_4_15_port);
   PGblock_3_23 : PG_4_0 port map( gleft => Gsignal_3_23_port, gright => n13, 
                           pleft => Psignal_3_23_port, pright => 
                           Psignal_3_19_port, pout => Psignal_4_23_port, gout 
                           => n15);
   PGblock_3_31 : PG_29 port map( gleft => Gsignal_3_31_port, gright => n12, 
                           pleft => Psignal_3_31_port, pright => 
                           Psignal_3_27_port, pout => Psignal_4_31_port, gout 
                           => Gsignal_4_31_port);
   Gblock_4_11 : G_6_0 port map( gleft => n10, gright => Cout_2_port, pleft => 
                           n8, gout => Cout_3_port);
   Gblock_4_15 : G_5_0 port map( gleft => Gsignal_4_15_port, gright => 
                           Cout_2_port, pleft => Psignal_4_15_port, gout => 
                           Cout_4_port);
   PGblock_4_27 : PG_28 port map( gleft => n12, gright => n15, pleft => 
                           Psignal_3_27_port, pright => Psignal_4_23_port, pout
                           => Psignal_5_27_port, gout => Gsignal_5_27_port);
   PGblock_4_31 : PG_27 port map( gleft => Gsignal_4_31_port, gright => n15, 
                           pleft => Psignal_4_31_port, pright => 
                           Psignal_4_23_port, pout => Psignal_5_31_port, gout 
                           => Gsignal_5_31_port);
   Gblock_5_19 : G_13 port map( gleft => n13, gright => Cout_4_port, pleft => 
                           Psignal_3_19_port, gout => Cout_5_port);
   Gblock_5_23 : G_12 port map( gleft => n15, gright => Cout_4_port, pleft => 
                           Psignal_4_23_port, gout => Cout_6_port);
   Gblock_5_27 : G_11 port map( gleft => Gsignal_5_27_port, gright => 
                           Cout_4_port, pleft => Psignal_5_27_port, gout => 
                           Cout_7_port);
   Gblock_5_31 : G_10 port map( gleft => Gsignal_5_31_port, gright => 
                           Cout_4_port, pleft => Psignal_5_31_port, gout => 
                           Cout_8_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_1;

architecture SYN_behav of xor_gate_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_2;

architecture SYN_behav of xor_gate_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_3;

architecture SYN_behav of xor_gate_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_4;

architecture SYN_behav of xor_gate_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_5;

architecture SYN_behav of xor_gate_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_6;

architecture SYN_behav of xor_gate_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_7;

architecture SYN_behav of xor_gate_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_8;

architecture SYN_behav of xor_gate_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_9;

architecture SYN_behav of xor_gate_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_10;

architecture SYN_behav of xor_gate_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_11;

architecture SYN_behav of xor_gate_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_12;

architecture SYN_behav of xor_gate_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_13;

architecture SYN_behav of xor_gate_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_14;

architecture SYN_behav of xor_gate_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_15;

architecture SYN_behav of xor_gate_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_16;

architecture SYN_behav of xor_gate_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_17;

architecture SYN_behav of xor_gate_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_18;

architecture SYN_behav of xor_gate_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_19;

architecture SYN_behav of xor_gate_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_20;

architecture SYN_behav of xor_gate_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_21;

architecture SYN_behav of xor_gate_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_22;

architecture SYN_behav of xor_gate_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_23;

architecture SYN_behav of xor_gate_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_24;

architecture SYN_behav of xor_gate_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_25;

architecture SYN_behav of xor_gate_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_26;

architecture SYN_behav of xor_gate_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_27;

architecture SYN_behav of xor_gate_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_28;

architecture SYN_behav of xor_gate_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_29;

architecture SYN_behav of xor_gate_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_30;

architecture SYN_behav of xor_gate_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_31;

architecture SYN_behav of xor_gate_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity xor_gate_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_0;

architecture SYN_behav of xor_gate_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH1 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_select_N4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4;

architecture SYN_STRUCTURAL of carry_select_N4 is

   component MUX21_GENERIC_N4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net61103, 
      net61104 : std_logic;

begin
   
   RCA0 : rca_generic_N4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net61104);
   RCA1 : rca_generic_N4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net61103);
   MUX : MUX21_GENERIC_N4 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PG is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG;

architecture SYN_STRUCTURAL of PG is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0 : std_logic;

begin
   
   C7 : GTECH_OR2 port map( A => gleft, B => N0, Z => gout);
   C8 : GTECH_AND2 port map( A => gright, B => pleft, Z => N0);
   C9 : GTECH_AND2 port map( A => pleft, B => pright, Z => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity G is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G;

architecture SYN_STRUCTURAL of G is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0 : std_logic;

begin
   
   C6 : GTECH_OR2 port map( A => gleft, B => N0, Z => gout);
   C7 : GTECH_AND2 port map( A => gright, B => pleft, Z => N0);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PGnet_block is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block;

architecture SYN_STRUCTURAL of PGnet_block is

   component GTECH_XOR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   C7 : GTECH_AND2 port map( A => A, B => B, Z => gout);
   C8 : GTECH_XOR2 port map( A => A, B => B, Z => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_thirdLevel is

   port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector (38 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end shift_thirdLevel;

architecture SYN_behav of shift_thirdLevel is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n40, n41, n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
      n56, n57, n58, n59, n60, n61, n62, n63, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(2), A2 => n148, ZN => n149);
   U2 : INV_X1 port map( A => n157, ZN => n156);
   U3 : INV_X1 port map( A => n149, ZN => n154);
   U4 : INV_X1 port map( A => n161, ZN => n158);
   U5 : INV_X1 port map( A => n153, ZN => n152);
   U6 : INV_X1 port map( A => n149, ZN => n155);
   U7 : OAI22_X1 port map( A1 => n165, A2 => n126, B1 => sel(0), B2 => n123, ZN
                           => Y(15));
   U8 : OAI22_X1 port map( A1 => n166, A2 => n129, B1 => sel(0), B2 => n126, ZN
                           => Y(14));
   U9 : OAI22_X1 port map( A1 => n166, A2 => n132, B1 => sel(0), B2 => n129, ZN
                           => Y(13));
   U10 : OAI22_X1 port map( A1 => n166, A2 => n135, B1 => sel(0), B2 => n132, 
                           ZN => Y(12));
   U11 : OAI22_X1 port map( A1 => n166, A2 => n138, B1 => sel(0), B2 => n135, 
                           ZN => Y(11));
   U12 : INV_X1 port map( A => n151, ZN => n150);
   U13 : OAI22_X1 port map( A1 => sel(0), A2 => n40, B1 => n41, B2 => n159, ZN 
                           => Y(9));
   U14 : OAI22_X1 port map( A1 => n161, A2 => n83, B1 => n158, B2 => n74, ZN =>
                           Y(29));
   U15 : OAI22_X1 port map( A1 => n162, A2 => n86, B1 => n158, B2 => n83, ZN =>
                           Y(28));
   U16 : OAI22_X1 port map( A1 => n162, A2 => n89, B1 => n158, B2 => n86, ZN =>
                           Y(27));
   U17 : OAI22_X1 port map( A1 => n162, A2 => n91, B1 => n158, B2 => n89, ZN =>
                           Y(26));
   U18 : OAI22_X1 port map( A1 => n162, A2 => n93, B1 => n158, B2 => n91, ZN =>
                           Y(25));
   U19 : OAI22_X1 port map( A1 => n163, A2 => n96, B1 => n158, B2 => n93, ZN =>
                           Y(24));
   U20 : OAI22_X1 port map( A1 => n163, A2 => n99, B1 => n158, B2 => n96, ZN =>
                           Y(23));
   U21 : OAI22_X1 port map( A1 => n163, A2 => n102, B1 => n158, B2 => n99, ZN 
                           => Y(22));
   U22 : OAI22_X1 port map( A1 => n164, A2 => n105, B1 => n158, B2 => n102, ZN 
                           => Y(21));
   U23 : OAI22_X1 port map( A1 => n164, A2 => n108, B1 => n158, B2 => n105, ZN 
                           => Y(20));
   U24 : OAI22_X1 port map( A1 => n164, A2 => n114, B1 => n158, B2 => n108, ZN 
                           => Y(19));
   U25 : OAI22_X1 port map( A1 => n165, A2 => n117, B1 => n158, B2 => n114, ZN 
                           => Y(18));
   U26 : OAI22_X1 port map( A1 => n165, A2 => n120, B1 => n158, B2 => n117, ZN 
                           => Y(17));
   U27 : OAI22_X1 port map( A1 => n165, A2 => n123, B1 => n158, B2 => n120, ZN 
                           => Y(16));
   U28 : OAI22_X1 port map( A1 => n159, A2 => n43, B1 => n158, B2 => n41, ZN =>
                           Y(8));
   U29 : OAI22_X1 port map( A1 => sel(0), A2 => n138, B1 => n159, B2 => n40, ZN
                           => Y(10));
   U30 : OAI221_X1 port map( B1 => A(13), B2 => n154, C1 => A(11), C2 => n44, A
                           => n142, ZN => n138);
   U31 : AOI22_X1 port map( A1 => n47, A2 => n50, B1 => n150, B2 => n137, ZN =>
                           n142);
   U32 : OAI221_X1 port map( B1 => A(20), B2 => n155, C1 => A(18), C2 => n156, 
                           A => n121, ZN => n117);
   U33 : AOI22_X1 port map( A1 => n152, A2 => n122, B1 => n150, B2 => n116, ZN 
                           => n121);
   U34 : OAI221_X1 port map( B1 => A(19), B2 => n154, C1 => A(17), C2 => n156, 
                           A => n124, ZN => n120);
   U35 : AOI22_X1 port map( A1 => n152, A2 => n125, B1 => n150, B2 => n119, ZN 
                           => n124);
   U36 : OAI221_X1 port map( B1 => A(18), B2 => n155, C1 => A(16), C2 => n156, 
                           A => n127, ZN => n123);
   U37 : AOI22_X1 port map( A1 => n152, A2 => n128, B1 => n150, B2 => n122, ZN 
                           => n127);
   U38 : OAI221_X1 port map( B1 => A(16), B2 => n154, C1 => A(14), C2 => n156, 
                           A => n133, ZN => n129);
   U39 : AOI22_X1 port map( A1 => n152, A2 => n134, B1 => n150, B2 => n128, ZN 
                           => n133);
   U40 : OAI221_X1 port map( B1 => A(15), B2 => n155, C1 => A(13), C2 => n156, 
                           A => n136, ZN => n132);
   U41 : AOI22_X1 port map( A1 => n152, A2 => n137, B1 => n150, B2 => n131, ZN 
                           => n136);
   U42 : OAI221_X1 port map( B1 => A(14), B2 => n154, C1 => A(12), C2 => n156, 
                           A => n139, ZN => n135);
   U43 : AOI22_X1 port map( A1 => n152, A2 => n140, B1 => n150, B2 => n134, ZN 
                           => n139);
   U44 : OAI221_X1 port map( B1 => A(12), B2 => n154, C1 => A(10), C2 => n156, 
                           A => n141, ZN => n40);
   U45 : AOI22_X1 port map( A1 => n152, A2 => n54, B1 => n150, B2 => n140, ZN 
                           => n141);
   U46 : OAI221_X1 port map( B1 => A(8), B2 => n44, C1 => A(10), C2 => n154, A 
                           => n52, ZN => n43);
   U47 : AOI22_X1 port map( A1 => n152, A2 => n53, B1 => n49, B2 => n54, ZN => 
                           n52);
   U48 : OAI221_X1 port map( B1 => A(32), B2 => n154, C1 => A(30), C2 => n156, 
                           A => n84, ZN => n74);
   U49 : AOI22_X1 port map( A1 => n152, A2 => n72, B1 => n49, B2 => n85, ZN => 
                           n84);
   U50 : INV_X1 port map( A => A(36), ZN => n85);
   U51 : OAI221_X1 port map( B1 => A(31), B2 => n155, C1 => A(29), C2 => n44, A
                           => n87, ZN => n83);
   U52 : AOI22_X1 port map( A1 => n152, A2 => n79, B1 => n49, B2 => n88, ZN => 
                           n87);
   U53 : INV_X1 port map( A => A(35), ZN => n88);
   U54 : OAI221_X1 port map( B1 => A(30), B2 => n155, C1 => A(28), C2 => n156, 
                           A => n90, ZN => n86);
   U55 : AOI22_X1 port map( A1 => n47, A2 => n73, B1 => n49, B2 => n72, ZN => 
                           n90);
   U56 : OAI221_X1 port map( B1 => A(29), B2 => n155, C1 => A(27), C2 => n44, A
                           => n92, ZN => n89);
   U57 : AOI22_X1 port map( A1 => n47, A2 => n77, B1 => n49, B2 => n79, ZN => 
                           n92);
   U58 : OAI221_X1 port map( B1 => A(28), B2 => n155, C1 => A(26), C2 => n156, 
                           A => n94, ZN => n91);
   U59 : AOI22_X1 port map( A1 => n47, A2 => n95, B1 => n49, B2 => n73, ZN => 
                           n94);
   U60 : OAI221_X1 port map( B1 => A(27), B2 => n155, C1 => A(25), C2 => n44, A
                           => n97, ZN => n93);
   U61 : AOI22_X1 port map( A1 => n47, A2 => n98, B1 => n49, B2 => n77, ZN => 
                           n97);
   U62 : OAI221_X1 port map( B1 => A(26), B2 => n155, C1 => A(24), C2 => n156, 
                           A => n100, ZN => n96);
   U63 : AOI22_X1 port map( A1 => n47, A2 => n101, B1 => n49, B2 => n95, ZN => 
                           n100);
   U64 : OAI221_X1 port map( B1 => A(25), B2 => n155, C1 => A(23), C2 => n44, A
                           => n103, ZN => n99);
   U65 : AOI22_X1 port map( A1 => n47, A2 => n104, B1 => n150, B2 => n98, ZN =>
                           n103);
   U66 : OAI221_X1 port map( B1 => A(24), B2 => n155, C1 => A(22), C2 => n156, 
                           A => n106, ZN => n102);
   U67 : AOI22_X1 port map( A1 => n47, A2 => n107, B1 => n150, B2 => n101, ZN 
                           => n106);
   U68 : OAI221_X1 port map( B1 => A(23), B2 => n155, C1 => A(21), C2 => n156, 
                           A => n109, ZN => n105);
   U69 : AOI22_X1 port map( A1 => n152, A2 => n110, B1 => n150, B2 => n104, ZN 
                           => n109);
   U70 : OAI221_X1 port map( B1 => A(22), B2 => n155, C1 => A(20), C2 => n156, 
                           A => n115, ZN => n108);
   U71 : AOI22_X1 port map( A1 => n152, A2 => n116, B1 => n150, B2 => n107, ZN 
                           => n115);
   U72 : OAI221_X1 port map( B1 => A(21), B2 => n155, C1 => A(19), C2 => n156, 
                           A => n118, ZN => n114);
   U73 : AOI22_X1 port map( A1 => n152, A2 => n119, B1 => n150, B2 => n110, ZN 
                           => n118);
   U74 : OAI221_X1 port map( B1 => A(17), B2 => n155, C1 => A(15), C2 => n156, 
                           A => n130, ZN => n126);
   U75 : AOI22_X1 port map( A1 => n152, A2 => n131, B1 => n150, B2 => n125, ZN 
                           => n130);
   U76 : OAI221_X1 port map( B1 => A(9), B2 => n44, C1 => A(11), C2 => n154, A 
                           => n46, ZN => n41);
   U77 : AOI22_X1 port map( A1 => n152, A2 => n48, B1 => n150, B2 => n50, ZN =>
                           n46);
   U78 : OAI22_X1 port map( A1 => n163, A2 => n74, B1 => n158, B2 => n69, ZN =>
                           Y(30));
   U79 : OAI22_X1 port map( A1 => n160, A2 => n51, B1 => n158, B2 => n43, ZN =>
                           Y(7));
   U80 : OAI22_X1 port map( A1 => n160, A2 => n55, B1 => n158, B2 => n51, ZN =>
                           Y(6));
   U81 : OAI22_X1 port map( A1 => n160, A2 => n58, B1 => n158, B2 => n55, ZN =>
                           Y(5));
   U82 : OAI22_X1 port map( A1 => n160, A2 => n61, B1 => n158, B2 => n58, ZN =>
                           Y(4));
   U83 : OAI22_X1 port map( A1 => n161, A2 => n66, B1 => sel(0), B2 => n61, ZN 
                           => Y(3));
   U84 : OAI22_X1 port map( A1 => n161, A2 => n80, B1 => sel(0), B2 => n66, ZN 
                           => Y(2));
   U85 : OAI22_X1 port map( A1 => n164, A2 => n111, B1 => n158, B2 => n80, ZN 
                           => Y(1));
   U86 : BUF_X1 port map( A => n167, Z => n160);
   U87 : BUF_X1 port map( A => n167, Z => n161);
   U88 : BUF_X1 port map( A => n165, Z => n162);
   U89 : INV_X1 port map( A => A(31), ZN => n77);
   U90 : INV_X1 port map( A => A(32), ZN => n73);
   U91 : BUF_X1 port map( A => n167, Z => n159);
   U92 : BUF_X1 port map( A => n166, Z => n163);
   U93 : BUF_X1 port map( A => n167, Z => n165);
   U94 : BUF_X1 port map( A => n167, Z => n166);
   U95 : BUF_X1 port map( A => n167, Z => n164);
   U96 : INV_X1 port map( A => A(30), ZN => n95);
   U97 : INV_X1 port map( A => A(29), ZN => n98);
   U98 : INV_X1 port map( A => A(28), ZN => n101);
   U99 : INV_X1 port map( A => A(27), ZN => n104);
   U100 : INV_X1 port map( A => A(26), ZN => n107);
   U101 : INV_X1 port map( A => A(25), ZN => n110);
   U102 : INV_X1 port map( A => A(24), ZN => n116);
   U103 : INV_X1 port map( A => A(23), ZN => n119);
   U104 : INV_X1 port map( A => A(22), ZN => n122);
   U105 : INV_X1 port map( A => A(21), ZN => n125);
   U106 : INV_X1 port map( A => A(20), ZN => n128);
   U107 : INV_X1 port map( A => A(19), ZN => n131);
   U108 : INV_X1 port map( A => A(18), ZN => n134);
   U109 : INV_X1 port map( A => A(17), ZN => n137);
   U110 : INV_X1 port map( A => A(16), ZN => n140);
   U111 : INV_X1 port map( A => A(15), ZN => n50);
   U112 : INV_X1 port map( A => A(14), ZN => n54);
   U113 : INV_X1 port map( A => A(13), ZN => n48);
   U114 : INV_X1 port map( A => A(12), ZN => n53);
   U115 : OAI221_X1 port map( B1 => A(1), B2 => n44, C1 => A(3), C2 => n154, A 
                           => n146, ZN => n111);
   U116 : INV_X1 port map( A => n147, ZN => n146);
   U117 : OAI22_X1 port map( A1 => n153, A2 => A(5), B1 => n151, B2 => A(7), ZN
                           => n147);
   U118 : OAI221_X1 port map( B1 => A(3), B2 => n44, C1 => A(5), C2 => n154, A 
                           => n81, ZN => n66);
   U119 : INV_X1 port map( A => n82, ZN => n81);
   U120 : OAI22_X1 port map( A1 => n153, A2 => A(7), B1 => n151, B2 => A(9), ZN
                           => n82);
   U121 : OAI221_X1 port map( B1 => A(2), B2 => n44, C1 => A(4), C2 => n154, A 
                           => n112, ZN => n80);
   U122 : INV_X1 port map( A => n113, ZN => n112);
   U123 : OAI22_X1 port map( A1 => n153, A2 => A(6), B1 => n151, B2 => A(8), ZN
                           => n113);
   U124 : OAI221_X1 port map( B1 => A(9), B2 => n154, C1 => A(7), C2 => n44, A 
                           => n56, ZN => n51);
   U125 : AOI22_X1 port map( A1 => n47, A2 => n57, B1 => n49, B2 => n48, ZN => 
                           n56);
   U126 : INV_X1 port map( A => A(11), ZN => n57);
   U127 : OAI221_X1 port map( B1 => A(8), B2 => n154, C1 => A(6), C2 => n44, A 
                           => n59, ZN => n55);
   U128 : AOI22_X1 port map( A1 => n152, A2 => n60, B1 => n150, B2 => n53, ZN 
                           => n59);
   U129 : INV_X1 port map( A => A(10), ZN => n60);
   U130 : OAI221_X1 port map( B1 => A(7), B2 => n154, C1 => A(5), C2 => n44, A 
                           => n62, ZN => n58);
   U131 : INV_X1 port map( A => n63, ZN => n62);
   U132 : OAI22_X1 port map( A1 => n153, A2 => A(9), B1 => n151, B2 => A(11), 
                           ZN => n63);
   U133 : OAI221_X1 port map( B1 => A(6), B2 => n154, C1 => A(4), C2 => n44, A 
                           => n67, ZN => n61);
   U134 : INV_X1 port map( A => n68, ZN => n67);
   U135 : OAI22_X1 port map( A1 => n153, A2 => A(8), B1 => n151, B2 => A(10), 
                           ZN => n68);
   U136 : OAI221_X1 port map( B1 => A(35), B2 => n153, C1 => A(37), C2 => n151,
                           A => n75, ZN => n69);
   U137 : AOI22_X1 port map( A1 => n157, A2 => n77, B1 => n149, B2 => n79, ZN 
                           => n75);
   U138 : OAI22_X1 port map( A1 => n161, A2 => n69, B1 => n158, B2 => n70, ZN 
                           => Y(31));
   U139 : AOI221_X1 port map( B1 => A(36), B2 => n47, C1 => A(38), C2 => n49, A
                           => n71, ZN => n70);
   U140 : OAI22_X1 port map( A1 => n154, A2 => n72, B1 => n44, B2 => n73, ZN =>
                           n71);
   U141 : OAI22_X1 port map( A1 => sel(0), A2 => n111, B1 => n143, B2 => n159, 
                           ZN => Y(0));
   U142 : AOI221_X1 port map( B1 => A(0), B2 => n157, C1 => A(2), C2 => n149, A
                           => n144, ZN => n143);
   U143 : INV_X1 port map( A => n145, ZN => n144);
   U144 : NOR2_X1 port map( A1 => sel(1), A2 => sel(2), ZN => n49);
   U145 : NOR2_X1 port map( A1 => n148, A2 => sel(2), ZN => n47);
   U146 : AOI22_X1 port map( A1 => n49, A2 => A(6), B1 => n47, B2 => A(4), ZN 
                           => n145);
   U147 : NAND2_X1 port map( A1 => sel(2), A2 => sel(1), ZN => n44);
   U148 : INV_X1 port map( A => A(33), ZN => n79);
   U149 : INV_X1 port map( A => A(34), ZN => n72);
   U150 : INV_X1 port map( A => sel(1), ZN => n148);
   U151 : INV_X1 port map( A => sel(0), ZN => n167);
   U152 : INV_X1 port map( A => n49, ZN => n151);
   U153 : INV_X1 port map( A => n47, ZN => n153);
   U154 : INV_X1 port map( A => n44, ZN => n157);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_secondLevel is

   port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : in 
         std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 downto 
         0));

end shift_secondLevel;

architecture SYN_behav of shift_secondLevel is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
      n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n90, Z => n93);
   U3 : BUF_X1 port map( A => n91, Z => n94);
   U4 : BUF_X1 port map( A => n90, Z => n92);
   U5 : BUF_X1 port map( A => n84, Z => n87);
   U6 : BUF_X1 port map( A => n85, Z => n88);
   U7 : BUF_X1 port map( A => n84, Z => n86);
   U8 : BUF_X1 port map( A => n96, Z => n99);
   U9 : BUF_X1 port map( A => n97, Z => n100);
   U10 : BUF_X1 port map( A => n96, Z => n98);
   U11 : BUF_X1 port map( A => n91, Z => n95);
   U12 : BUF_X1 port map( A => n85, Z => n89);
   U13 : BUF_X1 port map( A => n97, Z => n101);
   U14 : INV_X1 port map( A => n71, ZN => Y(1));
   U15 : INV_X1 port map( A => n52, ZN => Y(37));
   U16 : AOI222_X1 port map( A1 => mask00(37), A2 => n100, B1 => mask16(37), B2
                           => n94, C1 => mask08(37), C2 => n88, ZN => n52);
   U17 : INV_X1 port map( A => n51, ZN => Y(38));
   U18 : INV_X1 port map( A => n82, ZN => Y(0));
   U19 : INV_X1 port map( A => n41, ZN => Y(9));
   U20 : AOI222_X1 port map( A1 => mask00(9), A2 => n101, B1 => mask16(9), B2 
                           => n95, C1 => mask08(9), C2 => n89, ZN => n41);
   U21 : INV_X1 port map( A => n45, ZN => Y(8));
   U22 : AOI222_X1 port map( A1 => mask00(8), A2 => n101, B1 => mask16(8), B2 
                           => n95, C1 => mask08(8), C2 => n89, ZN => n45);
   U23 : INV_X1 port map( A => n80, ZN => Y(11));
   U24 : AOI222_X1 port map( A1 => mask00(11), A2 => n98, B1 => mask16(11), B2 
                           => n92, C1 => mask08(11), C2 => n86, ZN => n80);
   U25 : INV_X1 port map( A => n81, ZN => Y(10));
   U26 : AOI222_X1 port map( A1 => mask00(10), A2 => n98, B1 => mask16(10), B2 
                           => n92, C1 => mask08(10), C2 => n86, ZN => n81);
   U27 : INV_X1 port map( A => n59, ZN => Y(30));
   U28 : AOI222_X1 port map( A1 => mask00(30), A2 => n99, B1 => mask16(30), B2 
                           => n93, C1 => mask08(30), C2 => n87, ZN => n59);
   U29 : INV_X1 port map( A => n61, ZN => Y(29));
   U30 : AOI222_X1 port map( A1 => mask00(29), A2 => n99, B1 => mask16(29), B2 
                           => n93, C1 => mask08(29), C2 => n87, ZN => n61);
   U31 : INV_X1 port map( A => n62, ZN => Y(28));
   U32 : AOI222_X1 port map( A1 => mask00(28), A2 => n99, B1 => mask16(28), B2 
                           => n93, C1 => mask08(28), C2 => n87, ZN => n62);
   U33 : INV_X1 port map( A => n63, ZN => Y(27));
   U34 : AOI222_X1 port map( A1 => mask00(27), A2 => n99, B1 => mask16(27), B2 
                           => n93, C1 => mask08(27), C2 => n87, ZN => n63);
   U35 : INV_X1 port map( A => n64, ZN => Y(26));
   U36 : AOI222_X1 port map( A1 => mask00(26), A2 => n99, B1 => mask16(26), B2 
                           => n93, C1 => mask08(26), C2 => n87, ZN => n64);
   U37 : INV_X1 port map( A => n65, ZN => Y(25));
   U38 : AOI222_X1 port map( A1 => mask00(25), A2 => n99, B1 => mask16(25), B2 
                           => n93, C1 => mask08(25), C2 => n87, ZN => n65);
   U39 : INV_X1 port map( A => n66, ZN => Y(24));
   U40 : AOI222_X1 port map( A1 => mask00(24), A2 => n99, B1 => mask16(24), B2 
                           => n93, C1 => mask08(24), C2 => n87, ZN => n66);
   U41 : INV_X1 port map( A => n67, ZN => Y(23));
   U42 : AOI222_X1 port map( A1 => mask00(23), A2 => n99, B1 => mask16(23), B2 
                           => n93, C1 => mask08(23), C2 => n87, ZN => n67);
   U43 : INV_X1 port map( A => n68, ZN => Y(22));
   U44 : AOI222_X1 port map( A1 => mask00(22), A2 => n99, B1 => mask16(22), B2 
                           => n93, C1 => mask08(22), C2 => n87, ZN => n68);
   U45 : INV_X1 port map( A => n69, ZN => Y(21));
   U46 : AOI222_X1 port map( A1 => mask00(21), A2 => n99, B1 => mask16(21), B2 
                           => n93, C1 => mask08(21), C2 => n87, ZN => n69);
   U47 : INV_X1 port map( A => n70, ZN => Y(20));
   U48 : AOI222_X1 port map( A1 => mask00(20), A2 => n99, B1 => mask16(20), B2 
                           => n93, C1 => mask08(20), C2 => n87, ZN => n70);
   U49 : INV_X1 port map( A => n72, ZN => Y(19));
   U50 : AOI222_X1 port map( A1 => mask00(19), A2 => n98, B1 => mask16(19), B2 
                           => n92, C1 => mask08(19), C2 => n86, ZN => n72);
   U51 : INV_X1 port map( A => n73, ZN => Y(18));
   U52 : AOI222_X1 port map( A1 => mask00(18), A2 => n98, B1 => mask16(18), B2 
                           => n92, C1 => mask08(18), C2 => n86, ZN => n73);
   U53 : INV_X1 port map( A => n74, ZN => Y(17));
   U54 : AOI222_X1 port map( A1 => mask00(17), A2 => n98, B1 => mask16(17), B2 
                           => n92, C1 => mask08(17), C2 => n86, ZN => n74);
   U55 : INV_X1 port map( A => n75, ZN => Y(16));
   U56 : AOI222_X1 port map( A1 => mask00(16), A2 => n98, B1 => mask16(16), B2 
                           => n92, C1 => mask08(16), C2 => n86, ZN => n75);
   U57 : INV_X1 port map( A => n76, ZN => Y(15));
   U58 : AOI222_X1 port map( A1 => mask00(15), A2 => n98, B1 => mask16(15), B2 
                           => n92, C1 => mask08(15), C2 => n86, ZN => n76);
   U59 : INV_X1 port map( A => n77, ZN => Y(14));
   U60 : AOI222_X1 port map( A1 => mask00(14), A2 => n98, B1 => mask16(14), B2 
                           => n92, C1 => mask08(14), C2 => n86, ZN => n77);
   U61 : INV_X1 port map( A => n78, ZN => Y(13));
   U62 : AOI222_X1 port map( A1 => mask00(13), A2 => n98, B1 => mask16(13), B2 
                           => n92, C1 => mask08(13), C2 => n86, ZN => n78);
   U63 : INV_X1 port map( A => n79, ZN => Y(12));
   U64 : AOI222_X1 port map( A1 => mask00(12), A2 => n98, B1 => mask16(12), B2 
                           => n92, C1 => mask08(12), C2 => n86, ZN => n79);
   U65 : INV_X1 port map( A => n56, ZN => Y(33));
   U66 : AOI222_X1 port map( A1 => mask00(33), A2 => n100, B1 => mask16(33), B2
                           => n94, C1 => mask08(33), C2 => n88, ZN => n56);
   U67 : INV_X1 port map( A => n55, ZN => Y(34));
   U68 : AOI222_X1 port map( A1 => mask00(34), A2 => n100, B1 => mask16(34), B2
                           => n94, C1 => mask08(34), C2 => n88, ZN => n55);
   U69 : INV_X1 port map( A => n54, ZN => Y(35));
   U70 : AOI222_X1 port map( A1 => mask00(35), A2 => n100, B1 => mask16(35), B2
                           => n94, C1 => mask08(35), C2 => n88, ZN => n54);
   U71 : INV_X1 port map( A => n57, ZN => Y(32));
   U72 : AOI222_X1 port map( A1 => mask00(32), A2 => n100, B1 => mask16(32), B2
                           => n94, C1 => mask08(32), C2 => n88, ZN => n57);
   U73 : INV_X1 port map( A => n58, ZN => Y(31));
   U74 : AOI222_X1 port map( A1 => mask00(31), A2 => n100, B1 => mask16(31), B2
                           => n94, C1 => mask08(31), C2 => n88, ZN => n58);
   U75 : INV_X1 port map( A => n53, ZN => Y(36));
   U76 : AOI222_X1 port map( A1 => mask00(36), A2 => n100, B1 => mask16(36), B2
                           => n94, C1 => mask08(36), C2 => n88, ZN => n53);
   U77 : BUF_X1 port map( A => n42, Z => n96);
   U78 : BUF_X1 port map( A => n43, Z => n90);
   U79 : BUF_X1 port map( A => n44, Z => n84);
   U80 : BUF_X1 port map( A => n42, Z => n97);
   U81 : BUF_X1 port map( A => n43, Z => n91);
   U82 : BUF_X1 port map( A => n44, Z => n85);
   U83 : AOI222_X1 port map( A1 => mask00(38), A2 => n100, B1 => mask16(38), B2
                           => n94, C1 => mask08(38), C2 => n88, ZN => n51);
   U84 : AOI222_X1 port map( A1 => mask00(1), A2 => n98, B1 => mask16(1), B2 =>
                           n92, C1 => mask08(1), C2 => n86, ZN => n71);
   U85 : AOI222_X1 port map( A1 => mask00(0), A2 => n98, B1 => mask16(0), B2 =>
                           n92, C1 => mask08(0), C2 => n86, ZN => n82);
   U86 : INV_X1 port map( A => n47, ZN => Y(6));
   U87 : AOI222_X1 port map( A1 => mask00(6), A2 => n100, B1 => mask16(6), B2 
                           => n94, C1 => mask08(6), C2 => n88, ZN => n47);
   U88 : INV_X1 port map( A => n46, ZN => Y(7));
   U89 : AOI222_X1 port map( A1 => mask00(7), A2 => n101, B1 => mask16(7), B2 
                           => n95, C1 => mask08(7), C2 => n89, ZN => n46);
   U90 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n42);
   U91 : NOR2_X1 port map( A1 => n83, A2 => sel(0), ZN => n43);
   U92 : INV_X1 port map( A => n49, ZN => Y(4));
   U93 : AOI222_X1 port map( A1 => mask00(4), A2 => n100, B1 => mask16(4), B2 
                           => n94, C1 => mask08(4), C2 => n88, ZN => n49);
   U94 : INV_X1 port map( A => n48, ZN => Y(5));
   U95 : AOI222_X1 port map( A1 => mask00(5), A2 => n100, B1 => mask16(5), B2 
                           => n94, C1 => mask08(5), C2 => n88, ZN => n48);
   U96 : INV_X1 port map( A => n60, ZN => Y(2));
   U97 : AOI222_X1 port map( A1 => mask00(2), A2 => n99, B1 => mask16(2), B2 =>
                           n93, C1 => mask08(2), C2 => n87, ZN => n60);
   U98 : INV_X1 port map( A => n50, ZN => Y(3));
   U99 : AOI222_X1 port map( A1 => mask00(3), A2 => n100, B1 => mask16(3), B2 
                           => n94, C1 => mask08(3), C2 => n88, ZN => n50);
   U100 : INV_X1 port map( A => sel(1), ZN => n83);
   U101 : AND2_X1 port map( A1 => sel(0), A2 => n83, ZN => n44);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_firstLevel is

   port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector (1 
         downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 downto 
         0));

end shift_firstLevel;

architecture SYN_behav of shift_firstLevel is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask08_23_port, mask08_22_port, mask08_21_port, mask08_20_port, 
      mask08_19_port, mask08_18_port, mask08_17_port, mask08_16_port, 
      mask08_15_port, mask08_7_port, mask08_6_port, mask08_5_port, 
      mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port, mask08_0_port
      , mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n98, n116, n117, mask16_22_port, n119, n120, n121 : std_logic
      ;

begin
   mask08 <= ( mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask08_23_port, 
      mask08_22_port, mask08_21_port, mask08_20_port, mask08_19_port, 
      mask08_18_port, mask08_17_port, mask08_16_port, mask08_15_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port, mask08_7_port, mask08_6_port, 
      mask08_5_port, mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port
      , mask08_0_port );
   mask16 <= ( mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_22_port, mask16_22_port, mask16_22_port, mask16_22_port, 
      mask16_22_port, mask16_22_port, mask16_22_port, mask16_15_port, 
      mask16_14_port, mask16_13_port, mask16_12_port, mask16_11_port, 
      mask16_10_port, mask16_9_port, mask16_8_port, mask16_7_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port );
   
   U161 : NAND3_X1 port map( A1 => sel(1), A2 => n108, A3 => A(31), ZN => n61);
   U2 : INV_X1 port map( A => n116, ZN => n98);
   U3 : INV_X1 port map( A => mask16_22_port, ZN => n117);
   U4 : BUF_X1 port map( A => n59, Z => n121);
   U5 : BUF_X1 port map( A => n59, Z => n120);
   U6 : BUF_X1 port map( A => n59, Z => n119);
   U7 : INV_X1 port map( A => mask16_7_port, ZN => n94);
   U8 : INV_X1 port map( A => mask08_6_port, ZN => n111);
   U9 : INV_X1 port map( A => mask08_1_port, ZN => n96);
   U10 : INV_X1 port map( A => mask08_5_port, ZN => n112);
   U11 : INV_X1 port map( A => mask08_4_port, ZN => n113);
   U12 : INV_X1 port map( A => mask08_3_port, ZN => n114);
   U13 : INV_X1 port map( A => mask08_2_port, ZN => n115);
   U14 : OAI21_X1 port map( B1 => n120, B2 => n60, A => n117, ZN => 
                           mask16_38_port);
   U15 : OAI21_X1 port map( B1 => n120, B2 => n63, A => n117, ZN => 
                           mask16_36_port);
   U16 : OAI21_X1 port map( B1 => n120, B2 => n64, A => n117, ZN => 
                           mask16_35_port);
   U17 : OAI21_X1 port map( B1 => n120, B2 => n65, A => n117, ZN => 
                           mask16_34_port);
   U18 : OAI21_X1 port map( B1 => n120, B2 => n66, A => n117, ZN => 
                           mask16_33_port);
   U19 : OAI21_X1 port map( B1 => n120, B2 => n67, A => n117, ZN => 
                           mask16_32_port);
   U20 : OAI21_X1 port map( B1 => n120, B2 => n62, A => n117, ZN => 
                           mask16_37_port);
   U21 : NOR2_X1 port map( A1 => n86, A2 => n116, ZN => mask16_7_port);
   U22 : NOR2_X1 port map( A1 => n60, A2 => n116, ZN => mask08_7_port);
   U23 : NOR2_X1 port map( A1 => n62, A2 => n116, ZN => mask08_6_port);
   U24 : NOR2_X1 port map( A1 => n67, A2 => n116, ZN => mask08_1_port);
   U25 : NOR2_X1 port map( A1 => n65, A2 => n116, ZN => mask08_3_port);
   U26 : NOR2_X1 port map( A1 => n66, A2 => n116, ZN => mask08_2_port);
   U27 : NOR2_X1 port map( A1 => n63, A2 => n116, ZN => mask08_5_port);
   U28 : NOR2_X1 port map( A1 => n64, A2 => n116, ZN => mask08_4_port);
   U29 : INV_X1 port map( A => n61, ZN => mask16_22_port);
   U30 : INV_X1 port map( A => n53, ZN => mask16_9_port);
   U31 : NAND2_X1 port map( A1 => n96, A2 => n75, ZN => mask00(9));
   U32 : INV_X1 port map( A => n54, ZN => mask16_8_port);
   U33 : NAND2_X1 port map( A1 => n95, A2 => n76, ZN => mask00(8));
   U34 : INV_X1 port map( A => n83, ZN => mask16_11_port);
   U35 : NAND2_X1 port map( A1 => n114, A2 => n73, ZN => mask00(11));
   U36 : INV_X1 port map( A => n84, ZN => mask16_10_port);
   U37 : NAND2_X1 port map( A1 => n115, A2 => n74, ZN => mask00(10));
   U38 : OAI21_X1 port map( B1 => n121, B2 => n93, A => n94, ZN => mask00(23));
   U39 : OAI21_X1 port map( B1 => n87, B2 => n119, A => n117, ZN => 
                           mask08_37_port);
   U40 : INV_X1 port map( A => n97, ZN => n59);
   U41 : NAND2_X1 port map( A1 => n61, A2 => n69, ZN => mask16_30_port);
   U42 : OAI21_X1 port map( B1 => n86, B2 => n119, A => n80, ZN => mask00(30));
   U43 : NAND2_X1 port map( A1 => n61, A2 => n71, ZN => mask16_29_port);
   U44 : OAI21_X1 port map( B1 => n87, B2 => n119, A => n81, ZN => mask00(29));
   U45 : NAND2_X1 port map( A1 => n61, A2 => n72, ZN => mask16_28_port);
   U46 : OAI21_X1 port map( B1 => n88, B2 => n119, A => n82, ZN => mask00(28));
   U47 : NAND2_X1 port map( A1 => n61, A2 => n73, ZN => mask16_27_port);
   U48 : OAI21_X1 port map( B1 => n89, B2 => n119, A => n83, ZN => mask00(27));
   U49 : NAND2_X1 port map( A1 => n61, A2 => n74, ZN => mask16_26_port);
   U50 : OAI21_X1 port map( B1 => n90, B2 => n119, A => n84, ZN => mask00(26));
   U51 : NAND2_X1 port map( A1 => n61, A2 => n75, ZN => mask16_25_port);
   U52 : OAI21_X1 port map( B1 => n121, B2 => n91, A => n53, ZN => mask00(25));
   U53 : NAND2_X1 port map( A1 => n117, A2 => n76, ZN => mask16_24_port);
   U54 : OAI21_X1 port map( B1 => n121, B2 => n92, A => n54, ZN => mask00(24));
   U55 : NAND2_X1 port map( A1 => n79, A2 => n68, ZN => mask08_23_port);
   U56 : NAND2_X1 port map( A1 => n61, A2 => n77, ZN => mask16_23_port);
   U57 : NAND2_X1 port map( A1 => n80, A2 => n69, ZN => mask08_22_port);
   U58 : OAI21_X1 port map( B1 => n121, B2 => n60, A => n55, ZN => mask00(22));
   U59 : NAND2_X1 port map( A1 => n81, A2 => n71, ZN => mask08_21_port);
   U60 : OAI21_X1 port map( B1 => n121, B2 => n62, A => n56, ZN => mask00(21));
   U61 : NAND2_X1 port map( A1 => n82, A2 => n72, ZN => mask08_20_port);
   U62 : OAI21_X1 port map( B1 => n121, B2 => n63, A => n57, ZN => mask00(20));
   U63 : NAND2_X1 port map( A1 => n83, A2 => n73, ZN => mask08_19_port);
   U64 : OAI21_X1 port map( B1 => n121, B2 => n64, A => n58, ZN => mask00(19));
   U65 : NAND2_X1 port map( A1 => n84, A2 => n74, ZN => mask08_18_port);
   U66 : OAI21_X1 port map( B1 => n121, B2 => n65, A => n70, ZN => mask00(18));
   U67 : NAND2_X1 port map( A1 => n53, A2 => n75, ZN => mask08_17_port);
   U68 : OAI21_X1 port map( B1 => n121, B2 => n66, A => n78, ZN => mask00(17));
   U69 : NAND2_X1 port map( A1 => n54, A2 => n76, ZN => mask08_16_port);
   U70 : OAI21_X1 port map( B1 => n120, B2 => n67, A => n85, ZN => mask00(16));
   U71 : INV_X1 port map( A => n79, ZN => mask16_15_port);
   U72 : NAND2_X1 port map( A1 => n94, A2 => n77, ZN => mask08_15_port);
   U73 : INV_X1 port map( A => n80, ZN => mask16_14_port);
   U74 : NAND2_X1 port map( A1 => n111, A2 => n69, ZN => mask00(14));
   U75 : INV_X1 port map( A => n81, ZN => mask16_13_port);
   U76 : NAND2_X1 port map( A1 => n112, A2 => n71, ZN => mask00(13));
   U77 : INV_X1 port map( A => n82, ZN => mask16_12_port);
   U78 : NAND2_X1 port map( A1 => n113, A2 => n72, ZN => mask00(12));
   U79 : OAI21_X1 port map( B1 => n120, B2 => n91, A => n61, ZN => 
                           mask08_33_port);
   U80 : OAI21_X1 port map( B1 => n90, B2 => n119, A => n117, ZN => 
                           mask08_34_port);
   U81 : OAI21_X1 port map( B1 => n89, B2 => n119, A => n117, ZN => 
                           mask08_35_port);
   U82 : OAI21_X1 port map( B1 => n121, B2 => n104, A => n61, ZN => mask00(35))
                           ;
   U83 : OAI21_X1 port map( B1 => n120, B2 => n92, A => n117, ZN => 
                           mask08_32_port);
   U84 : OAI21_X1 port map( B1 => n107, B2 => n119, A => n117, ZN => mask00(32)
                           );
   U85 : NAND2_X1 port map( A1 => n61, A2 => n68, ZN => mask16_31_port);
   U86 : OAI21_X1 port map( B1 => n120, B2 => n93, A => n61, ZN => 
                           mask08_31_port);
   U87 : OAI21_X1 port map( B1 => n88, B2 => n119, A => n117, ZN => 
                           mask08_36_port);
   U88 : OAI21_X1 port map( B1 => n121, B2 => n103, A => n117, ZN => mask00(36)
                           );
   U89 : INV_X1 port map( A => n55, ZN => mask16_6_port);
   U90 : INV_X1 port map( A => n56, ZN => mask16_5_port);
   U91 : INV_X1 port map( A => n57, ZN => mask16_4_port);
   U92 : INV_X1 port map( A => n58, ZN => mask16_3_port);
   U93 : INV_X1 port map( A => n78, ZN => mask16_1_port);
   U94 : INV_X1 port map( A => n85, ZN => mask16_0_port);
   U95 : INV_X1 port map( A => n70, ZN => mask16_2_port);
   U96 : NAND2_X1 port map( A1 => n110, A2 => n68, ZN => mask00(15));
   U97 : INV_X1 port map( A => mask08_7_port, ZN => n110);
   U98 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n97);
   U99 : OAI21_X1 port map( B1 => n86, B2 => n119, A => n117, ZN => 
                           mask08_38_port);
   U100 : OAI21_X1 port map( B1 => n120, B2 => n101, A => n61, ZN => mask00(38)
                           );
   U101 : INV_X1 port map( A => A(31), ZN => n101);
   U102 : AND2_X1 port map( A1 => n99, A2 => A(1), ZN => mask00(1));
   U103 : INV_X1 port map( A => n95, ZN => mask08_0_port);
   U104 : AND2_X1 port map( A1 => n99, A2 => A(0), ZN => mask00(0));
   U105 : INV_X1 port map( A => sel(0), ZN => n108);
   U106 : AOI21_X1 port map( B1 => sel(0), B2 => sel(1), A => n97, ZN => n99);
   U107 : NAND2_X1 port map( A1 => A(8), A2 => n97, ZN => n68);
   U108 : NAND2_X1 port map( A1 => A(7), A2 => n97, ZN => n69);
   U109 : NAND2_X1 port map( A1 => A(2), A2 => n97, ZN => n75);
   U110 : NAND2_X1 port map( A1 => A(1), A2 => n97, ZN => n76);
   U111 : NAND2_X1 port map( A1 => A(6), A2 => n97, ZN => n71);
   U112 : NAND2_X1 port map( A1 => A(5), A2 => n97, ZN => n72);
   U113 : NAND2_X1 port map( A1 => A(4), A2 => n97, ZN => n73);
   U114 : NAND2_X1 port map( A1 => A(3), A2 => n97, ZN => n74);
   U115 : AND2_X1 port map( A1 => n99, A2 => A(6), ZN => mask00(6));
   U116 : NAND2_X1 port map( A1 => A(0), A2 => n97, ZN => n77);
   U117 : OAI21_X1 port map( B1 => n116, B2 => n100, A => n77, ZN => mask00(7))
                           ;
   U118 : INV_X1 port map( A => A(7), ZN => n100);
   U119 : NAND2_X1 port map( A1 => A(31), A2 => n98, ZN => n79);
   U120 : NAND2_X1 port map( A1 => A(30), A2 => n98, ZN => n80);
   U121 : NAND2_X1 port map( A1 => A(25), A2 => n98, ZN => n53);
   U122 : NAND2_X1 port map( A1 => A(24), A2 => n98, ZN => n54);
   U123 : NAND2_X1 port map( A1 => A(29), A2 => n98, ZN => n81);
   U124 : NAND2_X1 port map( A1 => A(28), A2 => n98, ZN => n82);
   U125 : NAND2_X1 port map( A1 => A(27), A2 => n98, ZN => n83);
   U126 : NAND2_X1 port map( A1 => A(26), A2 => n98, ZN => n84);
   U127 : OAI21_X1 port map( B1 => n109, B2 => n119, A => n79, ZN => mask00(31)
                           );
   U128 : INV_X1 port map( A => A(24), ZN => n109);
   U129 : OAI21_X1 port map( B1 => n121, B2 => n105, A => n61, ZN => mask00(34)
                           );
   U130 : INV_X1 port map( A => A(27), ZN => n105);
   U131 : OAI21_X1 port map( B1 => n121, B2 => n106, A => n61, ZN => mask00(33)
                           );
   U132 : INV_X1 port map( A => A(26), ZN => n106);
   U133 : OAI21_X1 port map( B1 => n120, B2 => n102, A => n61, ZN => mask00(37)
                           );
   U134 : INV_X1 port map( A => A(30), ZN => n102);
   U135 : NAND2_X1 port map( A1 => A(21), A2 => n98, ZN => n56);
   U136 : NAND2_X1 port map( A1 => A(20), A2 => n98, ZN => n57);
   U137 : NAND2_X1 port map( A1 => A(19), A2 => n98, ZN => n58);
   U138 : NAND2_X1 port map( A1 => A(22), A2 => n98, ZN => n55);
   U139 : AND2_X1 port map( A1 => n99, A2 => A(4), ZN => mask00(4));
   U140 : AND2_X1 port map( A1 => n99, A2 => A(5), ZN => mask00(5));
   U141 : INV_X1 port map( A => A(15), ZN => n60);
   U142 : INV_X1 port map( A => A(14), ZN => n62);
   U143 : INV_X1 port map( A => A(9), ZN => n67);
   U144 : INV_X1 port map( A => A(11), ZN => n65);
   U145 : INV_X1 port map( A => A(10), ZN => n66);
   U146 : INV_X1 port map( A => A(13), ZN => n63);
   U147 : INV_X1 port map( A => A(12), ZN => n64);
   U148 : INV_X1 port map( A => A(23), ZN => n86);
   U149 : NAND2_X1 port map( A1 => A(18), A2 => n99, ZN => n70);
   U150 : NAND2_X1 port map( A1 => A(17), A2 => n99, ZN => n78);
   U151 : NAND2_X1 port map( A1 => A(16), A2 => n99, ZN => n85);
   U152 : NAND2_X1 port map( A1 => A(8), A2 => n99, ZN => n95);
   U153 : AND2_X1 port map( A1 => n99, A2 => A(2), ZN => mask00(2));
   U154 : AND2_X1 port map( A1 => n99, A2 => A(3), ZN => mask00(3));
   U155 : INV_X1 port map( A => A(18), ZN => n91);
   U156 : INV_X1 port map( A => A(17), ZN => n92);
   U157 : INV_X1 port map( A => A(16), ZN => n93);
   U158 : INV_X1 port map( A => A(22), ZN => n87);
   U159 : INV_X1 port map( A => A(21), ZN => n88);
   U160 : INV_X1 port map( A => A(20), ZN => n89);
   U162 : INV_X1 port map( A => A(19), ZN => n90);
   U163 : INV_X1 port map( A => A(29), ZN => n103);
   U164 : INV_X1 port map( A => A(28), ZN => n104);
   U165 : INV_X1 port map( A => A(25), ZN => n107);
   U166 : INV_X1 port map( A => n99, ZN => n116);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity cla_adder_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end cla_adder_N32_1;

architecture SYN_struct of cla_adder_N32_1 is

   component sum_generator_Nbits32_Nblocks8_1
      port( A, B : in std_logic_vector (31 downto 0);  Carry : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_Nblocks8_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal Carry_8_port, Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port,
      Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port : std_logic;

begin
   
   CG : carry_generator_N32_Nblocks8_1 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci, Cout(8) => 
                           Carry_8_port, Cout(7) => Carry_7_port, Cout(6) => 
                           Carry_6_port, Cout(5) => Carry_5_port, Cout(4) => 
                           Carry_4_port, Cout(3) => Carry_3_port, Cout(2) => 
                           Carry_2_port, Cout(1) => Carry_1_port, Cout(0) => 
                           Carry_0_port);
   SG : sum_generator_Nbits32_Nblocks8_1 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Carry(8) => Carry_8_port, 
                           Carry(7) => Carry_7_port, Carry(6) => Carry_6_port, 
                           Carry(5) => Carry_5_port, Carry(4) => Carry_4_port, 
                           Carry(3) => Carry_3_port, Carry(2) => Carry_2_port, 
                           Carry(1) => Carry_1_port, Carry(0) => Carry_0_port, 
                           S(31) => Sum(31), S(30) => Sum(30), S(29) => Sum(29)
                           , S(28) => Sum(28), S(27) => Sum(27), S(26) => 
                           Sum(26), S(25) => Sum(25), S(24) => Sum(24), S(23) 
                           => Sum(23), S(22) => Sum(22), S(21) => Sum(21), 
                           S(20) => Sum(20), S(19) => Sum(19), S(18) => Sum(18)
                           , S(17) => Sum(17), S(16) => Sum(16), S(15) => 
                           Sum(15), S(14) => Sum(14), S(13) => Sum(13), S(12) 
                           => Sum(12), S(11) => Sum(11), S(10) => Sum(10), S(9)
                           => Sum(9), S(8) => Sum(8), S(7) => Sum(7), S(6) => 
                           Sum(6), S(5) => Sum(5), S(4) => Sum(4), S(3) => 
                           Sum(3), S(2) => Sum(2), S(1) => Sum(1), S(0) => 
                           Sum(0), Cout => Cout);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_1;

architecture SYN_struct of CSA_Nbits32_1 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_96 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co 
                           => Cout(1));
   FullAdd_1 : FA_95 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co 
                           => Cout(2));
   FullAdd_2 : FA_94 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co 
                           => Cout(3));
   FullAdd_3 : FA_93 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co 
                           => Cout(4));
   FullAdd_4 : FA_92 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co 
                           => Cout(5));
   FullAdd_5 : FA_91 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co 
                           => Cout(6));
   FullAdd_6 : FA_90 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co 
                           => Cout(7));
   FullAdd_7 : FA_89 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co 
                           => Cout(8));
   FullAdd_8 : FA_88 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co 
                           => Cout(9));
   FullAdd_9 : FA_87 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co 
                           => Cout(10));
   FullAdd_10 : FA_86 port map( A => A(10), B => B(10), Ci => C(10), S => S(10)
                           , Co => Cout(11));
   FullAdd_11 : FA_85 port map( A => A(11), B => B(11), Ci => C(11), S => S(11)
                           , Co => Cout(12));
   FullAdd_12 : FA_84 port map( A => A(12), B => B(12), Ci => C(12), S => S(12)
                           , Co => Cout(13));
   FullAdd_13 : FA_83 port map( A => A(13), B => B(13), Ci => C(13), S => S(13)
                           , Co => Cout(14));
   FullAdd_14 : FA_82 port map( A => A(14), B => B(14), Ci => C(14), S => S(14)
                           , Co => Cout(15));
   FullAdd_15 : FA_81 port map( A => A(15), B => B(15), Ci => C(15), S => S(15)
                           , Co => Cout(16));
   FullAdd_16 : FA_80 port map( A => A(16), B => B(16), Ci => C(16), S => S(16)
                           , Co => Cout(17));
   FullAdd_17 : FA_79 port map( A => A(17), B => B(17), Ci => C(17), S => S(17)
                           , Co => Cout(18));
   FullAdd_18 : FA_78 port map( A => A(18), B => B(18), Ci => C(18), S => S(18)
                           , Co => Cout(19));
   FullAdd_19 : FA_77 port map( A => A(19), B => B(19), Ci => C(19), S => S(19)
                           , Co => Cout(20));
   FullAdd_20 : FA_76 port map( A => A(20), B => B(20), Ci => C(20), S => S(20)
                           , Co => Cout(21));
   FullAdd_21 : FA_75 port map( A => A(21), B => B(21), Ci => C(21), S => S(21)
                           , Co => Cout(22));
   FullAdd_22 : FA_74 port map( A => A(22), B => B(22), Ci => C(22), S => S(22)
                           , Co => Cout(23));
   FullAdd_23 : FA_73 port map( A => A(23), B => B(23), Ci => C(23), S => S(23)
                           , Co => Cout(24));
   FullAdd_24 : FA_72 port map( A => A(24), B => B(24), Ci => C(24), S => S(24)
                           , Co => Cout(25));
   FullAdd_25 : FA_71 port map( A => A(25), B => B(25), Ci => C(25), S => S(25)
                           , Co => Cout(26));
   FullAdd_26 : FA_70 port map( A => A(26), B => B(26), Ci => C(26), S => S(26)
                           , Co => Cout(27));
   FullAdd_27 : FA_69 port map( A => A(27), B => B(27), Ci => C(27), S => S(27)
                           , Co => Cout(28));
   FullAdd_28 : FA_68 port map( A => A(28), B => B(28), Ci => C(28), S => S(28)
                           , Co => Cout(29));
   FullAdd_29 : FA_67 port map( A => A(29), B => B(29), Ci => C(29), S => S(29)
                           , Co => Cout(30));
   FullAdd_30 : FA_66 port map( A => A(30), B => B(30), Ci => C(30), S => S(30)
                           , Co => Cout(31));
   LastFA : FA_65 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), Co
                           => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_2;

architecture SYN_struct of CSA_Nbits32_2 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_128 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_127 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_126 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_125 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_124 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_123 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_122 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_121 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_120 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_119 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_118 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_117 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_116 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_115 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_114 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_113 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_112 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_111 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_110 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_109 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_108 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_107 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_106 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_105 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_104 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_103 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_102 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_101 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_100 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_99 port map( A => A(29), B => B(29), Ci => C(29), S => S(29)
                           , Co => Cout(30));
   FullAdd_30 : FA_98 port map( A => A(30), B => B(30), Ci => C(30), S => S(30)
                           , Co => Cout(31));
   LastFA : FA_97 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), Co
                           => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_3;

architecture SYN_struct of CSA_Nbits32_3 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_160 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_159 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_158 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_157 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_156 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_155 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_154 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_153 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_152 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_151 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_150 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_149 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_148 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_147 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_146 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_145 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_144 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_143 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_142 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_141 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_140 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_139 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_138 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_137 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_136 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_135 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_134 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_133 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_132 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_131 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_130 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_129 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_4 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_4;

architecture SYN_struct of CSA_Nbits32_4 is

   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_192 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_191 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_190 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_189 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_188 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_187 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_186 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_185 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_184 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_183 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_182 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_181 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_180 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_179 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_178 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_177 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_176 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_175 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_174 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_173 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_172 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_171 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_170 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_169 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_168 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_167 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_166 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_165 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_164 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_163 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_162 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_161 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_5 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_5;

architecture SYN_struct of CSA_Nbits32_5 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_224 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_223 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_222 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_221 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_220 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_219 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_218 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_217 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_216 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_215 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_214 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_213 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_212 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_211 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_210 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_209 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_208 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_207 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_206 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_205 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_204 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_203 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_202 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_201 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_200 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_199 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_198 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_197 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_196 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_195 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_194 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_193 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CSA_Nbits32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_0;

architecture SYN_struct of CSA_Nbits32_0 is

   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_64 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co 
                           => Cout(1));
   FullAdd_1 : FA_255 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_254 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_253 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_252 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_251 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_250 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_249 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_248 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_247 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_246 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_245 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_244 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_243 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_242 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_241 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_240 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_239 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_238 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_237 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_236 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_235 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_234 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_233 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_232 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_231 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_230 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_229 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_228 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_227 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_226 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_225 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_1 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_1;

architecture SYN_behav of mux_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n257);
   U2 : BUF_X1 port map( A => n10, Z => n256);
   U3 : BUF_X1 port map( A => n10, Z => n258);
   U4 : BUF_X1 port map( A => n6, Z => n269);
   U5 : BUF_X1 port map( A => n6, Z => n268);
   U6 : BUF_X1 port map( A => n9, Z => n260);
   U7 : BUF_X1 port map( A => n9, Z => n259);
   U8 : BUF_X1 port map( A => n7, Z => n266);
   U9 : BUF_X1 port map( A => n7, Z => n265);
   U10 : BUF_X1 port map( A => n8, Z => n263);
   U11 : BUF_X1 port map( A => n8, Z => n262);
   U12 : BUF_X1 port map( A => n9, Z => n261);
   U13 : BUF_X1 port map( A => n7, Z => n267);
   U14 : BUF_X1 port map( A => n8, Z => n264);
   U15 : BUF_X1 port map( A => n6, Z => n270);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U23 : AOI22_X1 port map( A1 => A(28), A2 => n260, B1 => B(28), B2 => n257, 
                           ZN => n31);
   U24 : AOI222_X1 port map( A1 => D(28), A2 => n269, B1 => E(28), B2 => n266, 
                           C1 => C(28), C2 => n263, ZN => n32);
   U25 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U26 : AOI22_X1 port map( A1 => A(14), A2 => n259, B1 => B(14), B2 => n256, 
                           ZN => n61);
   U27 : AOI222_X1 port map( A1 => D(14), A2 => n268, B1 => E(14), B2 => n265, 
                           C1 => C(14), C2 => n262, ZN => n62);
   U28 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U29 : AOI22_X1 port map( A1 => A(24), A2 => n260, B1 => B(24), B2 => n257, 
                           ZN => n39);
   U30 : AOI222_X1 port map( A1 => D(24), A2 => n269, B1 => E(24), B2 => n266, 
                           C1 => C(24), C2 => n263, ZN => n40);
   U31 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U32 : AOI22_X1 port map( A1 => A(18), A2 => n259, B1 => B(18), B2 => n256, 
                           ZN => n53);
   U33 : AOI222_X1 port map( A1 => D(18), A2 => n268, B1 => E(18), B2 => n265, 
                           C1 => C(18), C2 => n262, ZN => n54);
   U34 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n259, B1 => B(15), B2 => n256, 
                           ZN => n59);
   U36 : AOI222_X1 port map( A1 => D(15), A2 => n268, B1 => E(15), B2 => n265, 
                           C1 => C(15), C2 => n262, ZN => n60);
   U37 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U38 : AOI22_X1 port map( A1 => A(22), A2 => n260, B1 => B(22), B2 => n257, 
                           ZN => n43);
   U39 : AOI222_X1 port map( A1 => D(22), A2 => n269, B1 => E(22), B2 => n266, 
                           C1 => C(22), C2 => n263, ZN => n44);
   U40 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U41 : AOI22_X1 port map( A1 => A(16), A2 => n259, B1 => B(16), B2 => n256, 
                           ZN => n57);
   U42 : AOI222_X1 port map( A1 => D(16), A2 => n268, B1 => E(16), B2 => n265, 
                           C1 => C(16), C2 => n262, ZN => n58);
   U43 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U44 : AOI22_X1 port map( A1 => A(20), A2 => n260, B1 => B(20), B2 => n257, 
                           ZN => n47);
   U45 : AOI222_X1 port map( A1 => D(20), A2 => n269, B1 => E(20), B2 => n266, 
                           C1 => C(20), C2 => n263, ZN => n48);
   U46 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U47 : AOI22_X1 port map( A1 => A(27), A2 => n260, B1 => B(27), B2 => n257, 
                           ZN => n33);
   U48 : AOI222_X1 port map( A1 => D(27), A2 => n269, B1 => E(27), B2 => n266, 
                           C1 => C(27), C2 => n263, ZN => n34);
   U49 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U50 : AOI22_X1 port map( A1 => A(23), A2 => n260, B1 => B(23), B2 => n257, 
                           ZN => n41);
   U51 : AOI222_X1 port map( A1 => D(23), A2 => n269, B1 => E(23), B2 => n266, 
                           C1 => C(23), C2 => n263, ZN => n42);
   U52 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U53 : AOI22_X1 port map( A1 => A(17), A2 => n259, B1 => B(17), B2 => n256, 
                           ZN => n55);
   U54 : AOI222_X1 port map( A1 => D(17), A2 => n268, B1 => E(17), B2 => n265, 
                           C1 => C(17), C2 => n262, ZN => n56);
   U55 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U56 : AOI22_X1 port map( A1 => A(21), A2 => n260, B1 => B(21), B2 => n257, 
                           ZN => n45);
   U57 : AOI222_X1 port map( A1 => D(21), A2 => n269, B1 => E(21), B2 => n266, 
                           C1 => C(21), C2 => n263, ZN => n46);
   U58 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U59 : AOI22_X1 port map( A1 => A(19), A2 => n259, B1 => B(19), B2 => n256, 
                           ZN => n51);
   U60 : AOI222_X1 port map( A1 => D(19), A2 => n268, B1 => E(19), B2 => n265, 
                           C1 => C(19), C2 => n262, ZN => n52);
   U61 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U62 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U63 : AOI22_X1 port map( A1 => A(25), A2 => n260, B1 => B(25), B2 => n257, 
                           ZN => n37);
   U64 : AOI222_X1 port map( A1 => D(25), A2 => n269, B1 => E(25), B2 => n266, 
                           C1 => C(25), C2 => n263, ZN => n38);
   U65 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U66 : AOI22_X1 port map( A1 => A(29), A2 => n260, B1 => B(29), B2 => n257, 
                           ZN => n29);
   U67 : AOI222_X1 port map( A1 => D(29), A2 => n269, B1 => E(29), B2 => n266, 
                           C1 => C(29), C2 => n263, ZN => n30);
   U68 : INV_X1 port map( A => Sel(2), ZN => n74);
   U69 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U70 : AOI22_X1 port map( A1 => A(26), A2 => n260, B1 => B(26), B2 => n257, 
                           ZN => n35);
   U71 : AOI222_X1 port map( A1 => D(26), A2 => n269, B1 => E(26), B2 => n266, 
                           C1 => C(26), C2 => n263, ZN => n36);
   U72 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U73 : AOI22_X1 port map( A1 => A(6), A2 => n261, B1 => B(6), B2 => n258, ZN 
                           => n15);
   U74 : AOI222_X1 port map( A1 => D(6), A2 => n270, B1 => E(6), B2 => n267, C1
                           => C(6), C2 => n264, ZN => n16);
   U75 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U76 : AOI22_X1 port map( A1 => A(3), A2 => n261, B1 => B(3), B2 => n258, ZN 
                           => n21);
   U77 : AOI222_X1 port map( A1 => D(3), A2 => n270, B1 => E(3), B2 => n267, C1
                           => C(3), C2 => n264, ZN => n22);
   U78 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U79 : AOI22_X1 port map( A1 => A(7), A2 => n261, B1 => B(7), B2 => n258, ZN 
                           => n13);
   U80 : AOI222_X1 port map( A1 => D(7), A2 => n270, B1 => E(7), B2 => n267, C1
                           => C(7), C2 => n264, ZN => n14);
   U81 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U82 : AOI22_X1 port map( A1 => A(4), A2 => n261, B1 => B(4), B2 => n258, ZN 
                           => n19);
   U83 : AOI222_X1 port map( A1 => D(4), A2 => n270, B1 => E(4), B2 => n267, C1
                           => C(4), C2 => n264, ZN => n20);
   U84 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U85 : AOI22_X1 port map( A1 => A(8), A2 => n261, B1 => B(8), B2 => n258, ZN 
                           => n11);
   U86 : AOI222_X1 port map( A1 => D(8), A2 => n270, B1 => E(8), B2 => n267, C1
                           => C(8), C2 => n264, ZN => n12);
   U87 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U88 : AOI22_X1 port map( A1 => A(9), A2 => n261, B1 => B(9), B2 => n258, ZN 
                           => n4);
   U89 : AOI222_X1 port map( A1 => D(9), A2 => n270, B1 => E(9), B2 => n267, C1
                           => C(9), C2 => n264, ZN => n5);
   U90 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U91 : AOI22_X1 port map( A1 => A(5), A2 => n261, B1 => B(5), B2 => n258, ZN 
                           => n17);
   U92 : AOI222_X1 port map( A1 => D(5), A2 => n270, B1 => E(5), B2 => n267, C1
                           => C(5), C2 => n264, ZN => n18);
   U93 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U94 : AOI22_X1 port map( A1 => A(31), A2 => n261, B1 => B(31), B2 => n258, 
                           ZN => n23);
   U95 : AOI222_X1 port map( A1 => D(31), A2 => n270, B1 => E(31), B2 => n267, 
                           C1 => C(31), C2 => n264, ZN => n24);
   U96 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U97 : AOI22_X1 port map( A1 => A(2), A2 => n260, B1 => B(2), B2 => n257, ZN 
                           => n27);
   U98 : AOI222_X1 port map( A1 => D(2), A2 => n269, B1 => E(2), B2 => n266, C1
                           => C(2), C2 => n263, ZN => n28);
   U99 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U100 : AOI22_X1 port map( A1 => A(10), A2 => n259, B1 => B(10), B2 => n256, 
                           ZN => n69);
   U101 : AOI222_X1 port map( A1 => D(10), A2 => n268, B1 => E(10), B2 => n265,
                           C1 => C(10), C2 => n262, ZN => n70);
   U102 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U103 : AOI22_X1 port map( A1 => A(11), A2 => n259, B1 => B(11), B2 => n256, 
                           ZN => n67);
   U104 : AOI222_X1 port map( A1 => D(11), A2 => n268, B1 => E(11), B2 => n265,
                           C1 => C(11), C2 => n262, ZN => n68);
   U105 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U106 : AOI22_X1 port map( A1 => A(0), A2 => n259, B1 => B(0), B2 => n256, ZN
                           => n71);
   U107 : AOI222_X1 port map( A1 => D(0), A2 => n268, B1 => E(0), B2 => n265, 
                           C1 => C(0), C2 => n262, ZN => n72);
   U108 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U109 : AOI22_X1 port map( A1 => A(12), A2 => n259, B1 => B(12), B2 => n256, 
                           ZN => n65);
   U110 : AOI222_X1 port map( A1 => D(12), A2 => n268, B1 => E(12), B2 => n265,
                           C1 => C(12), C2 => n262, ZN => n66);
   U111 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U112 : AOI22_X1 port map( A1 => A(13), A2 => n259, B1 => B(13), B2 => n256, 
                           ZN => n63);
   U113 : AOI222_X1 port map( A1 => D(13), A2 => n268, B1 => E(13), B2 => n265,
                           C1 => C(13), C2 => n262, ZN => n64);
   U114 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U115 : AOI22_X1 port map( A1 => A(1), A2 => n259, B1 => B(1), B2 => n256, ZN
                           => n49);
   U116 : AOI222_X1 port map( A1 => D(1), A2 => n268, B1 => E(1), B2 => n265, 
                           C1 => C(1), C2 => n262, ZN => n50);
   U117 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U118 : AOI22_X1 port map( A1 => A(30), A2 => n260, B1 => B(30), B2 => n257, 
                           ZN => n25);
   U119 : AOI222_X1 port map( A1 => D(30), A2 => n269, B1 => E(30), B2 => n266,
                           C1 => C(30), C2 => n263, ZN => n26);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_2 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_2;

architecture SYN_behav of mux_N32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n269);
   U2 : BUF_X1 port map( A => n10, Z => n268);
   U3 : BUF_X1 port map( A => n10, Z => n270);
   U4 : BUF_X1 port map( A => n6, Z => n281);
   U5 : BUF_X1 port map( A => n6, Z => n280);
   U6 : BUF_X1 port map( A => n9, Z => n272);
   U7 : BUF_X1 port map( A => n9, Z => n271);
   U8 : BUF_X1 port map( A => n7, Z => n278);
   U9 : BUF_X1 port map( A => n7, Z => n277);
   U10 : BUF_X1 port map( A => n8, Z => n275);
   U11 : BUF_X1 port map( A => n8, Z => n274);
   U12 : BUF_X1 port map( A => n9, Z => n273);
   U13 : BUF_X1 port map( A => n7, Z => n279);
   U14 : BUF_X1 port map( A => n8, Z => n276);
   U15 : BUF_X1 port map( A => n6, Z => n282);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U24 : AOI22_X1 port map( A1 => A(26), A2 => n272, B1 => B(26), B2 => n269, 
                           ZN => n35);
   U25 : AOI222_X1 port map( A1 => D(26), A2 => n281, B1 => E(26), B2 => n278, 
                           C1 => C(26), C2 => n275, ZN => n36);
   U26 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U27 : AOI22_X1 port map( A1 => A(22), A2 => n272, B1 => B(22), B2 => n269, 
                           ZN => n43);
   U28 : AOI222_X1 port map( A1 => D(22), A2 => n281, B1 => E(22), B2 => n278, 
                           C1 => C(22), C2 => n275, ZN => n44);
   U29 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U30 : AOI22_X1 port map( A1 => A(28), A2 => n272, B1 => B(28), B2 => n269, 
                           ZN => n31);
   U31 : AOI222_X1 port map( A1 => D(28), A2 => n281, B1 => E(28), B2 => n278, 
                           C1 => C(28), C2 => n275, ZN => n32);
   U32 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U33 : AOI22_X1 port map( A1 => A(29), A2 => n272, B1 => B(29), B2 => n269, 
                           ZN => n29);
   U34 : AOI222_X1 port map( A1 => D(29), A2 => n281, B1 => E(29), B2 => n278, 
                           C1 => C(29), C2 => n275, ZN => n30);
   U35 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U36 : AOI22_X1 port map( A1 => A(30), A2 => n272, B1 => B(30), B2 => n269, 
                           ZN => n25);
   U37 : AOI222_X1 port map( A1 => D(30), A2 => n281, B1 => E(30), B2 => n278, 
                           C1 => C(30), C2 => n275, ZN => n26);
   U38 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U39 : AOI22_X1 port map( A1 => A(31), A2 => n273, B1 => B(31), B2 => n270, 
                           ZN => n23);
   U40 : AOI222_X1 port map( A1 => D(31), A2 => n282, B1 => E(31), B2 => n279, 
                           C1 => C(31), C2 => n276, ZN => n24);
   U41 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n271, B1 => B(16), B2 => n268, 
                           ZN => n57);
   U43 : AOI222_X1 port map( A1 => D(16), A2 => n280, B1 => E(16), B2 => n277, 
                           C1 => C(16), C2 => n274, ZN => n58);
   U44 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n272, B1 => B(20), B2 => n269, 
                           ZN => n47);
   U46 : AOI222_X1 port map( A1 => D(20), A2 => n281, B1 => E(20), B2 => n278, 
                           C1 => C(20), C2 => n275, ZN => n48);
   U47 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U48 : AOI22_X1 port map( A1 => A(14), A2 => n271, B1 => B(14), B2 => n268, 
                           ZN => n61);
   U49 : AOI222_X1 port map( A1 => D(14), A2 => n280, B1 => E(14), B2 => n277, 
                           C1 => C(14), C2 => n274, ZN => n62);
   U50 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U51 : AOI22_X1 port map( A1 => A(18), A2 => n271, B1 => B(18), B2 => n268, 
                           ZN => n53);
   U52 : AOI222_X1 port map( A1 => D(18), A2 => n280, B1 => E(18), B2 => n277, 
                           C1 => C(18), C2 => n274, ZN => n54);
   U53 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n272, B1 => B(25), B2 => n269, 
                           ZN => n37);
   U55 : AOI222_X1 port map( A1 => D(25), A2 => n281, B1 => E(25), B2 => n278, 
                           C1 => C(25), C2 => n275, ZN => n38);
   U56 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U57 : AOI22_X1 port map( A1 => A(21), A2 => n272, B1 => B(21), B2 => n269, 
                           ZN => n45);
   U58 : AOI222_X1 port map( A1 => D(21), A2 => n281, B1 => E(21), B2 => n278, 
                           C1 => C(21), C2 => n275, ZN => n46);
   U59 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U60 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U61 : AOI22_X1 port map( A1 => A(15), A2 => n271, B1 => B(15), B2 => n268, 
                           ZN => n59);
   U62 : AOI222_X1 port map( A1 => D(15), A2 => n280, B1 => E(15), B2 => n277, 
                           C1 => C(15), C2 => n274, ZN => n60);
   U63 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U64 : AOI22_X1 port map( A1 => A(19), A2 => n271, B1 => B(19), B2 => n268, 
                           ZN => n51);
   U65 : AOI222_X1 port map( A1 => D(19), A2 => n280, B1 => E(19), B2 => n277, 
                           C1 => C(19), C2 => n274, ZN => n52);
   U66 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U67 : AOI22_X1 port map( A1 => A(17), A2 => n271, B1 => B(17), B2 => n268, 
                           ZN => n55);
   U68 : AOI222_X1 port map( A1 => D(17), A2 => n280, B1 => E(17), B2 => n277, 
                           C1 => C(17), C2 => n274, ZN => n56);
   U69 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U70 : AOI22_X1 port map( A1 => A(12), A2 => n271, B1 => B(12), B2 => n268, 
                           ZN => n65);
   U71 : AOI222_X1 port map( A1 => D(12), A2 => n280, B1 => E(12), B2 => n277, 
                           C1 => C(12), C2 => n274, ZN => n66);
   U72 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U73 : AOI22_X1 port map( A1 => A(13), A2 => n271, B1 => B(13), B2 => n268, 
                           ZN => n63);
   U74 : AOI222_X1 port map( A1 => D(13), A2 => n280, B1 => E(13), B2 => n277, 
                           C1 => C(13), C2 => n274, ZN => n64);
   U75 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U76 : AOI22_X1 port map( A1 => A(23), A2 => n272, B1 => B(23), B2 => n269, 
                           ZN => n41);
   U77 : AOI222_X1 port map( A1 => D(23), A2 => n281, B1 => E(23), B2 => n278, 
                           C1 => C(23), C2 => n275, ZN => n42);
   U78 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U79 : AOI22_X1 port map( A1 => A(27), A2 => n272, B1 => B(27), B2 => n269, 
                           ZN => n33);
   U80 : AOI222_X1 port map( A1 => D(27), A2 => n281, B1 => E(27), B2 => n278, 
                           C1 => C(27), C2 => n275, ZN => n34);
   U81 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U82 : AOI22_X1 port map( A1 => A(24), A2 => n272, B1 => B(24), B2 => n269, 
                           ZN => n39);
   U83 : AOI222_X1 port map( A1 => D(24), A2 => n281, B1 => E(24), B2 => n278, 
                           C1 => C(24), C2 => n275, ZN => n40);
   U84 : INV_X1 port map( A => Sel(1), ZN => n75);
   U85 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U86 : AOI22_X1 port map( A1 => A(6), A2 => n273, B1 => B(6), B2 => n270, ZN 
                           => n15);
   U87 : AOI222_X1 port map( A1 => D(6), A2 => n282, B1 => E(6), B2 => n279, C1
                           => C(6), C2 => n276, ZN => n16);
   U88 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U89 : AOI22_X1 port map( A1 => A(3), A2 => n273, B1 => B(3), B2 => n270, ZN 
                           => n21);
   U90 : AOI222_X1 port map( A1 => D(3), A2 => n282, B1 => E(3), B2 => n279, C1
                           => C(3), C2 => n276, ZN => n22);
   U91 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U92 : AOI22_X1 port map( A1 => A(7), A2 => n273, B1 => B(7), B2 => n270, ZN 
                           => n13);
   U93 : AOI222_X1 port map( A1 => D(7), A2 => n282, B1 => E(7), B2 => n279, C1
                           => C(7), C2 => n276, ZN => n14);
   U94 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U95 : AOI22_X1 port map( A1 => A(4), A2 => n273, B1 => B(4), B2 => n270, ZN 
                           => n19);
   U96 : AOI222_X1 port map( A1 => D(4), A2 => n282, B1 => E(4), B2 => n279, C1
                           => C(4), C2 => n276, ZN => n20);
   U97 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U98 : AOI22_X1 port map( A1 => A(8), A2 => n273, B1 => B(8), B2 => n270, ZN 
                           => n11);
   U99 : AOI222_X1 port map( A1 => D(8), A2 => n282, B1 => E(8), B2 => n279, C1
                           => C(8), C2 => n276, ZN => n12);
   U100 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U101 : AOI22_X1 port map( A1 => A(9), A2 => n273, B1 => B(9), B2 => n270, ZN
                           => n4);
   U102 : AOI222_X1 port map( A1 => D(9), A2 => n282, B1 => E(9), B2 => n279, 
                           C1 => C(9), C2 => n276, ZN => n5);
   U103 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U104 : AOI22_X1 port map( A1 => A(5), A2 => n273, B1 => B(5), B2 => n270, ZN
                           => n17);
   U105 : AOI222_X1 port map( A1 => D(5), A2 => n282, B1 => E(5), B2 => n279, 
                           C1 => C(5), C2 => n276, ZN => n18);
   U106 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U107 : AOI22_X1 port map( A1 => A(2), A2 => n272, B1 => B(2), B2 => n269, ZN
                           => n27);
   U108 : AOI222_X1 port map( A1 => D(2), A2 => n281, B1 => E(2), B2 => n278, 
                           C1 => C(2), C2 => n275, ZN => n28);
   U109 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U110 : AOI22_X1 port map( A1 => A(10), A2 => n271, B1 => B(10), B2 => n268, 
                           ZN => n69);
   U111 : AOI222_X1 port map( A1 => D(10), A2 => n280, B1 => E(10), B2 => n277,
                           C1 => C(10), C2 => n274, ZN => n70);
   U112 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U113 : AOI22_X1 port map( A1 => A(11), A2 => n271, B1 => B(11), B2 => n268, 
                           ZN => n67);
   U114 : AOI222_X1 port map( A1 => D(11), A2 => n280, B1 => E(11), B2 => n277,
                           C1 => C(11), C2 => n274, ZN => n68);
   U115 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U116 : AOI22_X1 port map( A1 => A(0), A2 => n271, B1 => B(0), B2 => n268, ZN
                           => n71);
   U117 : AOI222_X1 port map( A1 => D(0), A2 => n280, B1 => E(0), B2 => n277, 
                           C1 => C(0), C2 => n274, ZN => n72);
   U118 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U119 : AOI22_X1 port map( A1 => A(1), A2 => n271, B1 => B(1), B2 => n268, ZN
                           => n49);
   U120 : AOI222_X1 port map( A1 => D(1), A2 => n280, B1 => E(1), B2 => n277, 
                           C1 => C(1), C2 => n274, ZN => n50);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_3 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_3;

architecture SYN_behav of mux_N32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n265);
   U2 : BUF_X1 port map( A => n10, Z => n266);
   U3 : BUF_X1 port map( A => n10, Z => n267);
   U4 : BUF_X1 port map( A => n6, Z => n277);
   U5 : BUF_X1 port map( A => n6, Z => n278);
   U6 : BUF_X1 port map( A => n9, Z => n268);
   U7 : BUF_X1 port map( A => n9, Z => n269);
   U8 : BUF_X1 port map( A => n7, Z => n274);
   U9 : BUF_X1 port map( A => n7, Z => n275);
   U10 : BUF_X1 port map( A => n8, Z => n271);
   U11 : BUF_X1 port map( A => n8, Z => n272);
   U12 : BUF_X1 port map( A => n9, Z => n270);
   U13 : BUF_X1 port map( A => n7, Z => n276);
   U14 : BUF_X1 port map( A => n8, Z => n273);
   U15 : BUF_X1 port map( A => n6, Z => n279);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U24 : AOI22_X1 port map( A1 => A(24), A2 => n269, B1 => B(24), B2 => n266, 
                           ZN => n39);
   U25 : AOI222_X1 port map( A1 => D(24), A2 => n278, B1 => E(24), B2 => n275, 
                           C1 => C(24), C2 => n272, ZN => n40);
   U26 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U27 : AOI22_X1 port map( A1 => A(20), A2 => n269, B1 => B(20), B2 => n266, 
                           ZN => n47);
   U28 : AOI222_X1 port map( A1 => D(20), A2 => n278, B1 => E(20), B2 => n275, 
                           C1 => C(20), C2 => n272, ZN => n48);
   U29 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U30 : AOI22_X1 port map( A1 => A(14), A2 => n268, B1 => B(14), B2 => n265, 
                           ZN => n61);
   U31 : AOI222_X1 port map( A1 => D(14), A2 => n277, B1 => E(14), B2 => n274, 
                           C1 => C(14), C2 => n271, ZN => n62);
   U32 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U33 : AOI22_X1 port map( A1 => A(18), A2 => n268, B1 => B(18), B2 => n265, 
                           ZN => n53);
   U34 : AOI222_X1 port map( A1 => D(18), A2 => n277, B1 => E(18), B2 => n274, 
                           C1 => C(18), C2 => n271, ZN => n54);
   U35 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U36 : AOI22_X1 port map( A1 => A(12), A2 => n268, B1 => B(12), B2 => n265, 
                           ZN => n65);
   U37 : AOI222_X1 port map( A1 => D(12), A2 => n277, B1 => E(12), B2 => n274, 
                           C1 => C(12), C2 => n271, ZN => n66);
   U38 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U39 : AOI22_X1 port map( A1 => A(16), A2 => n268, B1 => B(16), B2 => n265, 
                           ZN => n57);
   U40 : AOI222_X1 port map( A1 => D(16), A2 => n277, B1 => E(16), B2 => n274, 
                           C1 => C(16), C2 => n271, ZN => n58);
   U41 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U42 : AOI22_X1 port map( A1 => A(23), A2 => n269, B1 => B(23), B2 => n266, 
                           ZN => n41);
   U43 : AOI222_X1 port map( A1 => D(23), A2 => n278, B1 => E(23), B2 => n275, 
                           C1 => C(23), C2 => n272, ZN => n42);
   U44 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U45 : AOI22_X1 port map( A1 => A(19), A2 => n268, B1 => B(19), B2 => n265, 
                           ZN => n51);
   U46 : AOI222_X1 port map( A1 => D(19), A2 => n277, B1 => E(19), B2 => n274, 
                           C1 => C(19), C2 => n271, ZN => n52);
   U47 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U48 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U49 : AOI22_X1 port map( A1 => A(13), A2 => n268, B1 => B(13), B2 => n265, 
                           ZN => n63);
   U50 : AOI222_X1 port map( A1 => D(13), A2 => n277, B1 => E(13), B2 => n274, 
                           C1 => C(13), C2 => n271, ZN => n64);
   U51 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U52 : AOI22_X1 port map( A1 => A(17), A2 => n268, B1 => B(17), B2 => n265, 
                           ZN => n55);
   U53 : AOI222_X1 port map( A1 => D(17), A2 => n277, B1 => E(17), B2 => n274, 
                           C1 => C(17), C2 => n271, ZN => n56);
   U54 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U55 : AOI22_X1 port map( A1 => A(15), A2 => n268, B1 => B(15), B2 => n265, 
                           ZN => n59);
   U56 : AOI222_X1 port map( A1 => D(15), A2 => n277, B1 => E(15), B2 => n274, 
                           C1 => C(15), C2 => n271, ZN => n60);
   U57 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U58 : AOI22_X1 port map( A1 => A(10), A2 => n268, B1 => B(10), B2 => n265, 
                           ZN => n69);
   U59 : AOI222_X1 port map( A1 => D(10), A2 => n277, B1 => E(10), B2 => n274, 
                           C1 => C(10), C2 => n271, ZN => n70);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U61 : AOI22_X1 port map( A1 => A(11), A2 => n268, B1 => B(11), B2 => n265, 
                           ZN => n67);
   U62 : AOI222_X1 port map( A1 => D(11), A2 => n277, B1 => E(11), B2 => n274, 
                           C1 => C(11), C2 => n271, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U64 : AOI22_X1 port map( A1 => A(21), A2 => n269, B1 => B(21), B2 => n266, 
                           ZN => n45);
   U65 : AOI222_X1 port map( A1 => D(21), A2 => n278, B1 => E(21), B2 => n275, 
                           C1 => C(21), C2 => n272, ZN => n46);
   U66 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U67 : AOI22_X1 port map( A1 => A(25), A2 => n269, B1 => B(25), B2 => n266, 
                           ZN => n37);
   U68 : AOI222_X1 port map( A1 => D(25), A2 => n278, B1 => E(25), B2 => n275, 
                           C1 => C(25), C2 => n272, ZN => n38);
   U69 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U70 : AOI22_X1 port map( A1 => A(26), A2 => n269, B1 => B(26), B2 => n266, 
                           ZN => n35);
   U71 : AOI222_X1 port map( A1 => D(26), A2 => n278, B1 => E(26), B2 => n275, 
                           C1 => C(26), C2 => n272, ZN => n36);
   U72 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U73 : AOI22_X1 port map( A1 => A(27), A2 => n269, B1 => B(27), B2 => n266, 
                           ZN => n33);
   U74 : AOI222_X1 port map( A1 => D(27), A2 => n278, B1 => E(27), B2 => n275, 
                           C1 => C(27), C2 => n272, ZN => n34);
   U75 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U76 : AOI22_X1 port map( A1 => A(28), A2 => n269, B1 => B(28), B2 => n266, 
                           ZN => n31);
   U77 : AOI222_X1 port map( A1 => D(28), A2 => n278, B1 => E(28), B2 => n275, 
                           C1 => C(28), C2 => n272, ZN => n32);
   U78 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U79 : AOI22_X1 port map( A1 => A(29), A2 => n269, B1 => B(29), B2 => n266, 
                           ZN => n29);
   U80 : AOI222_X1 port map( A1 => D(29), A2 => n278, B1 => E(29), B2 => n275, 
                           C1 => C(29), C2 => n272, ZN => n30);
   U81 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U82 : AOI22_X1 port map( A1 => A(30), A2 => n269, B1 => B(30), B2 => n266, 
                           ZN => n25);
   U83 : AOI222_X1 port map( A1 => D(30), A2 => n278, B1 => E(30), B2 => n275, 
                           C1 => C(30), C2 => n272, ZN => n26);
   U84 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U85 : AOI22_X1 port map( A1 => A(31), A2 => n270, B1 => B(31), B2 => n267, 
                           ZN => n23);
   U86 : AOI222_X1 port map( A1 => D(31), A2 => n279, B1 => E(31), B2 => n276, 
                           C1 => C(31), C2 => n273, ZN => n24);
   U87 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U88 : AOI22_X1 port map( A1 => A(22), A2 => n269, B1 => B(22), B2 => n266, 
                           ZN => n43);
   U89 : AOI222_X1 port map( A1 => D(22), A2 => n278, B1 => E(22), B2 => n275, 
                           C1 => C(22), C2 => n272, ZN => n44);
   U90 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U91 : AOI22_X1 port map( A1 => A(9), A2 => n270, B1 => B(9), B2 => n267, ZN 
                           => n4);
   U92 : AOI222_X1 port map( A1 => D(9), A2 => n279, B1 => E(9), B2 => n276, C1
                           => C(9), C2 => n273, ZN => n5);
   U93 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U94 : AOI22_X1 port map( A1 => A(5), A2 => n270, B1 => B(5), B2 => n267, ZN 
                           => n17);
   U95 : AOI222_X1 port map( A1 => D(5), A2 => n279, B1 => E(5), B2 => n276, C1
                           => C(5), C2 => n273, ZN => n18);
   U96 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U97 : AOI22_X1 port map( A1 => A(6), A2 => n270, B1 => B(6), B2 => n267, ZN 
                           => n15);
   U98 : AOI222_X1 port map( A1 => D(6), A2 => n279, B1 => E(6), B2 => n276, C1
                           => C(6), C2 => n273, ZN => n16);
   U99 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U100 : AOI22_X1 port map( A1 => A(3), A2 => n270, B1 => B(3), B2 => n267, ZN
                           => n21);
   U101 : AOI222_X1 port map( A1 => D(3), A2 => n279, B1 => E(3), B2 => n276, 
                           C1 => C(3), C2 => n273, ZN => n22);
   U102 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U103 : AOI22_X1 port map( A1 => A(7), A2 => n270, B1 => B(7), B2 => n267, ZN
                           => n13);
   U104 : AOI222_X1 port map( A1 => D(7), A2 => n279, B1 => E(7), B2 => n276, 
                           C1 => C(7), C2 => n273, ZN => n14);
   U105 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U106 : AOI22_X1 port map( A1 => A(4), A2 => n270, B1 => B(4), B2 => n267, ZN
                           => n19);
   U107 : AOI222_X1 port map( A1 => D(4), A2 => n279, B1 => E(4), B2 => n276, 
                           C1 => C(4), C2 => n273, ZN => n20);
   U108 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U109 : AOI22_X1 port map( A1 => A(8), A2 => n270, B1 => B(8), B2 => n267, ZN
                           => n11);
   U110 : AOI222_X1 port map( A1 => D(8), A2 => n279, B1 => E(8), B2 => n276, 
                           C1 => C(8), C2 => n273, ZN => n12);
   U111 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U112 : AOI22_X1 port map( A1 => A(1), A2 => n268, B1 => B(1), B2 => n265, ZN
                           => n49);
   U113 : AOI222_X1 port map( A1 => D(1), A2 => n277, B1 => E(1), B2 => n274, 
                           C1 => C(1), C2 => n271, ZN => n50);
   U114 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U115 : AOI22_X1 port map( A1 => A(2), A2 => n269, B1 => B(2), B2 => n266, ZN
                           => n27);
   U116 : AOI222_X1 port map( A1 => D(2), A2 => n278, B1 => E(2), B2 => n275, 
                           C1 => C(2), C2 => n272, ZN => n28);
   U117 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U118 : AOI22_X1 port map( A1 => A(0), A2 => n268, B1 => B(0), B2 => n265, ZN
                           => n71);
   U119 : AOI222_X1 port map( A1 => D(0), A2 => n277, B1 => E(0), B2 => n274, 
                           C1 => C(0), C2 => n271, ZN => n72);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_4 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_4;

architecture SYN_behav of mux_N32_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n280);
   U2 : BUF_X1 port map( A => n10, Z => n281);
   U3 : BUF_X1 port map( A => n10, Z => n282);
   U4 : BUF_X1 port map( A => n6, Z => n292);
   U5 : BUF_X1 port map( A => n6, Z => n293);
   U6 : BUF_X1 port map( A => n9, Z => n283);
   U7 : BUF_X1 port map( A => n9, Z => n284);
   U8 : BUF_X1 port map( A => n7, Z => n289);
   U9 : BUF_X1 port map( A => n7, Z => n290);
   U10 : BUF_X1 port map( A => n8, Z => n286);
   U11 : BUF_X1 port map( A => n8, Z => n287);
   U12 : BUF_X1 port map( A => n9, Z => n285);
   U13 : BUF_X1 port map( A => n7, Z => n291);
   U14 : BUF_X1 port map( A => n8, Z => n288);
   U15 : BUF_X1 port map( A => n6, Z => n294);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U24 : AOI22_X1 port map( A1 => A(22), A2 => n284, B1 => B(22), B2 => n281, 
                           ZN => n43);
   U25 : AOI222_X1 port map( A1 => D(22), A2 => n293, B1 => E(22), B2 => n290, 
                           C1 => C(22), C2 => n287, ZN => n44);
   U26 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U27 : AOI22_X1 port map( A1 => A(8), A2 => n285, B1 => B(8), B2 => n282, ZN 
                           => n11);
   U28 : AOI222_X1 port map( A1 => D(8), A2 => n294, B1 => E(8), B2 => n291, C1
                           => C(8), C2 => n288, ZN => n12);
   U29 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U30 : AOI22_X1 port map( A1 => A(18), A2 => n283, B1 => B(18), B2 => n280, 
                           ZN => n53);
   U31 : AOI222_X1 port map( A1 => D(18), A2 => n292, B1 => E(18), B2 => n289, 
                           C1 => C(18), C2 => n286, ZN => n54);
   U32 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U33 : AOI22_X1 port map( A1 => A(25), A2 => n284, B1 => B(25), B2 => n281, 
                           ZN => n37);
   U34 : AOI222_X1 port map( A1 => D(25), A2 => n293, B1 => E(25), B2 => n290, 
                           C1 => C(25), C2 => n287, ZN => n38);
   U35 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U36 : AOI22_X1 port map( A1 => A(26), A2 => n284, B1 => B(26), B2 => n281, 
                           ZN => n35);
   U37 : AOI222_X1 port map( A1 => D(26), A2 => n293, B1 => E(26), B2 => n290, 
                           C1 => C(26), C2 => n287, ZN => n36);
   U38 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U39 : AOI22_X1 port map( A1 => A(27), A2 => n284, B1 => B(27), B2 => n281, 
                           ZN => n33);
   U40 : AOI222_X1 port map( A1 => D(27), A2 => n293, B1 => E(27), B2 => n290, 
                           C1 => C(27), C2 => n287, ZN => n34);
   U41 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U42 : AOI22_X1 port map( A1 => A(28), A2 => n284, B1 => B(28), B2 => n281, 
                           ZN => n31);
   U43 : AOI222_X1 port map( A1 => D(28), A2 => n293, B1 => E(28), B2 => n290, 
                           C1 => C(28), C2 => n287, ZN => n32);
   U44 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U45 : AOI22_X1 port map( A1 => A(24), A2 => n284, B1 => B(24), B2 => n281, 
                           ZN => n39);
   U46 : AOI222_X1 port map( A1 => D(24), A2 => n293, B1 => E(24), B2 => n290, 
                           C1 => C(24), C2 => n287, ZN => n40);
   U47 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U48 : AOI22_X1 port map( A1 => A(29), A2 => n284, B1 => B(29), B2 => n281, 
                           ZN => n29);
   U49 : AOI222_X1 port map( A1 => D(29), A2 => n293, B1 => E(29), B2 => n290, 
                           C1 => C(29), C2 => n287, ZN => n30);
   U50 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U51 : AOI22_X1 port map( A1 => A(30), A2 => n284, B1 => B(30), B2 => n281, 
                           ZN => n25);
   U52 : AOI222_X1 port map( A1 => D(30), A2 => n293, B1 => E(30), B2 => n290, 
                           C1 => C(30), C2 => n287, ZN => n26);
   U53 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U54 : AOI22_X1 port map( A1 => A(31), A2 => n285, B1 => B(31), B2 => n282, 
                           ZN => n23);
   U55 : AOI222_X1 port map( A1 => D(31), A2 => n294, B1 => E(31), B2 => n291, 
                           C1 => C(31), C2 => n288, ZN => n24);
   U56 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U57 : AOI22_X1 port map( A1 => A(12), A2 => n283, B1 => B(12), B2 => n280, 
                           ZN => n65);
   U58 : AOI222_X1 port map( A1 => D(12), A2 => n292, B1 => E(12), B2 => n289, 
                           C1 => C(12), C2 => n286, ZN => n66);
   U59 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U60 : AOI22_X1 port map( A1 => A(9), A2 => n285, B1 => B(9), B2 => n282, ZN 
                           => n4);
   U61 : AOI222_X1 port map( A1 => D(9), A2 => n294, B1 => E(9), B2 => n291, C1
                           => C(9), C2 => n288, ZN => n5);
   U62 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U63 : AOI22_X1 port map( A1 => A(16), A2 => n283, B1 => B(16), B2 => n280, 
                           ZN => n57);
   U64 : AOI222_X1 port map( A1 => D(16), A2 => n292, B1 => E(16), B2 => n289, 
                           C1 => C(16), C2 => n286, ZN => n58);
   U65 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U66 : AOI22_X1 port map( A1 => A(10), A2 => n283, B1 => B(10), B2 => n280, 
                           ZN => n69);
   U67 : AOI222_X1 port map( A1 => D(10), A2 => n292, B1 => E(10), B2 => n289, 
                           C1 => C(10), C2 => n286, ZN => n70);
   U68 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U69 : AOI22_X1 port map( A1 => A(14), A2 => n283, B1 => B(14), B2 => n280, 
                           ZN => n61);
   U70 : AOI222_X1 port map( A1 => D(14), A2 => n292, B1 => E(14), B2 => n289, 
                           C1 => C(14), C2 => n286, ZN => n62);
   U71 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U72 : AOI22_X1 port map( A1 => A(21), A2 => n284, B1 => B(21), B2 => n281, 
                           ZN => n45);
   U73 : AOI222_X1 port map( A1 => D(21), A2 => n293, B1 => E(21), B2 => n290, 
                           C1 => C(21), C2 => n287, ZN => n46);
   U74 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U75 : AOI22_X1 port map( A1 => A(17), A2 => n283, B1 => B(17), B2 => n280, 
                           ZN => n55);
   U76 : AOI222_X1 port map( A1 => D(17), A2 => n292, B1 => E(17), B2 => n289, 
                           C1 => C(17), C2 => n286, ZN => n56);
   U77 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U78 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U79 : AOI22_X1 port map( A1 => A(11), A2 => n283, B1 => B(11), B2 => n280, 
                           ZN => n67);
   U80 : AOI222_X1 port map( A1 => D(11), A2 => n292, B1 => E(11), B2 => n289, 
                           C1 => C(11), C2 => n286, ZN => n68);
   U81 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U82 : AOI22_X1 port map( A1 => A(15), A2 => n283, B1 => B(15), B2 => n280, 
                           ZN => n59);
   U83 : AOI222_X1 port map( A1 => D(15), A2 => n292, B1 => E(15), B2 => n289, 
                           C1 => C(15), C2 => n286, ZN => n60);
   U84 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U85 : AOI22_X1 port map( A1 => A(13), A2 => n283, B1 => B(13), B2 => n280, 
                           ZN => n63);
   U86 : AOI222_X1 port map( A1 => D(13), A2 => n292, B1 => E(13), B2 => n289, 
                           C1 => C(13), C2 => n286, ZN => n64);
   U87 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U88 : AOI22_X1 port map( A1 => A(20), A2 => n284, B1 => B(20), B2 => n281, 
                           ZN => n47);
   U89 : AOI222_X1 port map( A1 => D(20), A2 => n293, B1 => E(20), B2 => n290, 
                           C1 => C(20), C2 => n287, ZN => n48);
   U90 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U91 : AOI22_X1 port map( A1 => A(19), A2 => n283, B1 => B(19), B2 => n280, 
                           ZN => n51);
   U92 : AOI222_X1 port map( A1 => D(19), A2 => n292, B1 => E(19), B2 => n289, 
                           C1 => C(19), C2 => n286, ZN => n52);
   U93 : INV_X1 port map( A => Sel(1), ZN => n75);
   U94 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U95 : AOI22_X1 port map( A1 => A(5), A2 => n285, B1 => B(5), B2 => n282, ZN 
                           => n17);
   U96 : AOI222_X1 port map( A1 => D(5), A2 => n294, B1 => E(5), B2 => n291, C1
                           => C(5), C2 => n288, ZN => n18);
   U97 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U98 : AOI22_X1 port map( A1 => A(6), A2 => n285, B1 => B(6), B2 => n282, ZN 
                           => n15);
   U99 : AOI222_X1 port map( A1 => D(6), A2 => n294, B1 => E(6), B2 => n291, C1
                           => C(6), C2 => n288, ZN => n16);
   U100 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U101 : AOI22_X1 port map( A1 => A(3), A2 => n285, B1 => B(3), B2 => n282, ZN
                           => n21);
   U102 : AOI222_X1 port map( A1 => D(3), A2 => n294, B1 => E(3), B2 => n291, 
                           C1 => C(3), C2 => n288, ZN => n22);
   U103 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U104 : AOI22_X1 port map( A1 => A(7), A2 => n285, B1 => B(7), B2 => n282, ZN
                           => n13);
   U105 : AOI222_X1 port map( A1 => D(7), A2 => n294, B1 => E(7), B2 => n291, 
                           C1 => C(7), C2 => n288, ZN => n14);
   U106 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U107 : AOI22_X1 port map( A1 => A(4), A2 => n285, B1 => B(4), B2 => n282, ZN
                           => n19);
   U108 : AOI222_X1 port map( A1 => D(4), A2 => n294, B1 => E(4), B2 => n291, 
                           C1 => C(4), C2 => n288, ZN => n20);
   U109 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U110 : AOI22_X1 port map( A1 => A(1), A2 => n283, B1 => B(1), B2 => n280, ZN
                           => n49);
   U111 : AOI222_X1 port map( A1 => D(1), A2 => n292, B1 => E(1), B2 => n289, 
                           C1 => C(1), C2 => n286, ZN => n50);
   U112 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U113 : AOI22_X1 port map( A1 => A(2), A2 => n284, B1 => B(2), B2 => n281, ZN
                           => n27);
   U114 : AOI222_X1 port map( A1 => D(2), A2 => n293, B1 => E(2), B2 => n290, 
                           C1 => C(2), C2 => n287, ZN => n28);
   U115 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U116 : AOI22_X1 port map( A1 => A(23), A2 => n284, B1 => B(23), B2 => n281, 
                           ZN => n41);
   U117 : AOI222_X1 port map( A1 => D(23), A2 => n293, B1 => E(23), B2 => n290,
                           C1 => C(23), C2 => n287, ZN => n42);
   U118 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U119 : AOI22_X1 port map( A1 => A(0), A2 => n283, B1 => B(0), B2 => n280, ZN
                           => n71);
   U120 : AOI222_X1 port map( A1 => D(0), A2 => n292, B1 => E(0), B2 => n289, 
                           C1 => C(0), C2 => n286, ZN => n72);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_5 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_5;

architecture SYN_behav of mux_N32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n274);
   U2 : BUF_X1 port map( A => n10, Z => n275);
   U3 : BUF_X1 port map( A => n10, Z => n276);
   U4 : BUF_X1 port map( A => n6, Z => n286);
   U5 : BUF_X1 port map( A => n6, Z => n287);
   U6 : BUF_X1 port map( A => n9, Z => n277);
   U7 : BUF_X1 port map( A => n9, Z => n278);
   U8 : BUF_X1 port map( A => n7, Z => n283);
   U9 : BUF_X1 port map( A => n7, Z => n284);
   U10 : BUF_X1 port map( A => n8, Z => n280);
   U11 : BUF_X1 port map( A => n8, Z => n281);
   U12 : BUF_X1 port map( A => n9, Z => n279);
   U13 : BUF_X1 port map( A => n7, Z => n285);
   U14 : BUF_X1 port map( A => n8, Z => n282);
   U15 : BUF_X1 port map( A => n6, Z => n288);
   U16 : AND2_X1 port map( A1 => n74, A2 => n73, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n73, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n73, ZN => n8);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n74);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n73);
   U23 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U24 : AOI22_X1 port map( A1 => A(20), A2 => n278, B1 => B(20), B2 => n275, 
                           ZN => n47);
   U25 : AOI222_X1 port map( A1 => D(20), A2 => n287, B1 => C(20), B2 => n284, 
                           C1 => E(20), C2 => n281, ZN => n48);
   U26 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U27 : AOI22_X1 port map( A1 => A(16), A2 => n277, B1 => B(16), B2 => n274, 
                           ZN => n57);
   U28 : AOI222_X1 port map( A1 => D(16), A2 => n286, B1 => C(16), B2 => n283, 
                           C1 => E(16), C2 => n280, ZN => n58);
   U29 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n277, B1 => B(10), B2 => n274, 
                           ZN => n69);
   U31 : AOI222_X1 port map( A1 => D(10), A2 => n286, B1 => C(10), B2 => n283, 
                           C1 => E(10), C2 => n280, ZN => n70);
   U32 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n277, B1 => B(14), B2 => n274, 
                           ZN => n61);
   U34 : AOI222_X1 port map( A1 => D(14), A2 => n286, B1 => C(14), B2 => n283, 
                           C1 => E(14), C2 => n280, ZN => n62);
   U35 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n279, B1 => B(8), B2 => n276, ZN 
                           => n11);
   U37 : AOI222_X1 port map( A1 => D(8), A2 => n288, B1 => C(8), B2 => n285, C1
                           => E(8), C2 => n282, ZN => n12);
   U38 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U39 : AOI22_X1 port map( A1 => A(12), A2 => n277, B1 => B(12), B2 => n274, 
                           ZN => n65);
   U40 : AOI222_X1 port map( A1 => D(12), A2 => n286, B1 => C(12), B2 => n283, 
                           C1 => E(12), C2 => n280, ZN => n66);
   U41 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U42 : AOI22_X1 port map( A1 => A(19), A2 => n277, B1 => B(19), B2 => n274, 
                           ZN => n51);
   U43 : AOI222_X1 port map( A1 => D(19), A2 => n286, B1 => C(19), B2 => n283, 
                           C1 => E(19), C2 => n280, ZN => n52);
   U44 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U45 : AOI22_X1 port map( A1 => A(15), A2 => n277, B1 => B(15), B2 => n274, 
                           ZN => n59);
   U46 : AOI222_X1 port map( A1 => D(15), A2 => n286, B1 => C(15), B2 => n283, 
                           C1 => E(15), C2 => n280, ZN => n60);
   U47 : AND2_X1 port map( A1 => Sel(2), A2 => n74, ZN => n7);
   U48 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U49 : AOI22_X1 port map( A1 => A(9), A2 => n279, B1 => B(9), B2 => n276, ZN 
                           => n4);
   U50 : AOI222_X1 port map( A1 => D(9), A2 => n288, B1 => C(9), B2 => n285, C1
                           => E(9), C2 => n282, ZN => n5);
   U51 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U52 : AOI22_X1 port map( A1 => A(13), A2 => n277, B1 => B(13), B2 => n274, 
                           ZN => n63);
   U53 : AOI222_X1 port map( A1 => D(13), A2 => n286, B1 => C(13), B2 => n283, 
                           C1 => E(13), C2 => n280, ZN => n64);
   U54 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U55 : AOI22_X1 port map( A1 => A(7), A2 => n279, B1 => B(7), B2 => n276, ZN 
                           => n13);
   U56 : AOI222_X1 port map( A1 => D(7), A2 => n288, B1 => C(7), B2 => n285, C1
                           => E(7), C2 => n282, ZN => n14);
   U57 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U58 : AOI22_X1 port map( A1 => A(17), A2 => n277, B1 => B(17), B2 => n274, 
                           ZN => n55);
   U59 : AOI222_X1 port map( A1 => D(17), A2 => n286, B1 => C(17), B2 => n283, 
                           C1 => E(17), C2 => n280, ZN => n56);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U61 : AOI22_X1 port map( A1 => A(11), A2 => n277, B1 => B(11), B2 => n274, 
                           ZN => n67);
   U62 : AOI222_X1 port map( A1 => D(11), A2 => n286, B1 => C(11), B2 => n283, 
                           C1 => E(11), C2 => n280, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U64 : AOI22_X1 port map( A1 => A(6), A2 => n279, B1 => B(6), B2 => n276, ZN 
                           => n15);
   U65 : AOI222_X1 port map( A1 => D(6), A2 => n288, B1 => C(6), B2 => n285, C1
                           => E(6), C2 => n282, ZN => n16);
   U66 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U67 : AOI22_X1 port map( A1 => A(18), A2 => n277, B1 => B(18), B2 => n274, 
                           ZN => n53);
   U68 : AOI222_X1 port map( A1 => D(18), A2 => n286, B1 => C(18), B2 => n283, 
                           C1 => E(18), C2 => n280, ZN => n54);
   U69 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U70 : AOI22_X1 port map( A1 => A(21), A2 => n278, B1 => B(21), B2 => n275, 
                           ZN => n45);
   U71 : AOI222_X1 port map( A1 => D(21), A2 => n287, B1 => C(21), B2 => n284, 
                           C1 => E(21), C2 => n281, ZN => n46);
   U72 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U73 : AOI22_X1 port map( A1 => A(5), A2 => n279, B1 => B(5), B2 => n276, ZN 
                           => n17);
   U74 : AOI222_X1 port map( A1 => D(5), A2 => n288, B1 => C(5), B2 => n285, C1
                           => E(5), C2 => n282, ZN => n18);
   U75 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U76 : AOI22_X1 port map( A1 => A(3), A2 => n279, B1 => B(3), B2 => n276, ZN 
                           => n21);
   U77 : AOI222_X1 port map( A1 => D(3), A2 => n288, B1 => C(3), B2 => n285, C1
                           => E(3), C2 => n282, ZN => n22);
   U78 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U79 : AOI22_X1 port map( A1 => A(4), A2 => n279, B1 => B(4), B2 => n276, ZN 
                           => n19);
   U80 : AOI222_X1 port map( A1 => D(4), A2 => n288, B1 => C(4), B2 => n285, C1
                           => E(4), C2 => n282, ZN => n20);
   U81 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U82 : AOI22_X1 port map( A1 => A(31), A2 => n279, B1 => B(31), B2 => n276, 
                           ZN => n23);
   U83 : AOI222_X1 port map( A1 => D(31), A2 => n288, B1 => C(31), B2 => n285, 
                           C1 => E(31), C2 => n282, ZN => n24);
   U84 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U85 : AOI22_X1 port map( A1 => A(1), A2 => n277, B1 => B(1), B2 => n274, ZN 
                           => n49);
   U86 : AOI222_X1 port map( A1 => D(1), A2 => n286, B1 => C(1), B2 => n283, C1
                           => E(1), C2 => n280, ZN => n50);
   U87 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U88 : AOI22_X1 port map( A1 => A(25), A2 => n278, B1 => B(25), B2 => n275, 
                           ZN => n37);
   U89 : AOI222_X1 port map( A1 => D(25), A2 => n287, B1 => C(25), B2 => n284, 
                           C1 => E(25), C2 => n281, ZN => n38);
   U90 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U91 : AOI22_X1 port map( A1 => A(2), A2 => n278, B1 => B(2), B2 => n275, ZN 
                           => n27);
   U92 : AOI222_X1 port map( A1 => D(2), A2 => n287, B1 => C(2), B2 => n284, C1
                           => E(2), C2 => n281, ZN => n28);
   U93 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U94 : AOI22_X1 port map( A1 => A(26), A2 => n278, B1 => B(26), B2 => n275, 
                           ZN => n35);
   U95 : AOI222_X1 port map( A1 => D(26), A2 => n287, B1 => C(26), B2 => n284, 
                           C1 => E(26), C2 => n281, ZN => n36);
   U96 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U97 : AOI22_X1 port map( A1 => A(22), A2 => n278, B1 => B(22), B2 => n275, 
                           ZN => n43);
   U98 : AOI222_X1 port map( A1 => D(22), A2 => n287, B1 => C(22), B2 => n284, 
                           C1 => E(22), C2 => n281, ZN => n44);
   U99 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U100 : AOI22_X1 port map( A1 => A(27), A2 => n278, B1 => B(27), B2 => n275, 
                           ZN => n33);
   U101 : AOI222_X1 port map( A1 => D(27), A2 => n287, B1 => C(27), B2 => n284,
                           C1 => E(27), C2 => n281, ZN => n34);
   U102 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U103 : AOI22_X1 port map( A1 => A(23), A2 => n278, B1 => B(23), B2 => n275, 
                           ZN => n41);
   U104 : AOI222_X1 port map( A1 => D(23), A2 => n287, B1 => C(23), B2 => n284,
                           C1 => E(23), C2 => n281, ZN => n42);
   U105 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U106 : AOI22_X1 port map( A1 => A(0), A2 => n277, B1 => B(0), B2 => n274, ZN
                           => n71);
   U107 : AOI222_X1 port map( A1 => D(0), A2 => n286, B1 => C(0), B2 => n283, 
                           C1 => E(0), C2 => n280, ZN => n72);
   U108 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U109 : AOI22_X1 port map( A1 => A(28), A2 => n278, B1 => B(28), B2 => n275, 
                           ZN => n31);
   U110 : AOI222_X1 port map( A1 => D(28), A2 => n287, B1 => C(28), B2 => n284,
                           C1 => E(28), C2 => n281, ZN => n32);
   U111 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U112 : AOI22_X1 port map( A1 => A(24), A2 => n278, B1 => B(24), B2 => n275, 
                           ZN => n39);
   U113 : AOI222_X1 port map( A1 => D(24), A2 => n287, B1 => C(24), B2 => n284,
                           C1 => E(24), C2 => n281, ZN => n40);
   U114 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U115 : AOI22_X1 port map( A1 => A(29), A2 => n278, B1 => B(29), B2 => n275, 
                           ZN => n29);
   U116 : AOI222_X1 port map( A1 => D(29), A2 => n287, B1 => C(29), B2 => n284,
                           C1 => E(29), C2 => n281, ZN => n30);
   U117 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U118 : AOI22_X1 port map( A1 => A(30), A2 => n278, B1 => B(30), B2 => n275, 
                           ZN => n25);
   U119 : AOI222_X1 port map( A1 => D(30), A2 => n287, B1 => C(30), B2 => n284,
                           C1 => E(30), C2 => n281, ZN => n26);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_6 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_6;

architecture SYN_behav of mux_N32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n277);
   U2 : BUF_X1 port map( A => n10, Z => n278);
   U3 : BUF_X1 port map( A => n10, Z => n279);
   U4 : BUF_X1 port map( A => n6, Z => n289);
   U5 : BUF_X1 port map( A => n6, Z => n290);
   U6 : BUF_X1 port map( A => n9, Z => n280);
   U7 : BUF_X1 port map( A => n9, Z => n281);
   U8 : BUF_X1 port map( A => n7, Z => n286);
   U9 : BUF_X1 port map( A => n7, Z => n287);
   U10 : BUF_X1 port map( A => n8, Z => n283);
   U11 : BUF_X1 port map( A => n8, Z => n284);
   U12 : BUF_X1 port map( A => n9, Z => n282);
   U13 : BUF_X1 port map( A => n7, Z => n288);
   U14 : BUF_X1 port map( A => n8, Z => n285);
   U15 : BUF_X1 port map( A => n6, Z => n291);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U23 : AOI22_X1 port map( A1 => A(24), A2 => n281, B1 => B(24), B2 => n278, 
                           ZN => n39);
   U24 : AOI222_X1 port map( A1 => D(24), A2 => n290, B1 => E(24), B2 => n287, 
                           C1 => C(24), C2 => n284, ZN => n40);
   U25 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U26 : AOI22_X1 port map( A1 => A(25), A2 => n281, B1 => B(25), B2 => n278, 
                           ZN => n37);
   U27 : AOI222_X1 port map( A1 => D(25), A2 => n290, B1 => E(25), B2 => n287, 
                           C1 => C(25), C2 => n284, ZN => n38);
   U28 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U29 : AOI22_X1 port map( A1 => A(28), A2 => n281, B1 => B(28), B2 => n278, 
                           ZN => n31);
   U30 : AOI222_X1 port map( A1 => D(28), A2 => n290, B1 => E(28), B2 => n287, 
                           C1 => C(28), C2 => n284, ZN => n32);
   U31 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U32 : AOI22_X1 port map( A1 => A(29), A2 => n281, B1 => B(29), B2 => n278, 
                           ZN => n29);
   U33 : AOI222_X1 port map( A1 => D(29), A2 => n290, B1 => E(29), B2 => n287, 
                           C1 => C(29), C2 => n284, ZN => n30);
   U34 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U35 : AOI22_X1 port map( A1 => A(30), A2 => n281, B1 => B(30), B2 => n278, 
                           ZN => n25);
   U36 : AOI222_X1 port map( A1 => D(30), A2 => n290, B1 => E(30), B2 => n287, 
                           C1 => C(30), C2 => n284, ZN => n26);
   U37 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U38 : AOI22_X1 port map( A1 => A(31), A2 => n282, B1 => B(31), B2 => n279, 
                           ZN => n23);
   U39 : AOI222_X1 port map( A1 => D(31), A2 => n291, B1 => E(31), B2 => n288, 
                           C1 => C(31), C2 => n285, ZN => n24);
   U40 : INV_X1 port map( A => Sel(2), ZN => n74);
   U41 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U42 : AOI22_X1 port map( A1 => A(18), A2 => n280, B1 => B(18), B2 => n277, 
                           ZN => n53);
   U43 : AOI222_X1 port map( A1 => D(18), A2 => n289, B1 => E(18), B2 => n286, 
                           C1 => C(18), C2 => n283, ZN => n54);
   U44 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n282, B1 => B(4), B2 => n279, ZN 
                           => n19);
   U46 : AOI222_X1 port map( A1 => D(4), A2 => n291, B1 => E(4), B2 => n288, C1
                           => C(4), C2 => n285, ZN => n20);
   U47 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U48 : AOI22_X1 port map( A1 => A(14), A2 => n280, B1 => B(14), B2 => n277, 
                           ZN => n61);
   U49 : AOI222_X1 port map( A1 => D(14), A2 => n289, B1 => E(14), B2 => n286, 
                           C1 => C(14), C2 => n283, ZN => n62);
   U50 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U51 : AOI22_X1 port map( A1 => A(21), A2 => n281, B1 => B(21), B2 => n278, 
                           ZN => n45);
   U52 : AOI222_X1 port map( A1 => D(21), A2 => n290, B1 => E(21), B2 => n287, 
                           C1 => C(21), C2 => n284, ZN => n46);
   U53 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n281, B1 => B(22), B2 => n278, 
                           ZN => n43);
   U55 : AOI222_X1 port map( A1 => D(22), A2 => n290, B1 => E(22), B2 => n287, 
                           C1 => C(22), C2 => n284, ZN => n44);
   U56 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U57 : AOI22_X1 port map( A1 => A(8), A2 => n282, B1 => B(8), B2 => n279, ZN 
                           => n11);
   U58 : AOI222_X1 port map( A1 => D(8), A2 => n291, B1 => E(8), B2 => n288, C1
                           => C(8), C2 => n285, ZN => n12);
   U59 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U60 : AOI22_X1 port map( A1 => A(5), A2 => n282, B1 => B(5), B2 => n279, ZN 
                           => n17);
   U61 : AOI222_X1 port map( A1 => D(5), A2 => n291, B1 => E(5), B2 => n288, C1
                           => C(5), C2 => n285, ZN => n18);
   U62 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U63 : AOI22_X1 port map( A1 => A(20), A2 => n281, B1 => B(20), B2 => n278, 
                           ZN => n47);
   U64 : AOI222_X1 port map( A1 => D(20), A2 => n290, B1 => E(20), B2 => n287, 
                           C1 => C(20), C2 => n284, ZN => n48);
   U65 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U66 : AOI22_X1 port map( A1 => A(26), A2 => n281, B1 => B(26), B2 => n278, 
                           ZN => n35);
   U67 : AOI222_X1 port map( A1 => D(26), A2 => n290, B1 => E(26), B2 => n287, 
                           C1 => C(26), C2 => n284, ZN => n36);
   U68 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U69 : AOI22_X1 port map( A1 => A(27), A2 => n281, B1 => B(27), B2 => n278, 
                           ZN => n33);
   U70 : AOI222_X1 port map( A1 => D(27), A2 => n290, B1 => E(27), B2 => n287, 
                           C1 => C(27), C2 => n284, ZN => n34);
   U71 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U72 : AOI22_X1 port map( A1 => A(23), A2 => n281, B1 => B(23), B2 => n278, 
                           ZN => n41);
   U73 : AOI222_X1 port map( A1 => D(23), A2 => n290, B1 => E(23), B2 => n287, 
                           C1 => C(23), C2 => n284, ZN => n42);
   U74 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U75 : AOI22_X1 port map( A1 => A(6), A2 => n282, B1 => B(6), B2 => n279, ZN 
                           => n15);
   U76 : AOI222_X1 port map( A1 => D(6), A2 => n291, B1 => E(6), B2 => n288, C1
                           => C(6), C2 => n285, ZN => n16);
   U77 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U78 : AOI22_X1 port map( A1 => A(10), A2 => n280, B1 => B(10), B2 => n277, 
                           ZN => n69);
   U79 : AOI222_X1 port map( A1 => D(10), A2 => n289, B1 => E(10), B2 => n286, 
                           C1 => C(10), C2 => n283, ZN => n70);
   U80 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U81 : AOI22_X1 port map( A1 => A(17), A2 => n280, B1 => B(17), B2 => n277, 
                           ZN => n55);
   U82 : AOI222_X1 port map( A1 => D(17), A2 => n289, B1 => E(17), B2 => n286, 
                           C1 => C(17), C2 => n283, ZN => n56);
   U83 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U84 : AOI22_X1 port map( A1 => A(13), A2 => n280, B1 => B(13), B2 => n277, 
                           ZN => n63);
   U85 : AOI222_X1 port map( A1 => D(13), A2 => n289, B1 => E(13), B2 => n286, 
                           C1 => C(13), C2 => n283, ZN => n64);
   U86 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U87 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U88 : AOI22_X1 port map( A1 => A(7), A2 => n282, B1 => B(7), B2 => n279, ZN 
                           => n13);
   U89 : AOI222_X1 port map( A1 => D(7), A2 => n291, B1 => E(7), B2 => n288, C1
                           => C(7), C2 => n285, ZN => n14);
   U90 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U91 : AOI22_X1 port map( A1 => A(9), A2 => n282, B1 => B(9), B2 => n279, ZN 
                           => n4);
   U92 : AOI222_X1 port map( A1 => D(9), A2 => n291, B1 => E(9), B2 => n288, C1
                           => C(9), C2 => n285, ZN => n5);
   U93 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U94 : AOI22_X1 port map( A1 => A(12), A2 => n280, B1 => B(12), B2 => n277, 
                           ZN => n65);
   U95 : AOI222_X1 port map( A1 => D(12), A2 => n289, B1 => E(12), B2 => n286, 
                           C1 => C(12), C2 => n283, ZN => n66);
   U96 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U97 : AOI22_X1 port map( A1 => A(16), A2 => n280, B1 => B(16), B2 => n277, 
                           ZN => n57);
   U98 : AOI222_X1 port map( A1 => D(16), A2 => n289, B1 => E(16), B2 => n286, 
                           C1 => C(16), C2 => n283, ZN => n58);
   U99 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U100 : AOI22_X1 port map( A1 => A(15), A2 => n280, B1 => B(15), B2 => n277, 
                           ZN => n59);
   U101 : AOI222_X1 port map( A1 => D(15), A2 => n289, B1 => E(15), B2 => n286,
                           C1 => C(15), C2 => n283, ZN => n60);
   U102 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U103 : AOI22_X1 port map( A1 => A(11), A2 => n280, B1 => B(11), B2 => n277, 
                           ZN => n67);
   U104 : AOI222_X1 port map( A1 => D(11), A2 => n289, B1 => E(11), B2 => n286,
                           C1 => C(11), C2 => n283, ZN => n68);
   U105 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U106 : AOI22_X1 port map( A1 => A(3), A2 => n282, B1 => B(3), B2 => n279, ZN
                           => n21);
   U107 : AOI222_X1 port map( A1 => D(3), A2 => n291, B1 => E(3), B2 => n288, 
                           C1 => C(3), C2 => n285, ZN => n22);
   U108 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U109 : AOI22_X1 port map( A1 => A(0), A2 => n280, B1 => B(0), B2 => n277, ZN
                           => n71);
   U110 : AOI222_X1 port map( A1 => D(0), A2 => n289, B1 => E(0), B2 => n286, 
                           C1 => C(0), C2 => n283, ZN => n72);
   U111 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U112 : AOI22_X1 port map( A1 => A(1), A2 => n280, B1 => B(1), B2 => n277, ZN
                           => n49);
   U113 : AOI222_X1 port map( A1 => D(1), A2 => n289, B1 => E(1), B2 => n286, 
                           C1 => C(1), C2 => n283, ZN => n50);
   U114 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U115 : AOI22_X1 port map( A1 => A(2), A2 => n281, B1 => B(2), B2 => n278, ZN
                           => n27);
   U116 : AOI222_X1 port map( A1 => D(2), A2 => n290, B1 => E(2), B2 => n287, 
                           C1 => C(2), C2 => n284, ZN => n28);
   U117 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U118 : AOI22_X1 port map( A1 => A(19), A2 => n280, B1 => B(19), B2 => n277, 
                           ZN => n51);
   U119 : AOI222_X1 port map( A1 => D(19), A2 => n289, B1 => E(19), B2 => n286,
                           C1 => C(19), C2 => n283, ZN => n52);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_7 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_7;

architecture SYN_behav of mux_N32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n325);
   U2 : BUF_X1 port map( A => n10, Z => n326);
   U3 : BUF_X1 port map( A => n10, Z => n327);
   U4 : BUF_X1 port map( A => n6, Z => n337);
   U5 : BUF_X1 port map( A => n6, Z => n338);
   U6 : BUF_X1 port map( A => n9, Z => n328);
   U7 : BUF_X1 port map( A => n9, Z => n329);
   U8 : BUF_X1 port map( A => n7, Z => n334);
   U9 : BUF_X1 port map( A => n7, Z => n335);
   U10 : BUF_X1 port map( A => n8, Z => n331);
   U11 : BUF_X1 port map( A => n8, Z => n332);
   U12 : BUF_X1 port map( A => n9, Z => n330);
   U13 : BUF_X1 port map( A => n7, Z => n336);
   U14 : BUF_X1 port map( A => n8, Z => n333);
   U15 : BUF_X1 port map( A => n6, Z => n339);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U24 : AOI22_X1 port map( A1 => A(16), A2 => n328, B1 => B(16), B2 => n325, 
                           ZN => n57);
   U25 : AOI222_X1 port map( A1 => D(16), A2 => n337, B1 => E(16), B2 => n334, 
                           C1 => C(16), C2 => n331, ZN => n58);
   U26 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U27 : AOI22_X1 port map( A1 => A(2), A2 => n329, B1 => B(2), B2 => n326, ZN 
                           => n27);
   U28 : AOI222_X1 port map( A1 => D(2), A2 => n338, B1 => E(2), B2 => n335, C1
                           => C(2), C2 => n332, ZN => n28);
   U29 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U30 : AOI22_X1 port map( A1 => A(12), A2 => n328, B1 => B(12), B2 => n325, 
                           ZN => n65);
   U31 : AOI222_X1 port map( A1 => D(12), A2 => n337, B1 => E(12), B2 => n334, 
                           C1 => C(12), C2 => n331, ZN => n66);
   U32 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U33 : AOI22_X1 port map( A1 => A(6), A2 => n330, B1 => B(6), B2 => n327, ZN 
                           => n15);
   U34 : AOI222_X1 port map( A1 => D(6), A2 => n339, B1 => E(6), B2 => n336, C1
                           => C(6), C2 => n333, ZN => n16);
   U35 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U36 : AOI22_X1 port map( A1 => A(3), A2 => n330, B1 => B(3), B2 => n327, ZN 
                           => n21);
   U37 : AOI222_X1 port map( A1 => D(3), A2 => n339, B1 => E(3), B2 => n336, C1
                           => C(3), C2 => n333, ZN => n22);
   U38 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U39 : AOI22_X1 port map( A1 => A(10), A2 => n328, B1 => B(10), B2 => n325, 
                           ZN => n69);
   U40 : AOI222_X1 port map( A1 => D(10), A2 => n337, B1 => E(10), B2 => n334, 
                           C1 => C(10), C2 => n331, ZN => n70);
   U41 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n330, B1 => B(4), B2 => n327, ZN 
                           => n19);
   U43 : AOI222_X1 port map( A1 => D(4), A2 => n339, B1 => E(4), B2 => n336, C1
                           => C(4), C2 => n333, ZN => n20);
   U44 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U45 : AOI22_X1 port map( A1 => A(8), A2 => n330, B1 => B(8), B2 => n327, ZN 
                           => n11);
   U46 : AOI222_X1 port map( A1 => D(8), A2 => n339, B1 => E(8), B2 => n336, C1
                           => C(8), C2 => n333, ZN => n12);
   U47 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U48 : AOI22_X1 port map( A1 => A(15), A2 => n328, B1 => B(15), B2 => n325, 
                           ZN => n59);
   U49 : AOI222_X1 port map( A1 => D(15), A2 => n337, B1 => E(15), B2 => n334, 
                           C1 => C(15), C2 => n331, ZN => n60);
   U50 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U51 : AOI22_X1 port map( A1 => A(11), A2 => n328, B1 => B(11), B2 => n325, 
                           ZN => n67);
   U52 : AOI222_X1 port map( A1 => D(11), A2 => n337, B1 => E(11), B2 => n334, 
                           C1 => C(11), C2 => n331, ZN => n68);
   U53 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U54 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n329, B1 => B(25), B2 => n326, 
                           ZN => n37);
   U56 : AOI222_X1 port map( A1 => D(25), A2 => n338, B1 => E(25), B2 => n335, 
                           C1 => C(25), C2 => n332, ZN => n38);
   U57 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U58 : AOI22_X1 port map( A1 => A(26), A2 => n329, B1 => B(26), B2 => n326, 
                           ZN => n35);
   U59 : AOI222_X1 port map( A1 => D(26), A2 => n338, B1 => E(26), B2 => n335, 
                           C1 => C(26), C2 => n332, ZN => n36);
   U60 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U61 : AOI22_X1 port map( A1 => A(22), A2 => n329, B1 => B(22), B2 => n326, 
                           ZN => n43);
   U62 : AOI222_X1 port map( A1 => D(22), A2 => n338, B1 => E(22), B2 => n335, 
                           C1 => C(22), C2 => n332, ZN => n44);
   U63 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n329, B1 => B(27), B2 => n326, 
                           ZN => n33);
   U65 : AOI222_X1 port map( A1 => D(27), A2 => n338, B1 => E(27), B2 => n335, 
                           C1 => C(27), C2 => n332, ZN => n34);
   U66 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U67 : AOI22_X1 port map( A1 => A(19), A2 => n328, B1 => B(19), B2 => n325, 
                           ZN => n51);
   U68 : AOI222_X1 port map( A1 => D(19), A2 => n337, B1 => E(19), B2 => n334, 
                           C1 => C(19), C2 => n331, ZN => n52);
   U69 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U70 : AOI22_X1 port map( A1 => A(28), A2 => n329, B1 => B(28), B2 => n326, 
                           ZN => n31);
   U71 : AOI222_X1 port map( A1 => D(28), A2 => n338, B1 => E(28), B2 => n335, 
                           C1 => C(28), C2 => n332, ZN => n32);
   U72 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U73 : AOI22_X1 port map( A1 => A(29), A2 => n329, B1 => B(29), B2 => n326, 
                           ZN => n29);
   U74 : AOI222_X1 port map( A1 => D(29), A2 => n338, B1 => E(29), B2 => n335, 
                           C1 => C(29), C2 => n332, ZN => n30);
   U75 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U76 : AOI22_X1 port map( A1 => A(5), A2 => n330, B1 => B(5), B2 => n327, ZN 
                           => n17);
   U77 : AOI222_X1 port map( A1 => D(5), A2 => n339, B1 => E(5), B2 => n336, C1
                           => C(5), C2 => n333, ZN => n18);
   U78 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U79 : AOI22_X1 port map( A1 => A(9), A2 => n330, B1 => B(9), B2 => n327, ZN 
                           => n4);
   U80 : AOI222_X1 port map( A1 => D(9), A2 => n339, B1 => E(9), B2 => n336, C1
                           => C(9), C2 => n333, ZN => n5);
   U81 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U82 : AOI22_X1 port map( A1 => A(7), A2 => n330, B1 => B(7), B2 => n327, ZN 
                           => n13);
   U83 : AOI222_X1 port map( A1 => D(7), A2 => n339, B1 => E(7), B2 => n336, C1
                           => C(7), C2 => n333, ZN => n14);
   U84 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U85 : AOI22_X1 port map( A1 => A(13), A2 => n328, B1 => B(13), B2 => n325, 
                           ZN => n63);
   U86 : AOI222_X1 port map( A1 => D(13), A2 => n337, B1 => E(13), B2 => n334, 
                           C1 => C(13), C2 => n331, ZN => n64);
   U87 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U88 : AOI22_X1 port map( A1 => A(17), A2 => n328, B1 => B(17), B2 => n325, 
                           ZN => n55);
   U89 : AOI222_X1 port map( A1 => D(17), A2 => n337, B1 => E(17), B2 => n334, 
                           C1 => C(17), C2 => n331, ZN => n56);
   U90 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U91 : AOI22_X1 port map( A1 => A(14), A2 => n328, B1 => B(14), B2 => n325, 
                           ZN => n61);
   U92 : AOI222_X1 port map( A1 => D(14), A2 => n337, B1 => E(14), B2 => n334, 
                           C1 => C(14), C2 => n331, ZN => n62);
   U93 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U94 : AOI22_X1 port map( A1 => A(23), A2 => n329, B1 => B(23), B2 => n326, 
                           ZN => n41);
   U95 : AOI222_X1 port map( A1 => D(23), A2 => n338, B1 => E(23), B2 => n335, 
                           C1 => C(23), C2 => n332, ZN => n42);
   U96 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U97 : AOI22_X1 port map( A1 => A(24), A2 => n329, B1 => B(24), B2 => n326, 
                           ZN => n39);
   U98 : AOI222_X1 port map( A1 => D(24), A2 => n338, B1 => E(24), B2 => n335, 
                           C1 => C(24), C2 => n332, ZN => n40);
   U99 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U100 : AOI22_X1 port map( A1 => A(20), A2 => n329, B1 => B(20), B2 => n326, 
                           ZN => n47);
   U101 : AOI222_X1 port map( A1 => D(20), A2 => n338, B1 => E(20), B2 => n335,
                           C1 => C(20), C2 => n332, ZN => n48);
   U102 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U103 : AOI22_X1 port map( A1 => A(21), A2 => n329, B1 => B(21), B2 => n326, 
                           ZN => n45);
   U104 : AOI222_X1 port map( A1 => D(21), A2 => n338, B1 => E(21), B2 => n335,
                           C1 => C(21), C2 => n332, ZN => n46);
   U105 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U106 : AOI22_X1 port map( A1 => A(18), A2 => n328, B1 => B(18), B2 => n325, 
                           ZN => n53);
   U107 : AOI222_X1 port map( A1 => D(18), A2 => n337, B1 => E(18), B2 => n334,
                           C1 => C(18), C2 => n331, ZN => n54);
   U108 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U109 : AOI22_X1 port map( A1 => A(30), A2 => n329, B1 => B(30), B2 => n326, 
                           ZN => n25);
   U110 : AOI222_X1 port map( A1 => D(30), A2 => n338, B1 => E(30), B2 => n335,
                           C1 => C(30), C2 => n332, ZN => n26);
   U111 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U112 : AOI22_X1 port map( A1 => A(31), A2 => n330, B1 => B(31), B2 => n327, 
                           ZN => n23);
   U113 : AOI222_X1 port map( A1 => D(31), A2 => n339, B1 => E(31), B2 => n336,
                           C1 => C(31), C2 => n333, ZN => n24);
   U114 : INV_X1 port map( A => Sel(1), ZN => n75);
   U115 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U116 : AOI22_X1 port map( A1 => A(0), A2 => n328, B1 => B(0), B2 => n325, ZN
                           => n71);
   U117 : AOI222_X1 port map( A1 => D(0), A2 => n337, B1 => E(0), B2 => n334, 
                           C1 => C(0), C2 => n331, ZN => n72);
   U118 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U119 : AOI22_X1 port map( A1 => A(1), A2 => n328, B1 => B(1), B2 => n325, ZN
                           => n49);
   U120 : AOI222_X1 port map( A1 => D(1), A2 => n337, B1 => E(1), B2 => n334, 
                           C1 => C(1), C2 => n331, ZN => n50);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_N32_0 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_0;

architecture SYN_behav of mux_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286 : std_logic;

begin
   
   U105 : OAI33_X1 port map( A1 => n73, A2 => n75, A3 => n76, B1 => Sel(0), B2 
                           => Sel(2), B3 => Sel(1), ZN => n9);
   U1 : BUF_X1 port map( A => n10, Z => n272);
   U2 : BUF_X1 port map( A => n10, Z => n273);
   U3 : BUF_X1 port map( A => n10, Z => n274);
   U4 : BUF_X1 port map( A => n6, Z => n284);
   U5 : BUF_X1 port map( A => n6, Z => n285);
   U6 : BUF_X1 port map( A => n9, Z => n275);
   U7 : BUF_X1 port map( A => n9, Z => n276);
   U8 : BUF_X1 port map( A => n7, Z => n281);
   U9 : BUF_X1 port map( A => n7, Z => n282);
   U10 : BUF_X1 port map( A => n9, Z => n277);
   U11 : BUF_X1 port map( A => n8, Z => n278);
   U12 : BUF_X1 port map( A => n8, Z => n279);
   U13 : BUF_X1 port map( A => n7, Z => n283);
   U14 : BUF_X1 port map( A => n8, Z => n280);
   U15 : BUF_X1 port map( A => n6, Z => n286);
   U16 : AND2_X1 port map( A1 => n74, A2 => n73, ZN => n10);
   U17 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n73, ZN => n8);
   U18 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U19 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n74);
   U20 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U21 : AOI22_X1 port map( A1 => A(14), A2 => n275, B1 => B(14), B2 => n272, 
                           ZN => n61);
   U22 : AOI222_X1 port map( A1 => D(14), A2 => n284, B1 => C(14), B2 => n281, 
                           C1 => E(14), C2 => n278, ZN => n62);
   U23 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U24 : AOI22_X1 port map( A1 => A(1), A2 => n275, B1 => B(1), B2 => n272, ZN 
                           => n49);
   U25 : AOI222_X1 port map( A1 => D(1), A2 => n284, B1 => C(1), B2 => n281, C1
                           => E(1), C2 => n278, ZN => n50);
   U26 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U27 : AOI22_X1 port map( A1 => A(10), A2 => n275, B1 => B(10), B2 => n272, 
                           ZN => n69);
   U28 : AOI222_X1 port map( A1 => D(10), A2 => n284, B1 => C(10), B2 => n281, 
                           C1 => E(10), C2 => n278, ZN => n70);
   U29 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U30 : AOI22_X1 port map( A1 => A(4), A2 => n277, B1 => B(4), B2 => n274, ZN 
                           => n19);
   U31 : AOI222_X1 port map( A1 => D(4), A2 => n286, B1 => C(4), B2 => n283, C1
                           => E(4), C2 => n280, ZN => n20);
   U32 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U33 : AOI22_X1 port map( A1 => A(0), A2 => n275, B1 => B(0), B2 => n272, ZN 
                           => n71);
   U34 : AOI222_X1 port map( A1 => D(0), A2 => n284, B1 => C(0), B2 => n281, C1
                           => E(0), C2 => n278, ZN => n72);
   U35 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n277, B1 => B(8), B2 => n274, ZN 
                           => n11);
   U37 : AOI222_X1 port map( A1 => D(8), A2 => n286, B1 => C(8), B2 => n283, C1
                           => E(8), C2 => n280, ZN => n12);
   U38 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U39 : AOI22_X1 port map( A1 => A(2), A2 => n276, B1 => B(2), B2 => n273, ZN 
                           => n27);
   U40 : AOI222_X1 port map( A1 => D(2), A2 => n285, B1 => C(2), B2 => n282, C1
                           => E(2), C2 => n279, ZN => n28);
   U41 : INV_X1 port map( A => Sel(2), ZN => n73);
   U42 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U43 : AOI22_X1 port map( A1 => A(13), A2 => n275, B1 => B(13), B2 => n272, 
                           ZN => n63);
   U44 : AOI222_X1 port map( A1 => D(13), A2 => n284, B1 => C(13), B2 => n281, 
                           C1 => E(13), C2 => n278, ZN => n64);
   U45 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U46 : AOI22_X1 port map( A1 => A(9), A2 => n277, B1 => B(9), B2 => n274, ZN 
                           => n4);
   U47 : AOI222_X1 port map( A1 => D(9), A2 => n286, B1 => C(9), B2 => n283, C1
                           => E(9), C2 => n280, ZN => n5);
   U48 : AND2_X1 port map( A1 => Sel(2), A2 => n74, ZN => n7);
   U49 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U50 : AOI22_X1 port map( A1 => A(3), A2 => n277, B1 => B(3), B2 => n274, ZN 
                           => n21);
   U51 : AOI222_X1 port map( A1 => D(3), A2 => n286, B1 => C(3), B2 => n283, C1
                           => E(3), C2 => n280, ZN => n22);
   U52 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U53 : AOI22_X1 port map( A1 => A(7), A2 => n277, B1 => B(7), B2 => n274, ZN 
                           => n13);
   U54 : AOI222_X1 port map( A1 => D(7), A2 => n286, B1 => C(7), B2 => n283, C1
                           => E(7), C2 => n280, ZN => n14);
   U55 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U56 : AOI22_X1 port map( A1 => A(15), A2 => n275, B1 => B(15), B2 => n272, 
                           ZN => n59);
   U57 : AOI222_X1 port map( A1 => D(15), A2 => n284, B1 => C(15), B2 => n281, 
                           C1 => E(15), C2 => n278, ZN => n60);
   U58 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U59 : AOI22_X1 port map( A1 => A(11), A2 => n275, B1 => B(11), B2 => n272, 
                           ZN => n67);
   U60 : AOI222_X1 port map( A1 => D(11), A2 => n284, B1 => C(11), B2 => n281, 
                           C1 => E(11), C2 => n278, ZN => n68);
   U61 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U62 : AOI22_X1 port map( A1 => A(12), A2 => n275, B1 => B(12), B2 => n272, 
                           ZN => n65);
   U63 : AOI222_X1 port map( A1 => D(12), A2 => n284, B1 => C(12), B2 => n281, 
                           C1 => E(12), C2 => n278, ZN => n66);
   U64 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U65 : AOI22_X1 port map( A1 => A(6), A2 => n277, B1 => B(6), B2 => n274, ZN 
                           => n15);
   U66 : AOI222_X1 port map( A1 => D(6), A2 => n286, B1 => C(6), B2 => n283, C1
                           => E(6), C2 => n280, ZN => n16);
   U67 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U68 : AOI22_X1 port map( A1 => A(24), A2 => n276, B1 => B(24), B2 => n273, 
                           ZN => n39);
   U69 : AOI222_X1 port map( A1 => D(24), A2 => n285, B1 => C(24), B2 => n282, 
                           C1 => E(24), C2 => n279, ZN => n40);
   U70 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U71 : AOI22_X1 port map( A1 => A(20), A2 => n276, B1 => B(20), B2 => n273, 
                           ZN => n47);
   U72 : AOI222_X1 port map( A1 => D(20), A2 => n285, B1 => C(20), B2 => n282, 
                           C1 => E(20), C2 => n279, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U74 : AOI22_X1 port map( A1 => A(25), A2 => n276, B1 => B(25), B2 => n273, 
                           ZN => n37);
   U75 : AOI222_X1 port map( A1 => D(25), A2 => n285, B1 => C(25), B2 => n282, 
                           C1 => E(25), C2 => n279, ZN => n38);
   U76 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U77 : AOI22_X1 port map( A1 => A(21), A2 => n276, B1 => B(21), B2 => n273, 
                           ZN => n45);
   U78 : AOI222_X1 port map( A1 => D(21), A2 => n285, B1 => C(21), B2 => n282, 
                           C1 => E(21), C2 => n279, ZN => n46);
   U79 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U80 : AOI22_X1 port map( A1 => A(17), A2 => n275, B1 => B(17), B2 => n272, 
                           ZN => n55);
   U81 : AOI222_X1 port map( A1 => D(17), A2 => n284, B1 => C(17), B2 => n281, 
                           C1 => E(17), C2 => n278, ZN => n56);
   U82 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U83 : AOI22_X1 port map( A1 => A(26), A2 => n276, B1 => B(26), B2 => n273, 
                           ZN => n35);
   U84 : AOI222_X1 port map( A1 => D(26), A2 => n285, B1 => C(26), B2 => n282, 
                           C1 => E(26), C2 => n279, ZN => n36);
   U85 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U86 : AOI22_X1 port map( A1 => A(22), A2 => n276, B1 => B(22), B2 => n273, 
                           ZN => n43);
   U87 : AOI222_X1 port map( A1 => D(22), A2 => n285, B1 => C(22), B2 => n282, 
                           C1 => E(22), C2 => n279, ZN => n44);
   U88 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U89 : AOI22_X1 port map( A1 => A(18), A2 => n275, B1 => B(18), B2 => n272, 
                           ZN => n53);
   U90 : AOI222_X1 port map( A1 => D(18), A2 => n284, B1 => C(18), B2 => n281, 
                           C1 => E(18), C2 => n278, ZN => n54);
   U91 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U92 : AOI22_X1 port map( A1 => A(27), A2 => n276, B1 => B(27), B2 => n273, 
                           ZN => n33);
   U93 : AOI222_X1 port map( A1 => D(27), A2 => n285, B1 => C(27), B2 => n282, 
                           C1 => E(27), C2 => n279, ZN => n34);
   U94 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U95 : AOI22_X1 port map( A1 => A(23), A2 => n276, B1 => B(23), B2 => n273, 
                           ZN => n41);
   U96 : AOI222_X1 port map( A1 => D(23), A2 => n285, B1 => C(23), B2 => n282, 
                           C1 => E(23), C2 => n279, ZN => n42);
   U97 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U98 : AOI22_X1 port map( A1 => A(19), A2 => n275, B1 => B(19), B2 => n272, 
                           ZN => n51);
   U99 : AOI222_X1 port map( A1 => D(19), A2 => n284, B1 => C(19), B2 => n281, 
                           C1 => E(19), C2 => n278, ZN => n52);
   U100 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U101 : AOI22_X1 port map( A1 => A(28), A2 => n276, B1 => B(28), B2 => n273, 
                           ZN => n31);
   U102 : AOI222_X1 port map( A1 => D(28), A2 => n285, B1 => C(28), B2 => n282,
                           C1 => E(28), C2 => n279, ZN => n32);
   U103 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U104 : AOI22_X1 port map( A1 => A(29), A2 => n276, B1 => B(29), B2 => n273, 
                           ZN => n29);
   U106 : AOI222_X1 port map( A1 => D(29), A2 => n285, B1 => C(29), B2 => n282,
                           C1 => E(29), C2 => n279, ZN => n30);
   U107 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U108 : AOI22_X1 port map( A1 => A(30), A2 => n276, B1 => B(30), B2 => n273, 
                           ZN => n25);
   U109 : AOI222_X1 port map( A1 => D(30), A2 => n285, B1 => C(30), B2 => n282,
                           C1 => E(30), C2 => n279, ZN => n26);
   U110 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U111 : AOI22_X1 port map( A1 => A(31), A2 => n277, B1 => B(31), B2 => n274, 
                           ZN => n23);
   U112 : AOI222_X1 port map( A1 => D(31), A2 => n286, B1 => C(31), B2 => n283,
                           C1 => E(31), C2 => n280, ZN => n24);
   U113 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U114 : AOI22_X1 port map( A1 => A(16), A2 => n275, B1 => B(16), B2 => n272, 
                           ZN => n57);
   U115 : AOI222_X1 port map( A1 => D(16), A2 => n284, B1 => C(16), B2 => n281,
                           C1 => E(16), C2 => n278, ZN => n58);
   U116 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U117 : AOI22_X1 port map( A1 => A(5), A2 => n277, B1 => B(5), B2 => n274, ZN
                           => n17);
   U118 : AOI222_X1 port map( A1 => D(5), A2 => n286, B1 => C(5), B2 => n283, 
                           C1 => E(5), C2 => n280, ZN => n18);
   U119 : INV_X1 port map( A => Sel(1), ZN => n75);
   U120 : INV_X1 port map( A => Sel(0), ZN => n76);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S14 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S14;

architecture SYN_struct of shift_mul_N16_S14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_31_port, E_30_port, E_29_port, E_28_port, E_27_port,
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, n9, n10, n12, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n62, n63, 
      D_21_port, n65, D_23_port, n67, D_25_port, n69, D_27_port, n71, n72 : 
      std_logic;

begin
   B <= ( A(15), A(15), A(15), A(14), A(13), D_27_port, A(11), D_25_port, A(9),
      D_23_port, A(7), D_21_port, A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   C <= ( E_31_port, E_31_port, E_30_port, E_29_port, E_28_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   D <= ( A(15), A(15), A(14), A(13), D_27_port, A(11), D_25_port, A(9), 
      D_23_port, A(7), D_21_port, A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   E <= ( E_31_port, E_30_port, E_29_port, E_28_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n12, B => A(13), Z => E_28_port);
   U28 : XOR2_X1 port map( A => n14, B => n71, Z => E_27_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_26_port);
   U30 : XOR2_X1 port map( A => n17, B => n69, Z => E_25_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_24_port);
   U32 : XOR2_X1 port map( A => n20, B => n67, Z => E_23_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_22_port);
   U34 : XOR2_X1 port map( A => n23, B => n65, Z => E_21_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_20_port);
   U36 : XOR2_X1 port map( A => n26, B => n63, Z => E_19_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_18_port);
   U38 : XOR2_X1 port map( A => n29, B => n62, Z => E_17_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_16_port);
   U2 : INV_X1 port map( A => n9, ZN => E_31_port);
   U3 : OAI21_X1 port map( B1 => n10, B2 => n72, A => n9, ZN => E_30_port);
   U4 : NAND2_X1 port map( A1 => n14, A2 => n71, ZN => n12);
   U5 : NAND2_X1 port map( A1 => n17, A2 => n69, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n72, A2 => n10, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n26, A2 => n63, ZN => n25);
   U8 : NAND2_X1 port map( A1 => n20, A2 => n67, ZN => n19);
   U9 : NAND2_X1 port map( A1 => n23, A2 => n65, ZN => n22);
   U10 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U11 : XNOR2_X1 port map( A => A(14), B => n13, ZN => E_29_port);
   U12 : NOR2_X1 port map( A1 => A(13), A2 => n12, ZN => n13);
   U13 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U14 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U15 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U16 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U18 : INV_X1 port map( A => A(8), ZN => n67);
   U19 : INV_X1 port map( A => A(12), ZN => n71);
   U20 : INV_X1 port map( A => A(10), ZN => n69);
   U21 : INV_X1 port map( A => A(6), ZN => n65);
   U22 : INV_X1 port map( A => A(4), ZN => n63);
   U23 : INV_X1 port map( A => A(15), ZN => n72);
   U24 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n12, ZN => n10);
   U25 : NAND2_X1 port map( A1 => n29, A2 => n62, ZN => n28);
   U26 : INV_X1 port map( A => A(2), ZN => n62);
   U40 : INV_X1 port map( A => n65, ZN => D_21_port);
   U41 : INV_X1 port map( A => n67, ZN => D_23_port);
   U42 : INV_X1 port map( A => n69, ZN => D_25_port);
   U43 : INV_X1 port map( A => n71, ZN => D_27_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S12 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S12;

architecture SYN_struct of shift_mul_N16_S12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_28_port, E_27_port, E_26_port, E_25_port, E_24_port,
      E_23_port, E_22_port, E_21_port, E_20_port, E_19_port, E_18_port, 
      E_17_port, E_16_port, E_15_port, E_14_port, E_29_port, n9, n10, n11, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n66, n67, n68, 
      D_21_port, n70, n71, D_25_port, n73, n74, D_28_port : std_logic;

begin
   B <= ( D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), 
      D_25_port, A(11), A(10), A(9), D_21_port, A(7), A(6), A(5), A(4), A(3), 
      A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_29_port, E_29_port, E_29_port, E_29_port, E_28_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), D_25_port, 
      A(11), A(10), A(9), D_21_port, A(7), A(6), A(5), A(4), A(3), A(2), A(1), 
      A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_29_port, E_29_port, E_29_port, E_28_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U25 : NAND3_X1 port map( A1 => n11, A2 => n74, A3 => D_28_port, ZN => n10);
   U26 : XOR2_X1 port map( A => n11, B => n74, Z => E_27_port);
   U27 : XOR2_X1 port map( A => n13, B => A(13), Z => E_26_port);
   U28 : XOR2_X1 port map( A => n14, B => n73, Z => E_25_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_24_port);
   U30 : XOR2_X1 port map( A => n17, B => n71, Z => E_23_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_22_port);
   U32 : XOR2_X1 port map( A => n20, B => n70, Z => E_21_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_20_port);
   U34 : XOR2_X1 port map( A => n23, B => n68, Z => E_19_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_18_port);
   U36 : XOR2_X1 port map( A => n26, B => n67, Z => E_17_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_16_port);
   U38 : XOR2_X1 port map( A => n29, B => n66, Z => E_15_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_14_port);
   U2 : AOI21_X1 port map( B1 => n74, B2 => n11, A => D_28_port, ZN => 
                           E_29_port);
   U3 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => E_28_port);
   U4 : INV_X1 port map( A => E_29_port, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n17, A2 => n71, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n26, A2 => n67, ZN => n25);
   U7 : NAND2_X1 port map( A1 => n20, A2 => n70, ZN => n19);
   U8 : NAND2_X1 port map( A1 => n23, A2 => n68, ZN => n22);
   U9 : NAND2_X1 port map( A1 => n14, A2 => n73, ZN => n13);
   U10 : NOR2_X1 port map( A1 => n13, A2 => A(13), ZN => n11);
   U11 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U12 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U13 : BUF_X1 port map( A => A(15), Z => D_28_port);
   U14 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U15 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U16 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U18 : INV_X1 port map( A => A(8), ZN => n70);
   U19 : INV_X1 port map( A => A(12), ZN => n73);
   U20 : INV_X1 port map( A => A(10), ZN => n71);
   U21 : INV_X1 port map( A => A(6), ZN => n68);
   U22 : INV_X1 port map( A => A(4), ZN => n67);
   U23 : NAND2_X1 port map( A1 => n29, A2 => n66, ZN => n28);
   U24 : INV_X1 port map( A => A(2), ZN => n66);
   U40 : INV_X1 port map( A => n70, ZN => D_21_port);
   U41 : INV_X1 port map( A => n73, ZN => D_25_port);
   U42 : INV_X1 port map( A => A(14), ZN => n74);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S10 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S10;

architecture SYN_struct of shift_mul_N16_S10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port,
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_26_port, E_27_port, n9, n10, n12, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n81, n82, n83, n84
      , n85, n86, D_26_port, n88 : std_logic;

begin
   B <= ( D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, 
      D_26_port, A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, 
      A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), 
      A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n12, B => A(13), Z => E_24_port);
   U28 : XOR2_X1 port map( A => n14, B => n86, Z => E_23_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_22_port);
   U30 : XOR2_X1 port map( A => n17, B => n85, Z => E_21_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_20_port);
   U32 : XOR2_X1 port map( A => n20, B => n84, Z => E_19_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_18_port);
   U34 : XOR2_X1 port map( A => n23, B => n83, Z => E_17_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_16_port);
   U36 : XOR2_X1 port map( A => n26, B => n82, Z => E_15_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_14_port);
   U38 : XOR2_X1 port map( A => n29, B => n81, Z => E_13_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_12_port);
   U2 : INV_X1 port map( A => n9, ZN => E_27_port);
   U3 : INV_X1 port map( A => n88, ZN => D_26_port);
   U4 : OAI21_X1 port map( B1 => n10, B2 => n88, A => n9, ZN => E_26_port);
   U5 : NAND2_X1 port map( A1 => n14, A2 => n86, ZN => n12);
   U6 : NAND2_X1 port map( A1 => n17, A2 => n85, ZN => n16);
   U7 : NAND2_X1 port map( A1 => n88, A2 => n10, ZN => n9);
   U8 : NAND2_X1 port map( A1 => n26, A2 => n82, ZN => n25);
   U9 : NAND2_X1 port map( A1 => n20, A2 => n84, ZN => n19);
   U10 : NAND2_X1 port map( A1 => n23, A2 => n83, ZN => n22);
   U11 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U12 : XNOR2_X1 port map( A => A(14), B => n13, ZN => E_25_port);
   U13 : NOR2_X1 port map( A1 => A(13), A2 => n12, ZN => n13);
   U14 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U15 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U16 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U17 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U18 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U19 : INV_X1 port map( A => A(8), ZN => n84);
   U20 : INV_X1 port map( A => A(12), ZN => n86);
   U21 : INV_X1 port map( A => A(10), ZN => n85);
   U22 : INV_X1 port map( A => A(6), ZN => n83);
   U23 : INV_X1 port map( A => A(4), ZN => n82);
   U24 : INV_X1 port map( A => A(15), ZN => n88);
   U25 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n12, ZN => n10);
   U26 : NAND2_X1 port map( A1 => n29, A2 => n81, ZN => n28);
   U40 : INV_X1 port map( A => A(2), ZN => n81);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S8 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S8;

architecture SYN_struct of shift_mul_N16_S8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_23_port, E_22_port, E_21_port, E_20_port, E_19_port,
      E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, E_13_port, 
      E_12_port, E_11_port, E_10_port, E_25_port, E_24_port, n7, n8, n9, n11, 
      n13, n15, n17, n18, n19, n21, n22, n24, n25, n95, n96, D_11_port, n98, 
      D_13_port, n100, D_15_port, n102, D_20_port, n104, D_23_port, n106, 
      D_24_port, B_27_port : std_logic;

begin
   B <= ( B_27_port, B_27_port, B_27_port, B_27_port, B_27_port, D_24_port, 
      D_24_port, D_24_port, D_24_port, D_23_port, A(13), A(12), D_20_port, 
      A(10), A(9), A(8), A(7), D_15_port, A(5), D_13_port, A(3), D_11_port, 
      A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, 
      E_25_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_24_port, D_24_port, D_24_port, D_24_port, D_24_port, D_24_port, 
      D_24_port, D_24_port, D_23_port, A(13), A(12), D_20_port, A(10), A(9), 
      A(8), A(7), D_15_port, A(5), D_13_port, A(3), D_11_port, A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U29 : NAND3_X1 port map( A1 => n9, A2 => n106, A3 => B_27_port, ZN => n8);
   U31 : XOR2_X1 port map( A => n11, B => A(12), Z => E_21_port);
   U33 : XOR2_X1 port map( A => n15, B => A(9), Z => E_18_port);
   U34 : XOR2_X1 port map( A => n17, B => A(7), Z => E_16_port);
   U35 : XOR2_X1 port map( A => n21, B => A(5), Z => E_14_port);
   U36 : XOR2_X1 port map( A => n24, B => A(3), Z => E_12_port);
   U37 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_10_port);
   U2 : AOI21_X2 port map( B1 => n106, B2 => n9, A => B_27_port, ZN => 
                           E_25_port);
   U3 : XNOR2_X1 port map( A => n9, B => D_23_port, ZN => E_23_port);
   U4 : XNOR2_X1 port map( A => n13, B => D_20_port, ZN => E_20_port);
   U5 : XNOR2_X1 port map( A => n22, B => D_13_port, ZN => E_13_port);
   U6 : XNOR2_X1 port map( A => n25, B => D_11_port, ZN => E_11_port);
   U7 : XNOR2_X1 port map( A => n19, B => D_15_port, ZN => E_15_port);
   U8 : NAND2_X1 port map( A1 => n13, A2 => n104, ZN => n11);
   U9 : NAND2_X1 port map( A1 => n19, A2 => n102, ZN => n17);
   U10 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => E_24_port);
   U11 : INV_X1 port map( A => E_25_port, ZN => n7);
   U12 : NAND2_X1 port map( A1 => n22, A2 => n100, ZN => n21);
   U13 : NOR3_X1 port map( A1 => A(12), A2 => A(13), A3 => n11, ZN => n9);
   U14 : XNOR2_X1 port map( A => n95, B => A(13), ZN => E_22_port);
   U15 : NOR2_X1 port map( A1 => n11, A2 => A(12), ZN => n95);
   U16 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n15, ZN => n13);
   U17 : XNOR2_X1 port map( A => n96, B => A(10), ZN => E_19_port);
   U18 : NOR2_X1 port map( A1 => n15, A2 => A(9), ZN => n96);
   U19 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n25);
   U20 : BUF_X1 port map( A => A(15), Z => D_24_port);
   U21 : XNOR2_X1 port map( A => A(8), B => n18, ZN => E_17_port);
   U22 : NOR2_X1 port map( A1 => A(7), A2 => n17, ZN => n18);
   U23 : NOR2_X1 port map( A1 => n24, A2 => A(3), ZN => n22);
   U24 : NOR2_X1 port map( A1 => n21, A2 => A(5), ZN => n19);
   U25 : BUF_X1 port map( A => A(15), Z => B_27_port);
   U26 : NAND2_X1 port map( A1 => n25, A2 => n98, ZN => n24);
   U27 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n17, ZN => n15);
   U28 : INV_X1 port map( A => n98, ZN => D_11_port);
   U30 : INV_X1 port map( A => A(2), ZN => n98);
   U32 : INV_X1 port map( A => n100, ZN => D_13_port);
   U38 : INV_X1 port map( A => A(4), ZN => n100);
   U39 : INV_X1 port map( A => n102, ZN => D_15_port);
   U40 : INV_X1 port map( A => A(6), ZN => n102);
   U41 : INV_X1 port map( A => n104, ZN => D_20_port);
   U42 : INV_X1 port map( A => A(11), ZN => n104);
   U43 : INV_X1 port map( A => n106, ZN => D_23_port);
   U44 : INV_X1 port map( A => A(14), ZN => n106);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S6 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S6;

architecture SYN_struct of shift_mul_N16_S6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_21_port, E_20_port, E_19_port, E_18_port, E_17_port,
      E_16_port, E_15_port, E_14_port, E_13_port, E_12_port, E_11_port, 
      E_10_port, E_9_port, E_8_port, E_23_port, E_22_port, n4, n6, n7, n9, n10,
      n11, n13, n15, n16, n17, n19, n20, n87, n88, n89, n90, E_26_port, 
      E_30_port, C_31_port, C_30_port, C_24_port, C_28_port, C_22_port, 
      C_26_port, E_27_port, D_18_port, n101, n102, D_22_port, B_23_port : 
      std_logic;

begin
   B <= ( B_23_port, B_23_port, B_23_port, B_23_port, B_23_port, B_23_port, 
      B_23_port, B_23_port, B_23_port, D_22_port, D_22_port, A(14), A(13), 
      A(12), D_18_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), 
      A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   C <= ( C_31_port, C_30_port, C_24_port, C_28_port, C_22_port, C_26_port, 
      E_26_port, C_24_port, C_28_port, C_22_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   D <= ( D_22_port, D_22_port, D_22_port, D_22_port, D_22_port, D_22_port, 
      D_22_port, D_22_port, D_22_port, D_22_port, A(14), A(13), A(12), 
      D_18_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), 
      A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( C_26_port, E_30_port, E_26_port, E_27_port, E_27_port, E_26_port, 
      E_30_port, C_31_port, C_30_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U24 : XOR2_X1 port map( A => n4, B => A(2), Z => E_9_port);
   U25 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_8_port);
   U26 : NAND3_X1 port map( A1 => n7, A2 => n102, A3 => B_23_port, ZN => n6);
   U27 : XOR2_X1 port map( A => n9, B => A(13), Z => E_20_port);
   U28 : XOR2_X1 port map( A => n10, B => A(12), Z => E_19_port);
   U30 : XOR2_X1 port map( A => n13, B => A(9), Z => E_16_port);
   U31 : XOR2_X1 port map( A => n15, B => A(7), Z => E_14_port);
   U33 : XOR2_X1 port map( A => n17, B => A(5), Z => E_12_port);
   U34 : XOR2_X1 port map( A => n19, B => A(3), Z => E_10_port);
   U2 : AOI21_X1 port map( B1 => n102, B2 => n7, A => B_23_port, ZN => 
                           E_23_port);
   U3 : XNOR2_X1 port map( A => n7, B => A(14), ZN => E_21_port);
   U4 : XNOR2_X1 port map( A => n11, B => D_18_port, ZN => E_18_port);
   U5 : NAND2_X1 port map( A1 => n11, A2 => n101, ZN => n10);
   U6 : NAND2_X1 port map( A1 => n90, A2 => n6, ZN => E_22_port);
   U7 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n13, ZN => n11);
   U8 : XNOR2_X1 port map( A => n87, B => A(10), ZN => E_17_port);
   U9 : NOR2_X1 port map( A1 => n13, A2 => A(9), ZN => n87);
   U10 : XNOR2_X1 port map( A => n88, B => A(6), ZN => E_13_port);
   U11 : NOR2_X1 port map( A1 => n17, A2 => A(5), ZN => n88);
   U12 : NOR2_X1 port map( A1 => n9, A2 => A(13), ZN => n7);
   U13 : BUF_X1 port map( A => A(15), Z => D_22_port);
   U14 : XNOR2_X1 port map( A => A(8), B => n16, ZN => E_15_port);
   U15 : NOR2_X1 port map( A1 => A(7), A2 => n15, ZN => n16);
   U16 : BUF_X1 port map( A => A(15), Z => B_23_port);
   U17 : XNOR2_X1 port map( A => A(4), B => n20, ZN => E_11_port);
   U18 : NOR2_X1 port map( A1 => A(3), A2 => n19, ZN => n20);
   U19 : OR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n19, ZN => n17);
   U20 : OR3_X1 port map( A1 => A(5), A2 => A(6), A3 => n17, ZN => n15);
   U21 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n15, ZN => n13);
   U22 : OR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n4);
   U23 : OR2_X1 port map( A1 => n10, A2 => A(12), ZN => n9);
   U29 : OR2_X1 port map( A1 => n4, A2 => A(2), ZN => n19);
   U32 : INV_X1 port map( A => E_23_port, ZN => n89);
   U35 : INV_X1 port map( A => E_23_port, ZN => n90);
   U36 : INV_X1 port map( A => n89, ZN => E_26_port);
   U37 : INV_X1 port map( A => n89, ZN => E_30_port);
   U38 : INV_X1 port map( A => n89, ZN => C_31_port);
   U39 : INV_X1 port map( A => n89, ZN => C_30_port);
   U40 : INV_X1 port map( A => n90, ZN => C_24_port);
   U41 : INV_X1 port map( A => n90, ZN => C_28_port);
   U42 : INV_X1 port map( A => n90, ZN => C_22_port);
   U43 : INV_X1 port map( A => n90, ZN => C_26_port);
   U44 : INV_X1 port map( A => n89, ZN => E_27_port);
   U45 : INV_X1 port map( A => n101, ZN => D_18_port);
   U46 : INV_X1 port map( A => A(11), ZN => n101);
   U47 : INV_X1 port map( A => A(14), ZN => n102);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S4 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S4;

architecture SYN_struct of shift_mul_N16_S4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_20_port, E_19_port, E_18_port, E_17_port, E_16_port,
      E_15_port, E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, 
      E_9_port, E_8_port, E_7_port, E_6_port, E_23_port, E_21_port, n6, n7, n8,
      n10, n12, n13, n14, n15, n16, n19, n21, n22, n24, n25, n105, n106, n107, 
      n108, n109, D_19_port, n111, D_20_port, B_19_port, n114 : std_logic;

begin
   B <= ( B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, 
      B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, 
      B_19_port, D_19_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6),
      A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   C <= ( E_21_port, E_21_port, E_21_port, E_21_port, E_23_port, E_23_port, 
      E_21_port, E_21_port, E_23_port, E_23_port, E_23_port, E_23_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   D <= ( D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, 
      D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, 
      D_19_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4)
      , A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   E <= ( E_23_port, E_23_port, E_23_port, E_21_port, E_23_port, E_23_port, 
      E_23_port, E_23_port, E_23_port, E_21_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U26 : XOR2_X1 port map( A => n6, B => A(4), Z => E_9_port);
   U27 : XOR2_X1 port map( A => n7, B => A(3), Z => E_8_port);
   U28 : XOR2_X1 port map( A => n8, B => n107, Z => E_7_port);
   U29 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_6_port);
   U30 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n114, ZN => n13);
   U32 : XOR2_X1 port map( A => A(12), B => n16, Z => E_17_port);
   U33 : XOR2_X1 port map( A => n15, B => n109, Z => E_16_port);
   U35 : XOR2_X1 port map( A => n19, B => A(9), Z => E_14_port);
   U36 : XOR2_X1 port map( A => n21, B => A(8), Z => E_13_port);
   U37 : XOR2_X1 port map( A => n22, B => n108, Z => E_12_port);
   U38 : XOR2_X1 port map( A => n24, B => A(5), Z => E_10_port);
   U2 : AOI21_X1 port map( B1 => n15, B2 => n14, A => n114, ZN => E_21_port);
   U3 : AOI21_X2 port map( B1 => n10, B2 => n111, A => n114, ZN => E_23_port);
   U4 : XNOR2_X1 port map( A => n10, B => D_19_port, ZN => E_19_port);
   U5 : NAND2_X1 port map( A1 => n15, A2 => n109, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n22, A2 => n108, ZN => n21);
   U7 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => E_20_port);
   U8 : INV_X1 port map( A => E_21_port, ZN => n12);
   U9 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n19, ZN => n15);
   U10 : NOR3_X1 port map( A1 => A(12), A2 => A(13), A3 => n16, ZN => n10);
   U11 : NOR4_X1 port map( A1 => A(11), A2 => A(12), A3 => A(13), A4 => 
                           D_19_port, ZN => n14);
   U12 : XNOR2_X1 port map( A => n105, B => A(13), ZN => E_18_port);
   U13 : NOR2_X1 port map( A1 => n16, A2 => A(12), ZN => n105);
   U14 : XNOR2_X1 port map( A => n106, B => A(10), ZN => E_15_port);
   U15 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n106);
   U16 : NOR3_X1 port map( A1 => A(5), A2 => A(6), A3 => n24, ZN => n22);
   U17 : BUF_X1 port map( A => A(15), Z => B_19_port);
   U18 : BUF_X1 port map( A => A(15), Z => D_20_port);
   U19 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n8);
   U20 : XNOR2_X1 port map( A => A(6), B => n25, ZN => E_11_port);
   U21 : NOR2_X1 port map( A1 => A(5), A2 => n24, ZN => n25);
   U22 : INV_X1 port map( A => A(7), ZN => n108);
   U23 : INV_X1 port map( A => A(11), ZN => n109);
   U24 : OR2_X1 port map( A1 => n6, A2 => A(4), ZN => n24);
   U25 : OR2_X1 port map( A1 => n21, A2 => A(8), ZN => n19);
   U31 : BUF_X1 port map( A => A(15), Z => n114);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n107, ZN => n7);
   U39 : OR2_X1 port map( A1 => n7, A2 => A(3), ZN => n6);
   U40 : INV_X1 port map( A => A(2), ZN => n107);
   U41 : INV_X1 port map( A => n111, ZN => D_19_port);
   U42 : INV_X1 port map( A => A(14), ZN => n111);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S2 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S2;

architecture SYN_struct of shift_mul_N16_S2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port,
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, C_22_port, n7, n8, n9, n11, n12, n15, n16, 
      n17, n18, n19, n20, n21, n23, n24, n26, n27, n28, E_23_port, n118, n119, 
      n120, D_13_port, n122, D_15_port, n124, D_18_port, D_30_port, B_29_port :
      std_logic;

begin
   B <= ( B_29_port, B_29_port, B_29_port, B_29_port, B_29_port, D_30_port, 
      D_30_port, D_30_port, D_30_port, D_30_port, D_30_port, D_30_port, 
      D_30_port, D_30_port, D_30_port, A(14), A(13), D_15_port, A(11), 
      D_13_port, A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port );
   C <= ( C_22_port, E_23_port, C_22_port, C_22_port, C_22_port, C_22_port, 
      C_22_port, E_23_port, C_22_port, C_22_port, E_23_port, E_23_port, 
      C_22_port, E_23_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, E_5_port, E_4_port, A(0), X_Logic0_port, 
      X_Logic0_port );
   D <= ( D_30_port, D_30_port, D_18_port, D_18_port, D_18_port, D_18_port, 
      D_18_port, D_18_port, D_18_port, D_18_port, D_18_port, D_18_port, 
      D_18_port, D_18_port, A(14), A(13), D_15_port, A(11), D_13_port, A(9), 
      A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   E <= ( C_22_port, C_22_port, E_23_port, C_22_port, E_23_port, E_23_port, 
      E_23_port, E_23_port, E_23_port, E_23_port, E_23_port, E_23_port, 
      E_23_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n7, B => A(6), Z => E_9_port);
   U28 : XOR2_X1 port map( A => n8, B => A(5), Z => E_8_port);
   U29 : XOR2_X1 port map( A => n9, B => n120, Z => E_7_port);
   U30 : XOR2_X1 port map( A => n11, B => A(3), Z => E_6_port);
   U31 : XOR2_X1 port map( A => n12, B => n119, Z => E_5_port);
   U32 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_4_port);
   U33 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => B_29_port, ZN => n15);
   U34 : XOR2_X1 port map( A => n20, B => A(13), Z => E_16_port);
   U35 : XOR2_X1 port map( A => n124, B => n21, Z => E_15_port);
   U36 : XOR2_X1 port map( A => n23, B => A(11), Z => E_14_port);
   U37 : XOR2_X1 port map( A => n122, B => n24, Z => E_13_port);
   U38 : XOR2_X1 port map( A => n26, B => A(9), Z => E_12_port);
   U39 : XOR2_X1 port map( A => n27, B => A(7), Z => E_10_port);
   U2 : INV_X1 port map( A => n118, ZN => E_23_port);
   U3 : INV_X1 port map( A => C_22_port, ZN => n118);
   U4 : AOI21_X1 port map( B1 => n17, B2 => n16, A => B_29_port, ZN => 
                           C_22_port);
   U5 : NAND2_X1 port map( A1 => n118, A2 => n15, ZN => E_18_port);
   U6 : INV_X1 port map( A => n16, ZN => n26);
   U7 : NAND2_X1 port map( A1 => n24, A2 => n122, ZN => n23);
   U8 : NAND2_X1 port map( A1 => n21, A2 => n124, ZN => n20);
   U9 : NAND2_X1 port map( A1 => n9, A2 => n120, ZN => n8);
   U10 : NOR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n27, ZN => n16);
   U11 : NOR4_X1 port map( A1 => A(11), A2 => D_15_port, A3 => D_13_port, A4 =>
                           n18, ZN => n17);
   U12 : OR3_X1 port map( A1 => A(13), A2 => A(9), A3 => A(14), ZN => n18);
   U13 : BUF_X1 port map( A => A(15), Z => D_18_port);
   U14 : BUF_X1 port map( A => A(15), Z => D_30_port);
   U15 : XNOR2_X1 port map( A => A(8), B => n28, ZN => E_11_port);
   U16 : NOR2_X1 port map( A1 => A(7), A2 => n27, ZN => n28);
   U17 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n12);
   U18 : XNOR2_X1 port map( A => A(14), B => n19, ZN => E_17_port);
   U19 : NOR2_X1 port map( A1 => A(13), A2 => n20, ZN => n19);
   U20 : NOR2_X1 port map( A1 => n26, A2 => A(9), ZN => n24);
   U21 : NOR2_X1 port map( A1 => n11, A2 => A(3), ZN => n9);
   U22 : NOR2_X1 port map( A1 => n23, A2 => A(11), ZN => n21);
   U23 : INV_X1 port map( A => A(12), ZN => n124);
   U24 : INV_X1 port map( A => A(10), ZN => n122);
   U25 : BUF_X1 port map( A => A(15), Z => B_29_port);
   U26 : INV_X1 port map( A => A(4), ZN => n120);
   U40 : OR2_X1 port map( A1 => n7, A2 => A(6), ZN => n27);
   U41 : NAND2_X1 port map( A1 => n12, A2 => n119, ZN => n11);
   U42 : OR2_X1 port map( A1 => n8, A2 => A(5), ZN => n7);
   U43 : INV_X1 port map( A => A(2), ZN => n119);
   U44 : INV_X1 port map( A => n122, ZN => D_13_port);
   U45 : INV_X1 port map( A => n124, ZN => D_15_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shift_mul_N16_S0 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S0;

architecture SYN_struct of shift_mul_N16_S0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_16_port, E_15_port, E_14_port, E_13_port, E_12_port,
      E_11_port, E_10_port, E_9_port, E_8_port, E_7_port, E_6_port, E_5_port, 
      E_3_port, E_2_port, net25272, E_4_port, n6, n8, n9, n10, n11, n12, n13, 
      n14, n16, n18, n19, n21, n22, n99, n100, C_20_port, D_3_port, n103, n104,
      D_12_port, n106, D_28_port, n108 : std_logic;

begin
   B <= ( A(15), D_28_port, D_28_port, D_28_port, A(15), D_28_port, D_28_port, 
      D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, 
      D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), A(12), 
      D_12_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), D_3_port, 
      A(1), A(0) );
   C <= ( C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, E_5_port, E_4_port, E_3_port, E_2_port, A(0) );
   D <= ( D_28_port, D_28_port, D_28_port, D_28_port, A(15), D_28_port, A(15), 
      D_28_port, A(15), D_28_port, A(15), D_28_port, A(15), D_28_port, A(15), 
      D_28_port, A(14), A(13), A(12), D_12_port, A(10), A(9), A(8), A(7), A(6),
      A(5), A(4), A(3), D_3_port, A(1), A(0), X_Logic0_port );
   E <= ( C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, E_3_port, E_2_port, A(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U29 : XOR2_X1 port map( A => n8, B => A(7), Z => E_8_port);
   U30 : XOR2_X1 port map( A => n9, B => A(6), Z => E_7_port);
   U31 : XOR2_X1 port map( A => n12, B => A(3), Z => E_4_port);
   U32 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_2_port);
   U34 : XOR2_X1 port map( A => n16, B => A(13), Z => E_14_port);
   U35 : XOR2_X1 port map( A => n18, B => A(12), Z => E_13_port);
   U36 : XOR2_X1 port map( A => n21, B => A(9), Z => E_10_port);
   U2 : BUF_X2 port map( A => net25272, Z => C_20_port);
   U3 : INV_X1 port map( A => n6, ZN => net25272);
   U4 : INV_X1 port map( A => n108, ZN => D_28_port);
   U5 : XNOR2_X1 port map( A => n19, B => D_12_port, ZN => E_12_port);
   U6 : XNOR2_X1 port map( A => n10, B => A(5), ZN => E_6_port);
   U7 : XNOR2_X1 port map( A => n13, B => D_3_port, ZN => E_3_port);
   U8 : OAI21_X1 port map( B1 => n14, B2 => n108, A => n6, ZN => E_16_port);
   U9 : NAND2_X1 port map( A1 => n10, A2 => n104, ZN => n9);
   U10 : NAND2_X1 port map( A1 => n19, A2 => n106, ZN => n18);
   U11 : NAND2_X1 port map( A1 => n108, A2 => n14, ZN => n6);
   U12 : NOR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n12, ZN => n10);
   U13 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n21, ZN => n19);
   U14 : XNOR2_X1 port map( A => n99, B => A(8), ZN => E_9_port);
   U15 : NOR2_X1 port map( A1 => n8, A2 => A(7), ZN => n99);
   U16 : XNOR2_X1 port map( A => n100, B => A(14), ZN => E_15_port);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(13), ZN => n100);
   U18 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n13);
   U19 : XNOR2_X1 port map( A => A(10), B => n22, ZN => E_11_port);
   U20 : NOR2_X1 port map( A1 => A(9), A2 => n21, ZN => n22);
   U21 : XNOR2_X1 port map( A => A(4), B => n11, ZN => E_5_port);
   U22 : NOR2_X1 port map( A1 => A(3), A2 => n12, ZN => n11);
   U23 : NAND2_X1 port map( A1 => n13, A2 => n103, ZN => n12);
   U24 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n8, ZN => n21);
   U25 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n16, ZN => n14);
   U26 : OR2_X1 port map( A1 => n18, A2 => A(12), ZN => n16);
   U27 : OR2_X1 port map( A1 => n9, A2 => A(6), ZN => n8);
   U28 : INV_X1 port map( A => n103, ZN => D_3_port);
   U33 : INV_X1 port map( A => A(2), ZN => n103);
   U37 : INV_X1 port map( A => A(5), ZN => n104);
   U38 : INV_X1 port map( A => n106, ZN => D_12_port);
   U39 : INV_X1 port map( A => A(11), ZN => n106);
   U40 : INV_X1 port map( A => A(15), ZN => n108);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity cla_adder_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end cla_adder_N32_0;

architecture SYN_struct of cla_adder_N32_0 is

   component sum_generator_Nbits32_Nblocks8_0
      port( A, B : in std_logic_vector (31 downto 0);  Carry : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_Nblocks8_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal Carry_8_port, Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port,
      Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port : std_logic;

begin
   
   CG : carry_generator_N32_Nblocks8_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci, Cout(8) => 
                           Carry_8_port, Cout(7) => Carry_7_port, Cout(6) => 
                           Carry_6_port, Cout(5) => Carry_5_port, Cout(4) => 
                           Carry_4_port, Cout(3) => Carry_3_port, Cout(2) => 
                           Carry_2_port, Cout(1) => Carry_1_port, Cout(0) => 
                           Carry_0_port);
   SG : sum_generator_Nbits32_Nblocks8_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Carry(8) => Carry_8_port, 
                           Carry(7) => Carry_7_port, Carry(6) => Carry_6_port, 
                           Carry(5) => Carry_5_port, Carry(4) => Carry_4_port, 
                           Carry(3) => Carry_3_port, Carry(2) => Carry_2_port, 
                           Carry(1) => Carry_1_port, Carry(0) => Carry_0_port, 
                           S(31) => Sum(31), S(30) => Sum(30), S(29) => Sum(29)
                           , S(28) => Sum(28), S(27) => Sum(27), S(26) => 
                           Sum(26), S(25) => Sum(25), S(24) => Sum(24), S(23) 
                           => Sum(23), S(22) => Sum(22), S(21) => Sum(21), 
                           S(20) => Sum(20), S(19) => Sum(19), S(18) => Sum(18)
                           , S(17) => Sum(17), S(16) => Sum(16), S(15) => 
                           Sum(15), S(14) => Sum(14), S(13) => Sum(13), S(12) 
                           => Sum(12), S(11) => Sum(11), S(10) => Sum(10), S(9)
                           => Sum(9), S(8) => Sum(8), S(7) => Sum(7), S(6) => 
                           Sum(6), S(5) => Sum(5), S(4) => Sum(4), S(3) => 
                           Sum(3), S(2) => Sum(2), S(1) => Sum(1), S(0) => 
                           Sum(0), Cout => Cout);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity generic_xor_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end generic_xor_N32;

architecture SYN_struct of generic_xor_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component xor_gate_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   X_gate_0 : xor_gate_0 port map( A => A(0), B => n3, Y => Y(0));
   X_gate_1 : xor_gate_31 port map( A => A(1), B => n1, Y => Y(1));
   X_gate_2 : xor_gate_30 port map( A => A(2), B => n1, Y => Y(2));
   X_gate_3 : xor_gate_29 port map( A => A(3), B => n1, Y => Y(3));
   X_gate_4 : xor_gate_28 port map( A => A(4), B => n1, Y => Y(4));
   X_gate_5 : xor_gate_27 port map( A => A(5), B => n1, Y => Y(5));
   X_gate_6 : xor_gate_26 port map( A => A(6), B => n1, Y => Y(6));
   X_gate_7 : xor_gate_25 port map( A => A(7), B => n1, Y => Y(7));
   X_gate_8 : xor_gate_24 port map( A => A(8), B => n1, Y => Y(8));
   X_gate_9 : xor_gate_23 port map( A => A(9), B => n1, Y => Y(9));
   X_gate_10 : xor_gate_22 port map( A => A(10), B => n1, Y => Y(10));
   X_gate_11 : xor_gate_21 port map( A => A(11), B => n1, Y => Y(11));
   X_gate_12 : xor_gate_20 port map( A => A(12), B => n1, Y => Y(12));
   X_gate_13 : xor_gate_19 port map( A => A(13), B => n2, Y => Y(13));
   X_gate_14 : xor_gate_18 port map( A => A(14), B => n2, Y => Y(14));
   X_gate_15 : xor_gate_17 port map( A => A(15), B => n2, Y => Y(15));
   X_gate_16 : xor_gate_16 port map( A => A(16), B => n2, Y => Y(16));
   X_gate_17 : xor_gate_15 port map( A => A(17), B => n2, Y => Y(17));
   X_gate_18 : xor_gate_14 port map( A => A(18), B => n2, Y => Y(18));
   X_gate_19 : xor_gate_13 port map( A => A(19), B => n2, Y => Y(19));
   X_gate_20 : xor_gate_12 port map( A => A(20), B => n2, Y => Y(20));
   X_gate_21 : xor_gate_11 port map( A => A(21), B => n2, Y => Y(21));
   X_gate_22 : xor_gate_10 port map( A => A(22), B => n2, Y => Y(22));
   X_gate_23 : xor_gate_9 port map( A => A(23), B => n2, Y => Y(23));
   X_gate_24 : xor_gate_8 port map( A => A(24), B => n2, Y => Y(24));
   X_gate_25 : xor_gate_7 port map( A => A(25), B => n3, Y => Y(25));
   X_gate_26 : xor_gate_6 port map( A => A(26), B => n3, Y => Y(26));
   X_gate_27 : xor_gate_5 port map( A => A(27), B => n3, Y => Y(27));
   X_gate_28 : xor_gate_4 port map( A => A(28), B => n3, Y => Y(28));
   X_gate_29 : xor_gate_3 port map( A => A(29), B => n3, Y => Y(29));
   X_gate_30 : xor_gate_2 port map( A => A(30), B => n3, Y => Y(30));
   X_gate_31 : xor_gate_1 port map( A => A(31), B => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : BUF_X1 port map( A => B, Z => n2);
   U3 : BUF_X1 port map( A => B, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity counter_DW01_dec_0 is

   port( A : in std_logic_vector (30 downto 0);  SUM : out std_logic_vector (30
         downto 0));

end counter_DW01_dec_0;

architecture SYN_rpl of counter_DW01_dec_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, 
      SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, 
      SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, 
      SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, SUM_11_port, 
      SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port, 
      SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n20,
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n60, n61, n62, n63, n65, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88 : std_logic;

begin
   SUM <= ( SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, 
      SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, 
      SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, 
      SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, SUM_11_port, 
      SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port, 
      SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U48 : XOR2_X1 port map( A => A(30), B => n34, Z => SUM_30_port);
   U3 : OR2_X2 port map( A1 => n29, A2 => A(6), ZN => n1);
   U1 : OR2_X1 port map( A1 => n6, A2 => A(4), ZN => n7);
   U2 : OR2_X1 port map( A1 => n38, A2 => A(3), ZN => n6);
   U4 : AND2_X1 port map( A1 => n2, A2 => n3, ZN => n69);
   U5 : INV_X1 port map( A => n12, ZN => n57);
   U6 : INV_X1 port map( A => n50, ZN => n51);
   U7 : NAND2_X1 port map( A1 => n57, A2 => n15, ZN => n14);
   U8 : OR2_X1 port map( A1 => n77, A2 => n5, ZN => n73);
   U9 : AND2_X1 port map( A1 => n52, A2 => n53, ZN => n50);
   U10 : OAI21_X1 port map( B1 => n57, B2 => n15, A => n14, ZN => SUM_20_port);
   U11 : INV_X1 port map( A => A(6), ZN => n26);
   U12 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n54, ZN => SUM_21_port);
   U13 : INV_X1 port map( A => A(21), ZN => n56);
   U14 : INV_X1 port map( A => n14, ZN => n55);
   U15 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n73, ZN => SUM_12_port);
   U16 : INV_X1 port map( A => A(12), ZN => n75);
   U17 : NOR2_X1 port map( A1 => n77, A2 => A(11), ZN => n74);
   U18 : NOR2_X1 port map( A1 => n73, A2 => A(13), ZN => n71);
   U19 : NOR2_X1 port map( A1 => n14, A2 => A(21), ZN => n52);
   U20 : INV_X1 port map( A => n76, ZN => SUM_11_port);
   U21 : AOI21_X1 port map( B1 => n77, B2 => A(11), A => n74, ZN => n76);
   U22 : AND2_X1 port map( A1 => n79, A2 => n80, ZN => n60);
   U23 : NOR2_X1 port map( A1 => n10, A2 => A(16), ZN => n79);
   U24 : NOR2_X1 port map( A1 => A(18), A2 => A(17), ZN => n80);
   U25 : NOR2_X1 port map( A1 => n42, A2 => A(27), ZN => n39);
   U26 : NOR2_X1 port map( A1 => n1, A2 => A(7), ZN => n22);
   U27 : NOR2_X1 port map( A1 => n87, A2 => A(17), ZN => n62);
   U28 : OR2_X1 port map( A1 => n16, A2 => A(24), ZN => n81);
   U29 : NOR2_X1 port map( A1 => A(29), A2 => n35, ZN => n34);
   U30 : NOR2_X1 port map( A1 => A(14), A2 => A(13), ZN => n3);
   U31 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n2);
   U32 : OR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n88);
   U33 : INV_X1 port map( A => n45, ZN => SUM_25_port);
   U34 : INV_X1 port map( A => n41, ZN => SUM_27_port);
   U35 : INV_X1 port map( A => A(20), ZN => n15);
   U36 : NOR2_X1 port map( A1 => n82, A2 => n83, ZN => n43);
   U37 : NAND2_X1 port map( A1 => n50, A2 => n17, ZN => n82);
   U38 : OR2_X1 port map( A1 => A(25), A2 => A(24), ZN => n83);
   U39 : OAI21_X1 port map( B1 => n47, B2 => n48, A => n81, ZN => SUM_24_port);
   U40 : INV_X1 port map( A => A(24), ZN => n48);
   U41 : INV_X1 port map( A => A(10), ZN => n78);
   U42 : INV_X1 port map( A => A(16), ZN => n68);
   U43 : OR2_X1 port map( A1 => A(12), A2 => A(11), ZN => n5);
   U44 : INV_X1 port map( A => A(17), ZN => n65);
   U45 : OAI21_X1 port map( B1 => n71, B2 => n9, A => n70, ZN => SUM_14_port);
   U46 : INV_X1 port map( A => A(14), ZN => n9);
   U47 : INV_X1 port map( A => n69, ZN => n70);
   U49 : INV_X1 port map( A => A(8), ZN => n23);
   U50 : INV_X1 port map( A => n24, ZN => SUM_7_port);
   U51 : INV_X1 port map( A => n19, ZN => SUM_9_port);
   U52 : INV_X1 port map( A => n72, ZN => SUM_13_port);
   U53 : AOI21_X1 port map( B1 => n73, B2 => A(13), A => n71, ZN => n72);
   U54 : INV_X1 port map( A => A(18), ZN => n8);
   U55 : INV_X1 port map( A => A(22), ZN => n53);
   U56 : INV_X1 port map( A => A(19), ZN => n13);
   U57 : INV_X1 port map( A => A(15), ZN => n11);
   U58 : INV_X1 port map( A => A(1), ZN => n58);
   U59 : INV_X1 port map( A => A(3), ZN => n33);
   U60 : INV_X1 port map( A => A(5), ZN => n28);
   U61 : INV_X1 port map( A => n7, ZN => n27);
   U62 : INV_X1 port map( A => A(2), ZN => n37);
   U63 : INV_X1 port map( A => n88, ZN => n36);
   U64 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n7, ZN => SUM_4_port);
   U65 : INV_X1 port map( A => A(4), ZN => n31);
   U66 : INV_X1 port map( A => n6, ZN => n30);
   U67 : INV_X1 port map( A => A(23), ZN => n17);
   U68 : INV_X1 port map( A => A(28), ZN => n40);
   U69 : INV_X1 port map( A => A(26), ZN => n44);
   U70 : OAI21_X1 port map( B1 => n39, B2 => n40, A => n35, ZN => SUM_28_port);
   U71 : OAI21_X1 port map( B1 => n60, B2 => n13, A => n12, ZN => SUM_19_port);
   U72 : INV_X1 port map( A => n60, ZN => n61);
   U73 : AOI21_X1 port map( B1 => n42, B2 => A(27), A => n39, ZN => n41);
   U74 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n35);
   U75 : OAI21_X1 port map( B1 => SUM_0_port, B2 => n58, A => n88, ZN => 
                           SUM_1_port);
   U76 : OR2_X1 port map( A1 => n10, A2 => A(16), ZN => n87);
   U77 : NOR2_X1 port map( A1 => n88, A2 => A(2), ZN => n32);
   U78 : NOR2_X1 port map( A1 => n7, A2 => A(5), ZN => n25);
   U79 : NAND2_X1 port map( A1 => n60, A2 => n13, ZN => n12);
   U80 : NOR2_X1 port map( A1 => n1, A2 => A(7), ZN => n84);
   U81 : AND2_X2 port map( A1 => n84, A2 => n85, ZN => n21);
   U82 : AND2_X1 port map( A1 => n86, A2 => n23, ZN => n85);
   U83 : INV_X1 port map( A => A(9), ZN => n86);
   U84 : XNOR2_X1 port map( A => A(29), B => n35, ZN => SUM_29_port);
   U85 : NAND2_X1 port map( A1 => n69, A2 => n11, ZN => n10);
   U86 : OAI21_X1 port map( B1 => n69, B2 => n11, A => n10, ZN => SUM_15_port);
   U87 : OAI21_X1 port map( B1 => n43, B2 => n44, A => n42, ZN => SUM_26_port);
   U88 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n6, ZN => SUM_3_port);
   U89 : INV_X1 port map( A => n10, ZN => n67);
   U90 : AOI21_X1 port map( B1 => n81, B2 => A(25), A => n43, ZN => n45);
   U91 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n42);
   U92 : INV_X1 port map( A => n32, ZN => n38);
   U93 : NAND2_X1 port map( A1 => n50, A2 => n17, ZN => n16);
   U94 : OAI21_X1 port map( B1 => n25, B2 => n26, A => n1, ZN => SUM_6_port);
   U95 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n87, ZN => SUM_16_port);
   U96 : OAI21_X1 port map( B1 => n50, B2 => n17, A => n16, ZN => SUM_23_port);
   U97 : OAI21_X1 port map( B1 => n27, B2 => n28, A => n29, ZN => SUM_5_port);
   U98 : INV_X1 port map( A => n16, ZN => n47);
   U99 : INV_X1 port map( A => n25, ZN => n29);
   U100 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => SUM_2_port);
   U101 : OAI21_X1 port map( B1 => n79, B2 => n65, A => n63, ZN => SUM_17_port)
                           ;
   U102 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U103 : OAI21_X1 port map( B1 => n22, B2 => n23, A => n20, ZN => SUM_8_port);
   U104 : OAI21_X1 port map( B1 => n62, B2 => n8, A => n61, ZN => SUM_18_port);
   U105 : INV_X1 port map( A => n62, ZN => n63);
   U106 : OAI21_X1 port map( B1 => n52, B2 => n53, A => n51, ZN => SUM_22_port)
                           ;
   U107 : AOI21_X1 port map( B1 => n20, B2 => A(9), A => n21, ZN => n19);
   U108 : AOI21_X1 port map( B1 => n1, B2 => A(7), A => n22, ZN => n24);
   U109 : OAI21_X1 port map( B1 => n21, B2 => n78, A => n77, ZN => SUM_10_port)
                           ;
   U110 : INV_X1 port map( A => n52, ZN => n54);
   U111 : NAND2_X1 port map( A1 => n21, A2 => n78, ZN => n77);
   U112 : NAND2_X1 port map( A1 => n21, A2 => n78, ZN => n4);
   U113 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n20);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PC_incr_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end PC_incr_DW01_add_1;

architecture SYN_cla of PC_incr_DW01_add_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, SUM_2_port, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U5 : XOR2_X1 port map( A => A(28), B => n13, Z => SUM_28_port);
   U6 : XOR2_X1 port map( A => A(27), B => n14, Z => SUM_27_port);
   U7 : XOR2_X1 port map( A => A(26), B => n15, Z => SUM_26_port);
   U8 : XOR2_X1 port map( A => A(25), B => n16, Z => SUM_25_port);
   U9 : XOR2_X1 port map( A => A(24), B => n17, Z => SUM_24_port);
   U10 : XOR2_X1 port map( A => A(23), B => n18, Z => SUM_23_port);
   U11 : XOR2_X1 port map( A => A(21), B => n19, Z => SUM_21_port);
   U12 : XOR2_X1 port map( A => A(20), B => n21, Z => SUM_20_port);
   U13 : XOR2_X1 port map( A => A(19), B => n22, Z => SUM_19_port);
   U14 : XOR2_X1 port map( A => A(18), B => n23, Z => SUM_18_port);
   U15 : XOR2_X1 port map( A => A(29), B => n11, Z => SUM_29_port);
   U16 : XOR2_X1 port map( A => n10, B => A(30), Z => SUM_30_port);
   U34 : XOR2_X1 port map( A => A(7), B => n6, Z => SUM_7_port);
   U35 : XOR2_X1 port map( A => A(17), B => n24, Z => SUM_17_port);
   U36 : XOR2_X1 port map( A => A(13), B => n40, Z => SUM_13_port);
   U37 : XOR2_X1 port map( A => A(12), B => n43, Z => SUM_12_port);
   U38 : XOR2_X1 port map( A => n2, B => A(16), Z => SUM_16_port);
   U39 : XOR2_X1 port map( A => A(10), B => n46, Z => SUM_10_port);
   U40 : XOR2_X1 port map( A => A(9), B => n4, Z => SUM_9_port);
   U41 : XOR2_X1 port map( A => A(8), B => n5, Z => SUM_8_port);
   U42 : XOR2_X1 port map( A => A(5), B => n7, Z => SUM_5_port);
   U43 : XOR2_X1 port map( A => A(4), B => n33, Z => SUM_4_port);
   U2 : INV_X1 port map( A => n33, ZN => n8);
   U3 : INV_X1 port map( A => n5, ZN => n44);
   U4 : XNOR2_X1 port map( A => n41, B => n38, ZN => SUM_14_port);
   U17 : NOR2_X1 port map( A1 => n50, A2 => SUM_2_port, ZN => n33);
   U18 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => n38);
   U19 : INV_X1 port map( A => n40, ZN => n39);
   U20 : NOR2_X1 port map( A1 => n8, A2 => n34, ZN => n5);
   U21 : NOR2_X1 port map( A1 => n44, A2 => n31, ZN => n43);
   U22 : NOR2_X1 port map( A1 => n29, A2 => n42, ZN => n40);
   U23 : INV_X1 port map( A => n43, ZN => n42);
   U24 : NOR2_X1 port map( A1 => n30, A2 => n31, ZN => n27);
   U25 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => n30);
   U26 : INV_X1 port map( A => n34, ZN => n32);
   U27 : XOR2_X1 port map( A => n51, B => A(15), Z => SUM_15_port);
   U28 : AND2_X1 port map( A1 => n38, A2 => A(14), ZN => n51);
   U29 : XNOR2_X1 port map( A => n1, B => A(6), ZN => SUM_6_port);
   U30 : XNOR2_X1 port map( A => n45, B => A(11), ZN => SUM_11_port);
   U31 : NAND2_X1 port map( A1 => n46, A2 => A(10), ZN => n45);
   U32 : XNOR2_X1 port map( A => n9, B => A(31), ZN => SUM_31_port);
   U33 : NAND2_X1 port map( A1 => n10, A2 => A(30), ZN => n9);
   U44 : XNOR2_X1 port map( A => A(22), B => n3, ZN => SUM_22_port);
   U45 : NAND4_X1 port map( A1 => A(7), A2 => A(6), A3 => A(5), A4 => A(4), ZN 
                           => n34);
   U46 : NAND4_X1 port map( A1 => A(11), A2 => A(10), A3 => A(9), A4 => A(8), 
                           ZN => n31);
   U47 : NOR2_X1 port map( A1 => n8, A2 => n48, ZN => n7);
   U48 : INV_X1 port map( A => A(4), ZN => n48);
   U49 : NOR2_X1 port map( A1 => n20, A2 => n3, ZN => n18);
   U50 : INV_X1 port map( A => A(22), ZN => n20);
   U51 : NOR2_X1 port map( A1 => n44, A2 => n47, ZN => n4);
   U52 : INV_X1 port map( A => A(8), ZN => n47);
   U53 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U54 : NAND2_X1 port map( A1 => A(21), A2 => n19, ZN => n3);
   U55 : NAND2_X1 port map( A1 => A(5), A2 => n7, ZN => n1);
   U56 : NOR2_X1 port map( A1 => n49, A2 => n1, ZN => n6);
   U57 : INV_X1 port map( A => A(6), ZN => n49);
   U58 : INV_X1 port map( A => A(3), ZN => n50);
   U59 : INV_X1 port map( A => A(14), ZN => n41);
   U60 : AND2_X1 port map( A1 => A(20), A2 => n21, ZN => n19);
   U61 : AND2_X1 port map( A1 => n4, A2 => A(9), ZN => n46);
   U62 : INV_X1 port map( A => A(13), ZN => n35);
   U63 : INV_X1 port map( A => A(12), ZN => n29);
   U64 : AND2_X1 port map( A1 => A(29), A2 => n11, ZN => n10);
   U65 : AND2_X1 port map( A1 => A(23), A2 => n18, ZN => n17);
   U66 : AND2_X1 port map( A1 => A(16), A2 => n2, ZN => n24);
   U67 : AND2_X1 port map( A1 => A(17), A2 => n24, ZN => n23);
   U68 : AND2_X1 port map( A1 => A(18), A2 => n23, ZN => n22);
   U69 : AND2_X1 port map( A1 => A(19), A2 => n22, ZN => n21);
   U70 : AND2_X1 port map( A1 => A(24), A2 => n17, ZN => n16);
   U71 : AND2_X1 port map( A1 => A(25), A2 => n16, ZN => n15);
   U72 : AND2_X1 port map( A1 => A(26), A2 => n15, ZN => n14);
   U73 : AND2_X1 port map( A1 => A(27), A2 => n14, ZN => n13);
   U74 : AND2_X1 port map( A1 => A(28), A2 => n13, ZN => n11);
   U75 : AND2_X1 port map( A1 => n25, A2 => A(15), ZN => n2);
   U76 : NOR2_X1 port map( A1 => n26, A2 => n41, ZN => n25);
   U77 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => n26);
   U78 : NOR2_X1 port map( A1 => n29, A2 => n35, ZN => n28);
   U79 : XNOR2_X1 port map( A => A(2), B => n50, ZN => SUM_3_port);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_665 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_664 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0 is

   port( A : in std_logic_vector (5 downto 0);  SUM : out std_logic_vector (5 
         downto 0));

end w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0;

architecture SYN_rpl of w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_5_port, B => A(5), Z => SUM(5));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity w_reg_file_M8_N8_F4_Nbit32_DW01_add_1 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end w_reg_file_M8_N8_F4_Nbit32_DW01_add_1;

architecture SYN_rpl of w_reg_file_M8_N8_F4_Nbit32_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port 
      : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : XOR2_X1 port map( A => B(5), B => carry_5_port, Z => SUM(5));
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity w_reg_file_M8_N8_F4_Nbit32_DW01_add_0 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end w_reg_file_M8_N8_F4_Nbit32_DW01_add_0;

architecture SYN_rpl of w_reg_file_M8_N8_F4_Nbit32_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port 
      : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : XOR2_X1 port map( A => B(5), B => carry_5_port, Z => SUM(5));
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity sum_generator_Nbits32_Nblocks8 is

   port( A, B : in std_logic_vector (31 downto 0);  Carry : in std_logic_vector
         (8 downto 0);  S : out std_logic_vector (31 downto 0);  Cout : out 
         std_logic);

end sum_generator_Nbits32_Nblocks8;

architecture SYN_STRUCTURAL of sum_generator_Nbits32_Nblocks8 is

   component carry_select_N4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(8);
   
   CS_0 : carry_select_N4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Carry(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), 
                           A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), Ci => Carry(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9),
                           A(0) => A(8), B(3) => B(11), B(2) => B(10), B(1) => 
                           B(9), B(0) => B(8), Ci => Carry(2), S(3) => S(11), 
                           S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13)
                           , A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) 
                           => B(13), B(0) => B(12), Ci => Carry(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CS_4 : carry_select_N4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17)
                           , A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) 
                           => B(17), B(0) => B(16), Ci => Carry(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CS_5 : carry_select_N4 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21)
                           , A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) 
                           => B(21), B(0) => B(20), Ci => Carry(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CS_6 : carry_select_N4 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25)
                           , A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) 
                           => B(25), B(0) => B(24), Ci => Carry(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CS_7 : carry_select_N4 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29)
                           , A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) 
                           => B(29), B(0) => B(28), Ci => Carry(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity carry_generator_N32_Nblocks8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_Nblocks8;

architecture SYN_STRUCTURAL of carry_generator_N32_Nblocks8 is

   component G
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PGnet_block
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   signal Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, g_cin, p_cin, Gsignal_1_31_port, 
      Gsignal_1_30_port, Gsignal_1_29_port, Gsignal_1_28_port, 
      Gsignal_1_27_port, Gsignal_1_26_port, Gsignal_1_25_port, 
      Gsignal_1_24_port, Gsignal_1_23_port, Gsignal_1_22_port, 
      Gsignal_1_21_port, Gsignal_1_20_port, Gsignal_1_19_port, 
      Gsignal_1_18_port, Gsignal_1_17_port, Gsignal_1_16_port, 
      Gsignal_1_15_port, Gsignal_1_14_port, Gsignal_1_13_port, 
      Gsignal_1_12_port, Gsignal_1_11_port, Gsignal_1_10_port, Gsignal_1_9_port
      , Gsignal_1_8_port, Gsignal_1_7_port, Gsignal_1_6_port, Gsignal_1_5_port,
      Gsignal_1_4_port, Gsignal_1_3_port, Gsignal_1_2_port, Gsignal_1_1_port, 
      Gsignal_1_0_port, Gsignal_2_31_port, Gsignal_2_29_port, Gsignal_2_27_port
      , Gsignal_2_25_port, Gsignal_2_23_port, Gsignal_2_21_port, 
      Gsignal_2_19_port, Gsignal_2_17_port, Gsignal_2_15_port, 
      Gsignal_2_13_port, Gsignal_2_11_port, Gsignal_2_9_port, Gsignal_2_7_port,
      Gsignal_2_5_port, Gsignal_2_3_port, Gsignal_2_1_port, Gsignal_3_31_port, 
      Gsignal_3_27_port, Gsignal_3_23_port, Gsignal_3_19_port, 
      Gsignal_3_15_port, Gsignal_3_11_port, Gsignal_3_7_port, Gsignal_4_31_port
      , Gsignal_4_23_port, Gsignal_4_15_port, Gsignal_5_31_port, 
      Gsignal_5_27_port, Psignal_1_31_port, Psignal_1_30_port, 
      Psignal_1_29_port, Psignal_1_28_port, Psignal_1_27_port, 
      Psignal_1_26_port, Psignal_1_25_port, Psignal_1_24_port, 
      Psignal_1_23_port, Psignal_1_22_port, Psignal_1_21_port, 
      Psignal_1_20_port, Psignal_1_19_port, Psignal_1_18_port, 
      Psignal_1_17_port, Psignal_1_16_port, Psignal_1_15_port, 
      Psignal_1_14_port, Psignal_1_13_port, Psignal_1_12_port, 
      Psignal_1_11_port, Psignal_1_10_port, Psignal_1_9_port, Psignal_1_8_port,
      Psignal_1_7_port, Psignal_1_6_port, Psignal_1_5_port, Psignal_1_4_port, 
      Psignal_1_3_port, Psignal_1_2_port, Psignal_1_1_port, Psignal_2_31_port, 
      Psignal_2_29_port, Psignal_2_27_port, Psignal_2_25_port, 
      Psignal_2_23_port, Psignal_2_21_port, Psignal_2_19_port, 
      Psignal_2_17_port, Psignal_2_15_port, Psignal_2_13_port, 
      Psignal_2_11_port, Psignal_2_9_port, Psignal_2_7_port, Psignal_2_5_port, 
      Psignal_2_3_port, Psignal_3_31_port, Psignal_3_27_port, Psignal_3_23_port
      , Psignal_3_19_port, Psignal_3_15_port, Psignal_3_11_port, 
      Psignal_3_7_port, Psignal_4_31_port, Psignal_4_23_port, Psignal_4_15_port
      , Psignal_5_31_port, Psignal_5_27_port : std_logic;

begin
   Cout <= ( Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, Ci );
   
   PGnet_Cin_0 : PGnet_block port map( A => A(0), B => B(0), pout => p_cin, 
                           gout => g_cin);
   GCin_0 : G port map( gleft => g_cin, gright => Ci, pleft => p_cin, gout => 
                           Gsignal_1_0_port);
   PGnet_1 : PGnet_block port map( A => A(1), B => B(1), pout => 
                           Psignal_1_1_port, gout => Gsignal_1_1_port);
   PGnet_2 : PGnet_block port map( A => A(2), B => B(2), pout => 
                           Psignal_1_2_port, gout => Gsignal_1_2_port);
   PGnet_3 : PGnet_block port map( A => A(3), B => B(3), pout => 
                           Psignal_1_3_port, gout => Gsignal_1_3_port);
   PGnet_4 : PGnet_block port map( A => A(4), B => B(4), pout => 
                           Psignal_1_4_port, gout => Gsignal_1_4_port);
   PGnet_5 : PGnet_block port map( A => A(5), B => B(5), pout => 
                           Psignal_1_5_port, gout => Gsignal_1_5_port);
   PGnet_6 : PGnet_block port map( A => A(6), B => B(6), pout => 
                           Psignal_1_6_port, gout => Gsignal_1_6_port);
   PGnet_7 : PGnet_block port map( A => A(7), B => B(7), pout => 
                           Psignal_1_7_port, gout => Gsignal_1_7_port);
   PGnet_8 : PGnet_block port map( A => A(8), B => B(8), pout => 
                           Psignal_1_8_port, gout => Gsignal_1_8_port);
   PGnet_9 : PGnet_block port map( A => A(9), B => B(9), pout => 
                           Psignal_1_9_port, gout => Gsignal_1_9_port);
   PGnet_10 : PGnet_block port map( A => A(10), B => B(10), pout => 
                           Psignal_1_10_port, gout => Gsignal_1_10_port);
   PGnet_11 : PGnet_block port map( A => A(11), B => B(11), pout => 
                           Psignal_1_11_port, gout => Gsignal_1_11_port);
   PGnet_12 : PGnet_block port map( A => A(12), B => B(12), pout => 
                           Psignal_1_12_port, gout => Gsignal_1_12_port);
   PGnet_13 : PGnet_block port map( A => A(13), B => B(13), pout => 
                           Psignal_1_13_port, gout => Gsignal_1_13_port);
   PGnet_14 : PGnet_block port map( A => A(14), B => B(14), pout => 
                           Psignal_1_14_port, gout => Gsignal_1_14_port);
   PGnet_15 : PGnet_block port map( A => A(15), B => B(15), pout => 
                           Psignal_1_15_port, gout => Gsignal_1_15_port);
   PGnet_16 : PGnet_block port map( A => A(16), B => B(16), pout => 
                           Psignal_1_16_port, gout => Gsignal_1_16_port);
   PGnet_17 : PGnet_block port map( A => A(17), B => B(17), pout => 
                           Psignal_1_17_port, gout => Gsignal_1_17_port);
   PGnet_18 : PGnet_block port map( A => A(18), B => B(18), pout => 
                           Psignal_1_18_port, gout => Gsignal_1_18_port);
   PGnet_19 : PGnet_block port map( A => A(19), B => B(19), pout => 
                           Psignal_1_19_port, gout => Gsignal_1_19_port);
   PGnet_20 : PGnet_block port map( A => A(20), B => B(20), pout => 
                           Psignal_1_20_port, gout => Gsignal_1_20_port);
   PGnet_21 : PGnet_block port map( A => A(21), B => B(21), pout => 
                           Psignal_1_21_port, gout => Gsignal_1_21_port);
   PGnet_22 : PGnet_block port map( A => A(22), B => B(22), pout => 
                           Psignal_1_22_port, gout => Gsignal_1_22_port);
   PGnet_23 : PGnet_block port map( A => A(23), B => B(23), pout => 
                           Psignal_1_23_port, gout => Gsignal_1_23_port);
   PGnet_24 : PGnet_block port map( A => A(24), B => B(24), pout => 
                           Psignal_1_24_port, gout => Gsignal_1_24_port);
   PGnet_25 : PGnet_block port map( A => A(25), B => B(25), pout => 
                           Psignal_1_25_port, gout => Gsignal_1_25_port);
   PGnet_26 : PGnet_block port map( A => A(26), B => B(26), pout => 
                           Psignal_1_26_port, gout => Gsignal_1_26_port);
   PGnet_27 : PGnet_block port map( A => A(27), B => B(27), pout => 
                           Psignal_1_27_port, gout => Gsignal_1_27_port);
   PGnet_28 : PGnet_block port map( A => A(28), B => B(28), pout => 
                           Psignal_1_28_port, gout => Gsignal_1_28_port);
   PGnet_29 : PGnet_block port map( A => A(29), B => B(29), pout => 
                           Psignal_1_29_port, gout => Gsignal_1_29_port);
   PGnet_30 : PGnet_block port map( A => A(30), B => B(30), pout => 
                           Psignal_1_30_port, gout => Gsignal_1_30_port);
   PGnet_31 : PGnet_block port map( A => A(31), B => B(31), pout => 
                           Psignal_1_31_port, gout => Gsignal_1_31_port);
   Gblock_1_1 : G port map( gleft => Gsignal_1_1_port, gright => 
                           Gsignal_1_0_port, pleft => Psignal_1_1_port, gout =>
                           Gsignal_2_1_port);
   PGblock_1_3 : PG port map( gleft => Gsignal_1_3_port, gright => 
                           Gsignal_1_2_port, pleft => Psignal_1_3_port, pright 
                           => Psignal_1_2_port, pout => Psignal_2_3_port, gout 
                           => Gsignal_2_3_port);
   PGblock_1_5 : PG port map( gleft => Gsignal_1_5_port, gright => 
                           Gsignal_1_4_port, pleft => Psignal_1_5_port, pright 
                           => Psignal_1_4_port, pout => Psignal_2_5_port, gout 
                           => Gsignal_2_5_port);
   PGblock_1_7 : PG port map( gleft => Gsignal_1_7_port, gright => 
                           Gsignal_1_6_port, pleft => Psignal_1_7_port, pright 
                           => Psignal_1_6_port, pout => Psignal_2_7_port, gout 
                           => Gsignal_2_7_port);
   PGblock_1_9 : PG port map( gleft => Gsignal_1_9_port, gright => 
                           Gsignal_1_8_port, pleft => Psignal_1_9_port, pright 
                           => Psignal_1_8_port, pout => Psignal_2_9_port, gout 
                           => Gsignal_2_9_port);
   PGblock_1_11 : PG port map( gleft => Gsignal_1_11_port, gright => 
                           Gsignal_1_10_port, pleft => Psignal_1_11_port, 
                           pright => Psignal_1_10_port, pout => 
                           Psignal_2_11_port, gout => Gsignal_2_11_port);
   PGblock_1_13 : PG port map( gleft => Gsignal_1_13_port, gright => 
                           Gsignal_1_12_port, pleft => Psignal_1_13_port, 
                           pright => Psignal_1_12_port, pout => 
                           Psignal_2_13_port, gout => Gsignal_2_13_port);
   PGblock_1_15 : PG port map( gleft => Gsignal_1_15_port, gright => 
                           Gsignal_1_14_port, pleft => Psignal_1_15_port, 
                           pright => Psignal_1_14_port, pout => 
                           Psignal_2_15_port, gout => Gsignal_2_15_port);
   PGblock_1_17 : PG port map( gleft => Gsignal_1_17_port, gright => 
                           Gsignal_1_16_port, pleft => Psignal_1_17_port, 
                           pright => Psignal_1_16_port, pout => 
                           Psignal_2_17_port, gout => Gsignal_2_17_port);
   PGblock_1_19 : PG port map( gleft => Gsignal_1_19_port, gright => 
                           Gsignal_1_18_port, pleft => Psignal_1_19_port, 
                           pright => Psignal_1_18_port, pout => 
                           Psignal_2_19_port, gout => Gsignal_2_19_port);
   PGblock_1_21 : PG port map( gleft => Gsignal_1_21_port, gright => 
                           Gsignal_1_20_port, pleft => Psignal_1_21_port, 
                           pright => Psignal_1_20_port, pout => 
                           Psignal_2_21_port, gout => Gsignal_2_21_port);
   PGblock_1_23 : PG port map( gleft => Gsignal_1_23_port, gright => 
                           Gsignal_1_22_port, pleft => Psignal_1_23_port, 
                           pright => Psignal_1_22_port, pout => 
                           Psignal_2_23_port, gout => Gsignal_2_23_port);
   PGblock_1_25 : PG port map( gleft => Gsignal_1_25_port, gright => 
                           Gsignal_1_24_port, pleft => Psignal_1_25_port, 
                           pright => Psignal_1_24_port, pout => 
                           Psignal_2_25_port, gout => Gsignal_2_25_port);
   PGblock_1_27 : PG port map( gleft => Gsignal_1_27_port, gright => 
                           Gsignal_1_26_port, pleft => Psignal_1_27_port, 
                           pright => Psignal_1_26_port, pout => 
                           Psignal_2_27_port, gout => Gsignal_2_27_port);
   PGblock_1_29 : PG port map( gleft => Gsignal_1_29_port, gright => 
                           Gsignal_1_28_port, pleft => Psignal_1_29_port, 
                           pright => Psignal_1_28_port, pout => 
                           Psignal_2_29_port, gout => Gsignal_2_29_port);
   PGblock_1_31 : PG port map( gleft => Gsignal_1_31_port, gright => 
                           Gsignal_1_30_port, pleft => Psignal_1_31_port, 
                           pright => Psignal_1_30_port, pout => 
                           Psignal_2_31_port, gout => Gsignal_2_31_port);
   Gblock_2_3 : G port map( gleft => Gsignal_2_3_port, gright => 
                           Gsignal_2_1_port, pleft => Psignal_2_3_port, gout =>
                           Cout_1_port);
   PGblock_2_7 : PG port map( gleft => Gsignal_2_7_port, gright => 
                           Gsignal_2_5_port, pleft => Psignal_2_7_port, pright 
                           => Psignal_2_5_port, pout => Psignal_3_7_port, gout 
                           => Gsignal_3_7_port);
   PGblock_2_11 : PG port map( gleft => Gsignal_2_11_port, gright => 
                           Gsignal_2_9_port, pleft => Psignal_2_11_port, pright
                           => Psignal_2_9_port, pout => Psignal_3_11_port, gout
                           => Gsignal_3_11_port);
   PGblock_2_15 : PG port map( gleft => Gsignal_2_15_port, gright => 
                           Gsignal_2_13_port, pleft => Psignal_2_15_port, 
                           pright => Psignal_2_13_port, pout => 
                           Psignal_3_15_port, gout => Gsignal_3_15_port);
   PGblock_2_19 : PG port map( gleft => Gsignal_2_19_port, gright => 
                           Gsignal_2_17_port, pleft => Psignal_2_19_port, 
                           pright => Psignal_2_17_port, pout => 
                           Psignal_3_19_port, gout => Gsignal_3_19_port);
   PGblock_2_23 : PG port map( gleft => Gsignal_2_23_port, gright => 
                           Gsignal_2_21_port, pleft => Psignal_2_23_port, 
                           pright => Psignal_2_21_port, pout => 
                           Psignal_3_23_port, gout => Gsignal_3_23_port);
   PGblock_2_27 : PG port map( gleft => Gsignal_2_27_port, gright => 
                           Gsignal_2_25_port, pleft => Psignal_2_27_port, 
                           pright => Psignal_2_25_port, pout => 
                           Psignal_3_27_port, gout => Gsignal_3_27_port);
   PGblock_2_31 : PG port map( gleft => Gsignal_2_31_port, gright => 
                           Gsignal_2_29_port, pleft => Psignal_2_31_port, 
                           pright => Psignal_2_29_port, pout => 
                           Psignal_3_31_port, gout => Gsignal_3_31_port);
   Gblock_3_7 : G port map( gleft => Gsignal_3_7_port, gright => Cout_1_port, 
                           pleft => Psignal_3_7_port, gout => Cout_2_port);
   PGblock_3_15 : PG port map( gleft => Gsignal_3_15_port, gright => 
                           Gsignal_3_11_port, pleft => Psignal_3_15_port, 
                           pright => Psignal_3_11_port, pout => 
                           Psignal_4_15_port, gout => Gsignal_4_15_port);
   PGblock_3_23 : PG port map( gleft => Gsignal_3_23_port, gright => 
                           Gsignal_3_19_port, pleft => Psignal_3_23_port, 
                           pright => Psignal_3_19_port, pout => 
                           Psignal_4_23_port, gout => Gsignal_4_23_port);
   PGblock_3_31 : PG port map( gleft => Gsignal_3_31_port, gright => 
                           Gsignal_3_27_port, pleft => Psignal_3_31_port, 
                           pright => Psignal_3_27_port, pout => 
                           Psignal_4_31_port, gout => Gsignal_4_31_port);
   Gblock_4_11 : G port map( gleft => Gsignal_3_11_port, gright => Cout_2_port,
                           pleft => Psignal_3_11_port, gout => Cout_3_port);
   Gblock_4_15 : G port map( gleft => Gsignal_4_15_port, gright => Cout_2_port,
                           pleft => Psignal_4_15_port, gout => Cout_4_port);
   PGblock_4_27 : PG port map( gleft => Gsignal_3_27_port, gright => 
                           Gsignal_4_23_port, pleft => Psignal_3_27_port, 
                           pright => Psignal_4_23_port, pout => 
                           Psignal_5_27_port, gout => Gsignal_5_27_port);
   PGblock_4_31 : PG port map( gleft => Gsignal_4_31_port, gright => 
                           Gsignal_4_23_port, pleft => Psignal_4_31_port, 
                           pright => Psignal_4_23_port, pout => 
                           Psignal_5_31_port, gout => Gsignal_5_31_port);
   Gblock_5_19 : G port map( gleft => Gsignal_3_19_port, gright => Cout_4_port,
                           pleft => Psignal_3_19_port, gout => Cout_5_port);
   Gblock_5_23 : G port map( gleft => Gsignal_4_23_port, gright => Cout_4_port,
                           pleft => Psignal_4_23_port, gout => Cout_6_port);
   Gblock_5_27 : G port map( gleft => Gsignal_5_27_port, gright => Cout_4_port,
                           pleft => Psignal_5_27_port, gout => Cout_7_port);
   Gblock_5_31 : G port map( gleft => Gsignal_5_31_port, gright => Cout_4_port,
                           pleft => Psignal_5_31_port, gout => Cout_8_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_alu is

   port( addsub, mul, log, shift, lhi : in std_logic_vector (31 downto 0);  gt,
         get, lt, let, eq, neq : in std_logic;  sel : in std_logic_vector (0 to
         4);  out_mux : out std_logic_vector (31 downto 0));

end mux_alu;

architecture SYN_behav of mux_alu is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n2, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n144 : std_logic;

begin
   
   U128 : OAI33_X1 port map( A1 => n101, A2 => n30, A3 => n102, B1 => n103, B2 
                           => sel(0), B3 => sel(2), ZN => n16);
   out_mux_tri_0_inst : TBUF_X1 port map( A => n153, EN => n119, Z => 
                           out_mux(0));
   out_mux_tri_1_inst : TBUF_X1 port map( A => n152, EN => n119, Z => 
                           out_mux(1));
   out_mux_tri_2_inst : TBUF_X1 port map( A => n151, EN => n119, Z => 
                           out_mux(2));
   out_mux_tri_3_inst : TBUF_X1 port map( A => n150, EN => n119, Z => 
                           out_mux(3));
   out_mux_tri_4_inst : TBUF_X1 port map( A => n149, EN => n119, Z => 
                           out_mux(4));
   out_mux_tri_5_inst : TBUF_X1 port map( A => n148, EN => n119, Z => 
                           out_mux(5));
   out_mux_tri_6_inst : TBUF_X1 port map( A => n147, EN => n119, Z => 
                           out_mux(6));
   out_mux_tri_7_inst : TBUF_X1 port map( A => n146, EN => n119, Z => 
                           out_mux(7));
   out_mux_tri_8_inst : TBUF_X1 port map( A => n145, EN => n119, Z => 
                           out_mux(8));
   out_mux_tri_9_inst : TBUF_X1 port map( A => n143, EN => n119, Z => 
                           out_mux(9));
   out_mux_tri_10_inst : TBUF_X1 port map( A => n142, EN => n119, Z => 
                           out_mux(10));
   out_mux_tri_11_inst : TBUF_X1 port map( A => n141, EN => n119, Z => 
                           out_mux(11));
   out_mux_tri_12_inst : TBUF_X1 port map( A => n140, EN => n120, Z => 
                           out_mux(12));
   out_mux_tri_13_inst : TBUF_X1 port map( A => n139, EN => n120, Z => 
                           out_mux(13));
   out_mux_tri_14_inst : TBUF_X1 port map( A => n138, EN => n120, Z => 
                           out_mux(14));
   out_mux_tri_15_inst : TBUF_X1 port map( A => n137, EN => n120, Z => 
                           out_mux(15));
   out_mux_tri_16_inst : TBUF_X1 port map( A => n136, EN => n120, Z => 
                           out_mux(16));
   out_mux_tri_17_inst : TBUF_X1 port map( A => n135, EN => n120, Z => 
                           out_mux(17));
   out_mux_tri_18_inst : TBUF_X1 port map( A => n134, EN => n120, Z => 
                           out_mux(18));
   out_mux_tri_19_inst : TBUF_X1 port map( A => n133, EN => n120, Z => 
                           out_mux(19));
   out_mux_tri_20_inst : TBUF_X1 port map( A => n132, EN => n120, Z => 
                           out_mux(20));
   out_mux_tri_21_inst : TBUF_X1 port map( A => n131, EN => n120, Z => 
                           out_mux(21));
   out_mux_tri_22_inst : TBUF_X1 port map( A => n130, EN => n120, Z => 
                           out_mux(22));
   out_mux_tri_23_inst : TBUF_X1 port map( A => n129, EN => n120, Z => 
                           out_mux(23));
   out_mux_tri_24_inst : TBUF_X1 port map( A => n128, EN => n144, Z => 
                           out_mux(24));
   out_mux_tri_25_inst : TBUF_X1 port map( A => n127, EN => n144, Z => 
                           out_mux(25));
   out_mux_tri_26_inst : TBUF_X1 port map( A => n126, EN => n144, Z => 
                           out_mux(26));
   out_mux_tri_27_inst : TBUF_X1 port map( A => n125, EN => n144, Z => 
                           out_mux(27));
   out_mux_tri_28_inst : TBUF_X1 port map( A => n124, EN => n144, Z => 
                           out_mux(28));
   out_mux_tri_29_inst : TBUF_X1 port map( A => n123, EN => n144, Z => 
                           out_mux(29));
   out_mux_tri_30_inst : TBUF_X1 port map( A => n122, EN => n144, Z => 
                           out_mux(30));
   out_mux_tri_31_inst : TBUF_X1 port map( A => n121, EN => n144, Z => 
                           out_mux(31));
   U2 : BUF_X1 port map( A => n38, Z => n104);
   U3 : BUF_X1 port map( A => n38, Z => n105);
   U4 : BUF_X1 port map( A => n38, Z => n106);
   U5 : NOR3_X1 port map( A1 => n30, A2 => n25, A3 => n101, ZN => n38);
   U6 : BUF_X1 port map( A => n17, Z => n113);
   U7 : BUF_X1 port map( A => n17, Z => n114);
   U8 : BUF_X1 port map( A => n37, Z => n107);
   U9 : BUF_X1 port map( A => n37, Z => n108);
   U10 : BUF_X1 port map( A => n16, Z => n116);
   U11 : BUF_X1 port map( A => n16, Z => n117);
   U12 : BUF_X1 port map( A => n36, Z => n110);
   U13 : BUF_X1 port map( A => n36, Z => n111);
   U14 : BUF_X1 port map( A => n16, Z => n118);
   U15 : BUF_X1 port map( A => n36, Z => n112);
   U16 : AOI22_X1 port map( A1 => n24, A2 => gt, B1 => n25, B2 => let, ZN => 
                           n23);
   U17 : BUF_X1 port map( A => n2, Z => n120);
   U18 : BUF_X1 port map( A => n2, Z => n119);
   U19 : INV_X1 port map( A => n102, ZN => n25);
   U20 : BUF_X1 port map( A => n2, Z => n144);
   U21 : BUF_X1 port map( A => n17, Z => n115);
   U22 : NAND2_X1 port map( A1 => n10, A2 => n12, ZN => n101);
   U23 : BUF_X1 port map( A => n37, Z => n109);
   U24 : INV_X1 port map( A => n24, ZN => n13);
   U25 : INV_X1 port map( A => n35, ZN => n29);
   U26 : AOI22_X1 port map( A1 => get, A2 => n25, B1 => n26, B2 => gt, ZN => 
                           n35);
   U27 : NAND2_X1 port map( A1 => sel(1), A2 => n28, ZN => n103);
   U28 : NOR4_X1 port map( A1 => n13, A2 => n12, A3 => n30, A4 => sel(1), ZN =>
                           n17);
   U29 : NOR4_X1 port map( A1 => n101, A2 => n25, A3 => n24, A4 => sel(2), ZN 
                           => n36);
   U30 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n127);
   U31 : AOI22_X1 port map( A1 => log(25), A2 => n104, B1 => addsub(25), B2 => 
                           n110, ZN => n87);
   U32 : AOI222_X1 port map( A1 => mul(25), A2 => n108, B1 => shift(25), B2 => 
                           n116, C1 => lhi(25), C2 => n114, ZN => n88);
   U33 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => n128);
   U34 : AOI22_X1 port map( A1 => log(24), A2 => n104, B1 => addsub(24), B2 => 
                           n110, ZN => n85);
   U35 : AOI222_X1 port map( A1 => mul(24), A2 => n108, B1 => shift(24), B2 => 
                           n116, C1 => lhi(24), C2 => n114, ZN => n86);
   U36 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => n129);
   U37 : AOI22_X1 port map( A1 => log(23), A2 => n104, B1 => addsub(23), B2 => 
                           n110, ZN => n83);
   U38 : AOI222_X1 port map( A1 => mul(23), A2 => n108, B1 => shift(23), B2 => 
                           n116, C1 => lhi(23), C2 => n114, ZN => n84);
   U39 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n130);
   U40 : AOI22_X1 port map( A1 => log(22), A2 => n104, B1 => addsub(22), B2 => 
                           n110, ZN => n81);
   U41 : AOI222_X1 port map( A1 => mul(22), A2 => n108, B1 => shift(22), B2 => 
                           n116, C1 => lhi(22), C2 => n114, ZN => n82);
   U42 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n131);
   U43 : AOI22_X1 port map( A1 => log(21), A2 => n104, B1 => addsub(21), B2 => 
                           n110, ZN => n79);
   U44 : AOI222_X1 port map( A1 => mul(21), A2 => n108, B1 => shift(21), B2 => 
                           n116, C1 => lhi(21), C2 => n114, ZN => n80);
   U45 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n132);
   U46 : AOI22_X1 port map( A1 => log(20), A2 => n104, B1 => addsub(20), B2 => 
                           n110, ZN => n77);
   U47 : AOI222_X1 port map( A1 => mul(20), A2 => n108, B1 => shift(20), B2 => 
                           n116, C1 => lhi(20), C2 => n114, ZN => n78);
   U48 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => n133);
   U49 : AOI22_X1 port map( A1 => log(19), A2 => n105, B1 => addsub(19), B2 => 
                           n111, ZN => n75);
   U50 : AOI222_X1 port map( A1 => mul(19), A2 => n108, B1 => shift(19), B2 => 
                           n117, C1 => lhi(19), C2 => n114, ZN => n76);
   U51 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => n134);
   U52 : AOI22_X1 port map( A1 => log(18), A2 => n105, B1 => addsub(18), B2 => 
                           n111, ZN => n73);
   U53 : AOI222_X1 port map( A1 => mul(18), A2 => n108, B1 => shift(18), B2 => 
                           n117, C1 => lhi(18), C2 => n114, ZN => n74);
   U54 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n135);
   U55 : AOI22_X1 port map( A1 => log(17), A2 => n105, B1 => addsub(17), B2 => 
                           n111, ZN => n71);
   U56 : AOI222_X1 port map( A1 => mul(17), A2 => n108, B1 => shift(17), B2 => 
                           n117, C1 => lhi(17), C2 => n114, ZN => n72);
   U57 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => n136);
   U58 : AOI22_X1 port map( A1 => log(16), A2 => n105, B1 => addsub(16), B2 => 
                           n111, ZN => n69);
   U59 : AOI222_X1 port map( A1 => mul(16), A2 => n108, B1 => shift(16), B2 => 
                           n117, C1 => lhi(16), C2 => n114, ZN => n70);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => n137);
   U61 : AOI22_X1 port map( A1 => log(15), A2 => n105, B1 => addsub(15), B2 => 
                           n111, ZN => n67);
   U62 : AOI222_X1 port map( A1 => mul(15), A2 => n108, B1 => shift(15), B2 => 
                           n117, C1 => lhi(15), C2 => n114, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => n138);
   U64 : AOI22_X1 port map( A1 => log(14), A2 => n105, B1 => addsub(14), B2 => 
                           n111, ZN => n65);
   U65 : AOI222_X1 port map( A1 => mul(14), A2 => n108, B1 => shift(14), B2 => 
                           n117, C1 => lhi(14), C2 => n114, ZN => n66);
   U66 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n139);
   U67 : AOI22_X1 port map( A1 => log(13), A2 => n105, B1 => addsub(13), B2 => 
                           n111, ZN => n63);
   U68 : AOI222_X1 port map( A1 => mul(13), A2 => n108, B1 => shift(13), B2 => 
                           n117, C1 => lhi(13), C2 => n114, ZN => n64);
   U69 : NOR3_X1 port map( A1 => n102, A2 => sel(2), A3 => n101, ZN => n37);
   U70 : NOR2_X1 port map( A1 => sel(3), A2 => sel(4), ZN => n24);
   U71 : AOI21_X1 port map( B1 => n10, B2 => n11, A => n12, ZN => n2);
   U72 : NAND2_X1 port map( A1 => sel(2), A2 => n13, ZN => n11);
   U73 : NOR2_X1 port map( A1 => n28, A2 => sel(4), ZN => n26);
   U74 : INV_X1 port map( A => sel(2), ZN => n30);
   U75 : AOI21_X1 port map( B1 => n26, B2 => lt, A => n27, ZN => n22);
   U76 : AND3_X1 port map( A1 => get, A2 => n28, A3 => sel(4), ZN => n27);
   U77 : AOI21_X1 port map( B1 => n32, B2 => n33, A => n30, ZN => n31);
   U78 : AOI21_X1 port map( B1 => eq, B2 => n26, A => n34, ZN => n33);
   U79 : AOI22_X1 port map( A1 => neq, A2 => n25, B1 => n24, B2 => lt, ZN => 
                           n32);
   U80 : AND3_X1 port map( A1 => let, A2 => n28, A3 => sel(4), ZN => n34);
   U81 : INV_X1 port map( A => sel(0), ZN => n12);
   U82 : OAI21_X1 port map( B1 => n19, B2 => n10, A => n20, ZN => n18);
   U83 : INV_X1 port map( A => n21, ZN => n20);
   U84 : AOI21_X1 port map( B1 => n29, B2 => n30, A => n31, ZN => n19);
   U85 : AOI211_X1 port map( C1 => n22, C2 => n23, A => sel(2), B => n12, ZN =>
                           n21);
   U86 : NAND2_X1 port map( A1 => sel(3), A2 => sel(4), ZN => n102);
   U87 : INV_X1 port map( A => sel(3), ZN => n28);
   U88 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n153);
   U89 : AOI222_X1 port map( A1 => addsub(0), A2 => n112, B1 => mul(0), B2 => 
                           n107, C1 => log(0), C2 => n106, ZN => n14);
   U90 : AOI221_X1 port map( B1 => shift(0), B2 => n118, C1 => lhi(0), C2 => 
                           n113, A => n18, ZN => n15);
   U91 : INV_X1 port map( A => sel(1), ZN => n10);
   U92 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => n146);
   U93 : AOI22_X1 port map( A1 => log(7), A2 => n106, B1 => addsub(7), B2 => 
                           n112, ZN => n51);
   U94 : AOI222_X1 port map( A1 => mul(7), A2 => n107, B1 => shift(7), B2 => 
                           n118, C1 => lhi(7), C2 => n113, ZN => n52);
   U95 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n147);
   U96 : AOI22_X1 port map( A1 => log(6), A2 => n106, B1 => addsub(6), B2 => 
                           n112, ZN => n49);
   U97 : AOI222_X1 port map( A1 => mul(6), A2 => n107, B1 => shift(6), B2 => 
                           n118, C1 => lhi(6), C2 => n113, ZN => n50);
   U98 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => n148);
   U99 : AOI22_X1 port map( A1 => log(5), A2 => n106, B1 => addsub(5), B2 => 
                           n112, ZN => n47);
   U100 : AOI222_X1 port map( A1 => mul(5), A2 => n107, B1 => shift(5), B2 => 
                           n118, C1 => lhi(5), C2 => n113, ZN => n48);
   U101 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n149);
   U102 : AOI22_X1 port map( A1 => log(4), A2 => n106, B1 => addsub(4), B2 => 
                           n112, ZN => n45);
   U103 : AOI222_X1 port map( A1 => mul(4), A2 => n107, B1 => shift(4), B2 => 
                           n118, C1 => lhi(4), C2 => n113, ZN => n46);
   U104 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n150);
   U105 : AOI22_X1 port map( A1 => log(3), A2 => n106, B1 => addsub(3), B2 => 
                           n112, ZN => n43);
   U106 : AOI222_X1 port map( A1 => mul(3), A2 => n107, B1 => shift(3), B2 => 
                           n118, C1 => lhi(3), C2 => n113, ZN => n44);
   U107 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n151);
   U108 : AOI22_X1 port map( A1 => log(2), A2 => n106, B1 => addsub(2), B2 => 
                           n112, ZN => n41);
   U109 : AOI222_X1 port map( A1 => mul(2), A2 => n107, B1 => shift(2), B2 => 
                           n118, C1 => lhi(2), C2 => n113, ZN => n42);
   U110 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n152);
   U111 : AOI22_X1 port map( A1 => log(1), A2 => n106, B1 => addsub(1), B2 => 
                           n112, ZN => n39);
   U112 : AOI222_X1 port map( A1 => mul(1), A2 => n107, B1 => shift(1), B2 => 
                           n118, C1 => lhi(1), C2 => n113, ZN => n40);
   U113 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n121);
   U114 : AOI22_X1 port map( A1 => log(31), A2 => n104, B1 => addsub(31), B2 =>
                           n110, ZN => n99);
   U115 : AOI222_X1 port map( A1 => mul(31), A2 => n109, B1 => shift(31), B2 =>
                           n116, C1 => lhi(31), C2 => n115, ZN => n100);
   U116 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n122);
   U117 : AOI22_X1 port map( A1 => log(30), A2 => n104, B1 => addsub(30), B2 =>
                           n110, ZN => n97);
   U118 : AOI222_X1 port map( A1 => mul(30), A2 => n109, B1 => shift(30), B2 =>
                           n116, C1 => lhi(30), C2 => n115, ZN => n98);
   U119 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n123);
   U120 : AOI22_X1 port map( A1 => log(29), A2 => n104, B1 => addsub(29), B2 =>
                           n110, ZN => n95);
   U121 : AOI222_X1 port map( A1 => mul(29), A2 => n109, B1 => shift(29), B2 =>
                           n116, C1 => lhi(29), C2 => n115, ZN => n96);
   U122 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => n124);
   U123 : AOI22_X1 port map( A1 => log(28), A2 => n104, B1 => addsub(28), B2 =>
                           n110, ZN => n93);
   U124 : AOI222_X1 port map( A1 => mul(28), A2 => n109, B1 => shift(28), B2 =>
                           n116, C1 => lhi(28), C2 => n115, ZN => n94);
   U125 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => n125);
   U126 : AOI22_X1 port map( A1 => log(27), A2 => n104, B1 => addsub(27), B2 =>
                           n110, ZN => n91);
   U127 : AOI222_X1 port map( A1 => mul(27), A2 => n109, B1 => shift(27), B2 =>
                           n116, C1 => lhi(27), C2 => n115, ZN => n92);
   U129 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n126);
   U130 : AOI22_X1 port map( A1 => log(26), A2 => n104, B1 => addsub(26), B2 =>
                           n110, ZN => n89);
   U131 : AOI222_X1 port map( A1 => mul(26), A2 => n109, B1 => shift(26), B2 =>
                           n116, C1 => lhi(26), C2 => n115, ZN => n90);
   U132 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n140);
   U133 : AOI22_X1 port map( A1 => log(12), A2 => n105, B1 => addsub(12), B2 =>
                           n111, ZN => n61);
   U134 : AOI222_X1 port map( A1 => mul(12), A2 => n107, B1 => shift(12), B2 =>
                           n117, C1 => lhi(12), C2 => n113, ZN => n62);
   U135 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => n141);
   U136 : AOI22_X1 port map( A1 => log(11), A2 => n105, B1 => addsub(11), B2 =>
                           n111, ZN => n59);
   U137 : AOI222_X1 port map( A1 => mul(11), A2 => n107, B1 => shift(11), B2 =>
                           n117, C1 => lhi(11), C2 => n113, ZN => n60);
   U138 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n142);
   U139 : AOI22_X1 port map( A1 => log(10), A2 => n105, B1 => addsub(10), B2 =>
                           n111, ZN => n57);
   U140 : AOI222_X1 port map( A1 => mul(10), A2 => n107, B1 => shift(10), B2 =>
                           n117, C1 => lhi(10), C2 => n113, ZN => n58);
   U141 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n143);
   U142 : AOI22_X1 port map( A1 => log(9), A2 => n105, B1 => addsub(9), B2 => 
                           n111, ZN => n55);
   U143 : AOI222_X1 port map( A1 => mul(9), A2 => n107, B1 => shift(9), B2 => 
                           n117, C1 => lhi(9), C2 => n113, ZN => n56);
   U144 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n145);
   U145 : AOI22_X1 port map( A1 => log(8), A2 => n105, B1 => addsub(8), B2 => 
                           n111, ZN => n53);
   U146 : AOI222_X1 port map( A1 => mul(8), A2 => n107, B1 => shift(8), B2 => 
                           n117, C1 => lhi(8), C2 => n113, ZN => n54);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity comparator is

   port( C : in std_logic;  Sum : in std_logic_vector (31 downto 0);  sign : in
         std_logic;  gt, get, lt, let, eq, neq : out std_logic);

end comparator;

architecture SYN_behav of comparator is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal gt_port, get_port, lt_port, eq_port, n4, n5, n6, n7, n8, n9, n10, n11
      , n12, n13 : std_logic;

begin
   gt <= gt_port;
   get <= get_port;
   lt <= lt_port;
   eq <= eq_port;
   
   U16 : XOR2_X1 port map( A => sign, B => C, Z => get_port);
   U1 : INV_X1 port map( A => gt_port, ZN => let);
   U2 : INV_X1 port map( A => eq_port, ZN => neq);
   U3 : NOR4_X1 port map( A1 => Sum(23), A2 => Sum(22), A3 => Sum(21), A4 => 
                           Sum(20), ZN => n9);
   U4 : NOR4_X1 port map( A1 => Sum(9), A2 => Sum(8), A3 => Sum(7), A4 => 
                           Sum(6), ZN => n13);
   U5 : NOR4_X1 port map( A1 => Sum(16), A2 => Sum(15), A3 => Sum(14), A4 => 
                           Sum(13), ZN => n7);
   U6 : NOR2_X1 port map( A1 => lt_port, A2 => eq_port, ZN => gt_port);
   U7 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => eq_port);
   U8 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => n4
                           );
   U9 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U10 : NOR4_X1 port map( A1 => Sum(27), A2 => Sum(26), A3 => Sum(25), A4 => 
                           Sum(24), ZN => n10);
   U11 : NOR4_X1 port map( A1 => Sum(1), A2 => Sum(19), A3 => Sum(18), A4 => 
                           Sum(17), ZN => n8);
   U12 : NOR4_X1 port map( A1 => Sum(5), A2 => Sum(4), A3 => Sum(3), A4 => 
                           Sum(31), ZN => n12);
   U13 : NOR4_X1 port map( A1 => Sum(30), A2 => Sum(2), A3 => Sum(29), A4 => 
                           Sum(28), ZN => n11);
   U14 : NOR4_X1 port map( A1 => Sum(12), A2 => Sum(11), A3 => Sum(10), A4 => 
                           Sum(0), ZN => n6);
   U15 : INV_X1 port map( A => get_port, ZN => lt_port);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity shifter is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (1 downto 0);  C : out std_logic_vector (31 downto 0));

end shifter;

architecture SYN_struct of shifter is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_thirdLevel
      port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector 
            (38 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_secondLevel
      port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : 
            in std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 
            downto 0));
   end component;
   
   component shift_firstLevel
      port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
            (1 downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 
            downto 0));
   end component;
   
   signal s3_2_port, s3_1_port, s3_0_port, m0_38_port, m0_37_port, m0_36_port, 
      m0_35_port, m0_34_port, m0_33_port, m0_32_port, m0_31_port, m0_30_port, 
      m0_29_port, m0_28_port, m0_27_port, m0_26_port, m0_25_port, m0_24_port, 
      m0_23_port, m0_22_port, m0_21_port, m0_20_port, m0_19_port, m0_18_port, 
      m0_17_port, m0_16_port, m0_15_port, m0_14_port, m0_13_port, m0_12_port, 
      m0_11_port, m0_10_port, m0_9_port, m0_8_port, m0_7_port, m0_6_port, 
      m0_5_port, m0_4_port, m0_3_port, m0_2_port, m0_1_port, m0_0_port, 
      m8_38_port, m8_37_port, m8_36_port, m8_35_port, m8_34_port, m8_33_port, 
      m8_32_port, m8_31_port, m8_30_port, m8_29_port, m8_28_port, m8_27_port, 
      m8_26_port, m8_25_port, m8_24_port, m8_23_port, m8_22_port, m8_21_port, 
      m8_20_port, m8_19_port, m8_18_port, m8_17_port, m8_16_port, m8_15_port, 
      m8_14_port, m8_13_port, m8_12_port, m8_11_port, m8_10_port, m8_9_port, 
      m8_8_port, m8_7_port, m8_6_port, m8_5_port, m8_4_port, m8_3_port, 
      m8_2_port, m8_1_port, m8_0_port, m16_38_port, m16_37_port, m16_36_port, 
      m16_35_port, m16_34_port, m16_33_port, m16_32_port, m16_31_port, 
      m16_30_port, m16_29_port, m16_28_port, m16_27_port, m16_26_port, 
      m16_25_port, m16_24_port, m16_23_port, m16_22_port, m16_21_port, 
      m16_20_port, m16_19_port, m16_18_port, m16_17_port, m16_16_port, 
      m16_15_port, m16_14_port, m16_13_port, m16_12_port, m16_11_port, 
      m16_10_port, m16_9_port, m16_8_port, m16_7_port, m16_6_port, m16_5_port, 
      m16_4_port, m16_3_port, m16_2_port, m16_1_port, m16_0_port, y_38_port, 
      y_37_port, y_36_port, y_35_port, y_34_port, y_33_port, y_32_port, 
      y_31_port, y_30_port, y_29_port, y_28_port, y_27_port, y_26_port, 
      y_25_port, y_24_port, y_23_port, y_22_port, y_21_port, y_20_port, 
      y_19_port, y_18_port, y_17_port, y_16_port, y_15_port, y_14_port, 
      y_13_port, y_12_port, y_11_port, y_10_port, y_9_port, y_8_port, y_7_port,
      y_6_port, y_5_port, y_4_port, y_3_port, y_2_port, y_1_port, y_0_port, n6,
      n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   IL : shift_firstLevel port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), sel(1) => sel(1), sel(0) => sel(0), 
                           mask00(38) => m0_38_port, mask00(37) => m0_37_port, 
                           mask00(36) => m0_36_port, mask00(35) => m0_35_port, 
                           mask00(34) => m0_34_port, mask00(33) => m0_33_port, 
                           mask00(32) => m0_32_port, mask00(31) => m0_31_port, 
                           mask00(30) => m0_30_port, mask00(29) => m0_29_port, 
                           mask00(28) => m0_28_port, mask00(27) => m0_27_port, 
                           mask00(26) => m0_26_port, mask00(25) => m0_25_port, 
                           mask00(24) => m0_24_port, mask00(23) => m0_23_port, 
                           mask00(22) => m0_22_port, mask00(21) => m0_21_port, 
                           mask00(20) => m0_20_port, mask00(19) => m0_19_port, 
                           mask00(18) => m0_18_port, mask00(17) => m0_17_port, 
                           mask00(16) => m0_16_port, mask00(15) => m0_15_port, 
                           mask00(14) => m0_14_port, mask00(13) => m0_13_port, 
                           mask00(12) => m0_12_port, mask00(11) => m0_11_port, 
                           mask00(10) => m0_10_port, mask00(9) => m0_9_port, 
                           mask00(8) => m0_8_port, mask00(7) => m0_7_port, 
                           mask00(6) => m0_6_port, mask00(5) => m0_5_port, 
                           mask00(4) => m0_4_port, mask00(3) => m0_3_port, 
                           mask00(2) => m0_2_port, mask00(1) => m0_1_port, 
                           mask00(0) => m0_0_port, mask08(38) => m8_38_port, 
                           mask08(37) => m8_37_port, mask08(36) => m8_36_port, 
                           mask08(35) => m8_35_port, mask08(34) => m8_34_port, 
                           mask08(33) => m8_33_port, mask08(32) => m8_32_port, 
                           mask08(31) => m8_31_port, mask08(30) => m8_30_port, 
                           mask08(29) => m8_29_port, mask08(28) => m8_28_port, 
                           mask08(27) => m8_27_port, mask08(26) => m8_26_port, 
                           mask08(25) => m8_25_port, mask08(24) => m8_24_port, 
                           mask08(23) => m8_23_port, mask08(22) => m8_22_port, 
                           mask08(21) => m8_21_port, mask08(20) => m8_20_port, 
                           mask08(19) => m8_19_port, mask08(18) => m8_18_port, 
                           mask08(17) => m8_17_port, mask08(16) => m8_16_port, 
                           mask08(15) => m8_15_port, mask08(14) => m8_14_port, 
                           mask08(13) => m8_13_port, mask08(12) => m8_12_port, 
                           mask08(11) => m8_11_port, mask08(10) => m8_10_port, 
                           mask08(9) => m8_9_port, mask08(8) => m8_8_port, 
                           mask08(7) => m8_7_port, mask08(6) => m8_6_port, 
                           mask08(5) => m8_5_port, mask08(4) => m8_4_port, 
                           mask08(3) => m8_3_port, mask08(2) => m8_2_port, 
                           mask08(1) => m8_1_port, mask08(0) => m8_0_port, 
                           mask16(38) => m16_38_port, mask16(37) => m16_37_port
                           , mask16(36) => m16_36_port, mask16(35) => 
                           m16_35_port, mask16(34) => m16_34_port, mask16(33) 
                           => m16_33_port, mask16(32) => m16_32_port, 
                           mask16(31) => m16_31_port, mask16(30) => m16_30_port
                           , mask16(29) => m16_29_port, mask16(28) => 
                           m16_28_port, mask16(27) => m16_27_port, mask16(26) 
                           => m16_26_port, mask16(25) => m16_25_port, 
                           mask16(24) => m16_24_port, mask16(23) => m16_23_port
                           , mask16(22) => m16_22_port, mask16(21) => 
                           m16_21_port, mask16(20) => m16_20_port, mask16(19) 
                           => m16_19_port, mask16(18) => m16_18_port, 
                           mask16(17) => m16_17_port, mask16(16) => m16_16_port
                           , mask16(15) => m16_15_port, mask16(14) => 
                           m16_14_port, mask16(13) => m16_13_port, mask16(12) 
                           => m16_12_port, mask16(11) => m16_11_port, 
                           mask16(10) => m16_10_port, mask16(9) => m16_9_port, 
                           mask16(8) => m16_8_port, mask16(7) => m16_7_port, 
                           mask16(6) => m16_6_port, mask16(5) => m16_5_port, 
                           mask16(4) => m16_4_port, mask16(3) => m16_3_port, 
                           mask16(2) => m16_2_port, mask16(1) => m16_1_port, 
                           mask16(0) => m16_0_port);
   IIL : shift_secondLevel port map( sel(1) => B(4), sel(0) => B(3), mask00(38)
                           => m0_38_port, mask00(37) => m0_37_port, mask00(36) 
                           => m0_36_port, mask00(35) => m0_35_port, mask00(34) 
                           => m0_34_port, mask00(33) => m0_33_port, mask00(32) 
                           => m0_32_port, mask00(31) => m0_31_port, mask00(30) 
                           => m0_30_port, mask00(29) => m0_29_port, mask00(28) 
                           => m0_28_port, mask00(27) => m0_27_port, mask00(26) 
                           => m0_26_port, mask00(25) => m0_25_port, mask00(24) 
                           => m0_24_port, mask00(23) => m0_23_port, mask00(22) 
                           => m0_22_port, mask00(21) => m0_21_port, mask00(20) 
                           => m0_20_port, mask00(19) => m0_19_port, mask00(18) 
                           => m0_18_port, mask00(17) => m0_17_port, mask00(16) 
                           => m0_16_port, mask00(15) => m0_15_port, mask00(14) 
                           => m0_14_port, mask00(13) => m0_13_port, mask00(12) 
                           => m0_12_port, mask00(11) => m0_11_port, mask00(10) 
                           => m0_10_port, mask00(9) => m0_9_port, mask00(8) => 
                           m0_8_port, mask00(7) => m0_7_port, mask00(6) => 
                           m0_6_port, mask00(5) => m0_5_port, mask00(4) => 
                           m0_4_port, mask00(3) => m0_3_port, mask00(2) => 
                           m0_2_port, mask00(1) => m0_1_port, mask00(0) => 
                           m0_0_port, mask08(38) => m8_38_port, mask08(37) => 
                           m8_37_port, mask08(36) => m8_36_port, mask08(35) => 
                           m8_35_port, mask08(34) => m8_34_port, mask08(33) => 
                           m8_33_port, mask08(32) => m8_32_port, mask08(31) => 
                           m8_31_port, mask08(30) => m8_30_port, mask08(29) => 
                           m8_29_port, mask08(28) => m8_28_port, mask08(27) => 
                           m8_27_port, mask08(26) => m8_26_port, mask08(25) => 
                           m8_25_port, mask08(24) => m8_24_port, mask08(23) => 
                           m8_23_port, mask08(22) => m8_22_port, mask08(21) => 
                           m8_21_port, mask08(20) => m8_20_port, mask08(19) => 
                           m8_19_port, mask08(18) => m8_18_port, mask08(17) => 
                           m8_17_port, mask08(16) => m8_16_port, mask08(15) => 
                           m8_15_port, mask08(14) => m8_14_port, mask08(13) => 
                           m8_13_port, mask08(12) => m8_12_port, mask08(11) => 
                           m8_11_port, mask08(10) => m8_10_port, mask08(9) => 
                           m8_9_port, mask08(8) => m8_8_port, mask08(7) => 
                           m8_7_port, mask08(6) => m8_6_port, mask08(5) => 
                           m8_5_port, mask08(4) => m8_4_port, mask08(3) => 
                           m8_3_port, mask08(2) => m8_2_port, mask08(1) => 
                           m8_1_port, mask08(0) => m8_0_port, mask16(38) => 
                           m16_38_port, mask16(37) => m16_37_port, mask16(36) 
                           => m16_36_port, mask16(35) => m16_35_port, 
                           mask16(34) => m16_34_port, mask16(33) => m16_33_port
                           , mask16(32) => m16_32_port, mask16(31) => 
                           m16_31_port, mask16(30) => m16_30_port, mask16(29) 
                           => m16_29_port, mask16(28) => m16_28_port, 
                           mask16(27) => m16_27_port, mask16(26) => m16_26_port
                           , mask16(25) => m16_25_port, mask16(24) => 
                           m16_24_port, mask16(23) => m16_23_port, mask16(22) 
                           => m16_22_port, mask16(21) => m16_21_port, 
                           mask16(20) => m16_20_port, mask16(19) => m16_19_port
                           , mask16(18) => m16_18_port, mask16(17) => 
                           m16_17_port, mask16(16) => m16_16_port, mask16(15) 
                           => m16_15_port, mask16(14) => m16_14_port, 
                           mask16(13) => m16_13_port, mask16(12) => m16_12_port
                           , mask16(11) => m16_11_port, mask16(10) => 
                           m16_10_port, mask16(9) => m16_9_port, mask16(8) => 
                           m16_8_port, mask16(7) => m16_7_port, mask16(6) => 
                           m16_6_port, mask16(5) => m16_5_port, mask16(4) => 
                           m16_4_port, mask16(3) => m16_3_port, mask16(2) => 
                           m16_2_port, mask16(1) => m16_1_port, mask16(0) => 
                           m16_0_port, Y(38) => y_38_port, Y(37) => y_37_port, 
                           Y(36) => y_36_port, Y(35) => y_35_port, Y(34) => 
                           y_34_port, Y(33) => y_33_port, Y(32) => y_32_port, 
                           Y(31) => y_31_port, Y(30) => y_30_port, Y(29) => 
                           y_29_port, Y(28) => y_28_port, Y(27) => y_27_port, 
                           Y(26) => y_26_port, Y(25) => y_25_port, Y(24) => 
                           y_24_port, Y(23) => y_23_port, Y(22) => y_22_port, 
                           Y(21) => y_21_port, Y(20) => y_20_port, Y(19) => 
                           y_19_port, Y(18) => y_18_port, Y(17) => y_17_port, 
                           Y(16) => y_16_port, Y(15) => y_15_port, Y(14) => 
                           y_14_port, Y(13) => y_13_port, Y(12) => y_12_port, 
                           Y(11) => y_11_port, Y(10) => y_10_port, Y(9) => 
                           y_9_port, Y(8) => y_8_port, Y(7) => y_7_port, Y(6) 
                           => y_6_port, Y(5) => y_5_port, Y(4) => y_4_port, 
                           Y(3) => y_3_port, Y(2) => y_2_port, Y(1) => y_1_port
                           , Y(0) => y_0_port);
   IIIL : shift_thirdLevel port map( sel(2) => s3_2_port, sel(1) => s3_1_port, 
                           sel(0) => s3_0_port, A(38) => y_38_port, A(37) => 
                           y_37_port, A(36) => y_36_port, A(35) => y_35_port, 
                           A(34) => y_34_port, A(33) => y_33_port, A(32) => 
                           y_32_port, A(31) => y_31_port, A(30) => y_30_port, 
                           A(29) => y_29_port, A(28) => y_28_port, A(27) => 
                           y_27_port, A(26) => y_26_port, A(25) => y_25_port, 
                           A(24) => y_24_port, A(23) => y_23_port, A(22) => 
                           y_22_port, A(21) => y_21_port, A(20) => y_20_port, 
                           A(19) => y_19_port, A(18) => y_18_port, A(17) => 
                           y_17_port, A(16) => y_16_port, A(15) => y_15_port, 
                           A(14) => y_14_port, A(13) => y_13_port, A(12) => 
                           y_12_port, A(11) => y_11_port, A(10) => y_10_port, 
                           A(9) => y_9_port, A(8) => y_8_port, A(7) => y_7_port
                           , A(6) => y_6_port, A(5) => y_5_port, A(4) => 
                           y_4_port, A(3) => y_3_port, A(2) => y_2_port, A(1) 
                           => y_1_port, A(0) => y_0_port, Y(31) => C(31), Y(30)
                           => C(30), Y(29) => C(29), Y(28) => C(28), Y(27) => 
                           C(27), Y(26) => C(26), Y(25) => C(25), Y(24) => 
                           C(24), Y(23) => C(23), Y(22) => C(22), Y(21) => 
                           C(21), Y(20) => C(20), Y(19) => C(19), Y(18) => 
                           C(18), Y(17) => C(17), Y(16) => C(16), Y(15) => 
                           C(15), Y(14) => C(14), Y(13) => C(13), Y(12) => 
                           C(12), Y(11) => C(11), Y(10) => C(10), Y(9) => C(9),
                           Y(8) => C(8), Y(7) => C(7), Y(6) => C(6), Y(5) => 
                           C(5), Y(4) => C(4), Y(3) => C(3), Y(2) => C(2), Y(1)
                           => C(1), Y(0) => C(0));
   U1 : AOI221_X1 port map( B1 => n6, B2 => n7, C1 => sel(0), C2 => B(2), A => 
                           n8, ZN => s3_2_port);
   U2 : INV_X1 port map( A => n6, ZN => n11);
   U3 : INV_X1 port map( A => B(2), ZN => n7);
   U4 : INV_X1 port map( A => n9, ZN => n8);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => sel(0), A => sel(1), ZN => n9);
   U6 : OAI22_X1 port map( A1 => B(0), A2 => n10, B1 => n11, B2 => n13, ZN => 
                           s3_0_port);
   U7 : INV_X1 port map( A => B(0), ZN => n13);
   U8 : OAI22_X1 port map( A1 => B(1), A2 => n10, B1 => n11, B2 => n12, ZN => 
                           s3_1_port);
   U9 : INV_X1 port map( A => B(1), ZN => n12);
   U10 : XNOR2_X1 port map( A => sel(1), B => sel(0), ZN => n10);
   U11 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n6);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity logical is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (3 downto 0);  Y : out std_logic_vector (31 downto 0));

end logical;

architecture SYN_behav of logical is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201 : 
      std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n121, A2 => n122, B1 => B(25), B2 => n123, ZN 
                           => Y(25));
   U2 : OAI22_X1 port map( A1 => n125, A2 => n126, B1 => B(24), B2 => n127, ZN 
                           => Y(24));
   U3 : OAI22_X1 port map( A1 => n129, A2 => n130, B1 => B(23), B2 => n131, ZN 
                           => Y(23));
   U4 : OAI22_X1 port map( A1 => n133, A2 => n134, B1 => B(22), B2 => n135, ZN 
                           => Y(22));
   U5 : OAI22_X1 port map( A1 => n137, A2 => n138, B1 => B(21), B2 => n139, ZN 
                           => Y(21));
   U6 : OAI22_X1 port map( A1 => n141, A2 => n142, B1 => B(20), B2 => n143, ZN 
                           => Y(20));
   U7 : OAI22_X1 port map( A1 => n149, A2 => n150, B1 => B(19), B2 => n151, ZN 
                           => Y(19));
   U8 : OAI22_X1 port map( A1 => n153, A2 => n154, B1 => B(18), B2 => n155, ZN 
                           => Y(18));
   U9 : OAI22_X1 port map( A1 => n157, A2 => n158, B1 => B(17), B2 => n159, ZN 
                           => Y(17));
   U10 : OAI22_X1 port map( A1 => n161, A2 => n162, B1 => B(16), B2 => n163, ZN
                           => Y(16));
   U11 : OAI22_X1 port map( A1 => n165, A2 => n166, B1 => B(15), B2 => n167, ZN
                           => Y(15));
   U12 : OAI22_X1 port map( A1 => n169, A2 => n170, B1 => B(14), B2 => n171, ZN
                           => Y(14));
   U13 : OAI22_X1 port map( A1 => n173, A2 => n174, B1 => B(13), B2 => n175, ZN
                           => Y(13));
   U14 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => B(7), B2 => n75, ZN => 
                           Y(7));
   U15 : OAI22_X1 port map( A1 => n77, A2 => n78, B1 => B(6), B2 => n79, ZN => 
                           Y(6));
   U16 : OAI22_X1 port map( A1 => n81, A2 => n82, B1 => B(5), B2 => n83, ZN => 
                           Y(5));
   U17 : OAI22_X1 port map( A1 => n85, A2 => n86, B1 => B(4), B2 => n87, ZN => 
                           Y(4));
   U18 : OAI22_X1 port map( A1 => n89, A2 => n90, B1 => B(3), B2 => n91, ZN => 
                           Y(3));
   U19 : OAI22_X1 port map( A1 => n101, A2 => n102, B1 => B(2), B2 => n103, ZN 
                           => Y(2));
   U20 : OAI22_X1 port map( A1 => n145, A2 => n146, B1 => B(1), B2 => n147, ZN 
                           => Y(1));
   U21 : OAI22_X1 port map( A1 => n93, A2 => n94, B1 => B(31), B2 => n95, ZN =>
                           Y(31));
   U22 : OAI22_X1 port map( A1 => n97, A2 => n98, B1 => B(30), B2 => n99, ZN =>
                           Y(30));
   U23 : OAI22_X1 port map( A1 => n105, A2 => n106, B1 => B(29), B2 => n107, ZN
                           => Y(29));
   U24 : OAI22_X1 port map( A1 => n109, A2 => n110, B1 => B(28), B2 => n111, ZN
                           => Y(28));
   U25 : OAI22_X1 port map( A1 => n113, A2 => n114, B1 => B(27), B2 => n115, ZN
                           => Y(27));
   U26 : OAI22_X1 port map( A1 => n117, A2 => n118, B1 => B(26), B2 => n119, ZN
                           => Y(26));
   U27 : OAI22_X1 port map( A1 => n177, A2 => n178, B1 => B(12), B2 => n179, ZN
                           => Y(12));
   U28 : OAI22_X1 port map( A1 => n181, A2 => n182, B1 => B(11), B2 => n183, ZN
                           => Y(11));
   U29 : OAI22_X1 port map( A1 => n185, A2 => n186, B1 => B(10), B2 => n187, ZN
                           => Y(10));
   U30 : OAI22_X1 port map( A1 => n65, A2 => n66, B1 => B(9), B2 => n67, ZN => 
                           Y(9));
   U31 : OAI22_X1 port map( A1 => n69, A2 => n70, B1 => B(8), B2 => n71, ZN => 
                           Y(8));
   U32 : BUF_X1 port map( A => sel(1), Z => n197);
   U33 : BUF_X1 port map( A => sel(0), Z => n194);
   U34 : BUF_X1 port map( A => sel(1), Z => n196);
   U35 : BUF_X1 port map( A => sel(0), Z => n193);
   U36 : OAI22_X1 port map( A1 => n189, A2 => n190, B1 => B(0), B2 => n191, ZN 
                           => Y(0));
   U37 : INV_X1 port map( A => B(0), ZN => n190);
   U38 : AOI22_X1 port map( A1 => n199, A2 => n192, B1 => A(0), B2 => n193, ZN 
                           => n189);
   U39 : AOI22_X1 port map( A1 => sel(3), A2 => n192, B1 => A(0), B2 => n196, 
                           ZN => n191);
   U40 : BUF_X1 port map( A => sel(2), Z => n200);
   U41 : BUF_X1 port map( A => sel(2), Z => n199);
   U42 : BUF_X1 port map( A => sel(1), Z => n198);
   U43 : BUF_X1 port map( A => sel(0), Z => n195);
   U44 : BUF_X1 port map( A => sel(2), Z => n201);
   U45 : AOI22_X1 port map( A1 => sel(3), A2 => n96, B1 => A(31), B2 => n198, 
                           ZN => n95);
   U46 : AOI22_X1 port map( A1 => sel(3), A2 => n72, B1 => A(8), B2 => n198, ZN
                           => n71);
   U47 : AOI22_X1 port map( A1 => sel(3), A2 => n76, B1 => A(7), B2 => n198, ZN
                           => n75);
   U48 : AOI22_X1 port map( A1 => sel(3), A2 => n80, B1 => A(6), B2 => n198, ZN
                           => n79);
   U49 : AOI22_X1 port map( A1 => sel(3), A2 => n84, B1 => A(5), B2 => n198, ZN
                           => n83);
   U50 : AOI22_X1 port map( A1 => sel(3), A2 => n88, B1 => A(4), B2 => n198, ZN
                           => n87);
   U51 : AOI22_X1 port map( A1 => sel(3), A2 => n92, B1 => A(3), B2 => n198, ZN
                           => n91);
   U52 : AOI22_X1 port map( A1 => sel(3), A2 => n68, B1 => n198, B2 => A(9), ZN
                           => n67);
   U53 : AOI22_X1 port map( A1 => sel(3), A2 => n100, B1 => A(30), B2 => n197, 
                           ZN => n99);
   U54 : AOI22_X1 port map( A1 => sel(3), A2 => n108, B1 => A(29), B2 => n197, 
                           ZN => n107);
   U55 : AOI22_X1 port map( A1 => sel(3), A2 => n112, B1 => A(28), B2 => n197, 
                           ZN => n111);
   U56 : AOI22_X1 port map( A1 => sel(3), A2 => n116, B1 => A(27), B2 => n197, 
                           ZN => n115);
   U57 : AOI22_X1 port map( A1 => sel(3), A2 => n120, B1 => A(26), B2 => n197, 
                           ZN => n119);
   U58 : AOI22_X1 port map( A1 => sel(3), A2 => n124, B1 => A(25), B2 => n197, 
                           ZN => n123);
   U59 : AOI22_X1 port map( A1 => sel(3), A2 => n128, B1 => A(24), B2 => n197, 
                           ZN => n127);
   U60 : AOI22_X1 port map( A1 => sel(3), A2 => n132, B1 => A(23), B2 => n197, 
                           ZN => n131);
   U61 : AOI22_X1 port map( A1 => sel(3), A2 => n136, B1 => A(22), B2 => n197, 
                           ZN => n135);
   U62 : AOI22_X1 port map( A1 => sel(3), A2 => n140, B1 => A(21), B2 => n197, 
                           ZN => n139);
   U63 : AOI22_X1 port map( A1 => sel(3), A2 => n144, B1 => A(20), B2 => n197, 
                           ZN => n143);
   U64 : AOI22_X1 port map( A1 => sel(3), A2 => n152, B1 => A(19), B2 => n196, 
                           ZN => n151);
   U65 : AOI22_X1 port map( A1 => sel(3), A2 => n156, B1 => A(18), B2 => n196, 
                           ZN => n155);
   U66 : AOI22_X1 port map( A1 => sel(3), A2 => n160, B1 => A(17), B2 => n196, 
                           ZN => n159);
   U67 : AOI22_X1 port map( A1 => sel(3), A2 => n164, B1 => A(16), B2 => n196, 
                           ZN => n163);
   U68 : AOI22_X1 port map( A1 => sel(3), A2 => n168, B1 => A(15), B2 => n196, 
                           ZN => n167);
   U69 : AOI22_X1 port map( A1 => sel(3), A2 => n172, B1 => A(14), B2 => n196, 
                           ZN => n171);
   U70 : AOI22_X1 port map( A1 => sel(3), A2 => n176, B1 => A(13), B2 => n196, 
                           ZN => n175);
   U71 : AOI22_X1 port map( A1 => sel(3), A2 => n180, B1 => A(12), B2 => n196, 
                           ZN => n179);
   U72 : AOI22_X1 port map( A1 => sel(3), A2 => n184, B1 => A(11), B2 => n196, 
                           ZN => n183);
   U73 : AOI22_X1 port map( A1 => sel(3), A2 => n188, B1 => A(10), B2 => n196, 
                           ZN => n187);
   U74 : AOI22_X1 port map( A1 => sel(3), A2 => n104, B1 => A(2), B2 => n197, 
                           ZN => n103);
   U75 : AOI22_X1 port map( A1 => sel(3), A2 => n148, B1 => A(1), B2 => n196, 
                           ZN => n147);
   U76 : AOI22_X1 port map( A1 => n201, A2 => n96, B1 => A(31), B2 => n195, ZN 
                           => n93);
   U77 : AOI22_X1 port map( A1 => n201, A2 => n72, B1 => A(8), B2 => n195, ZN 
                           => n69);
   U78 : AOI22_X1 port map( A1 => n201, A2 => n76, B1 => A(7), B2 => n195, ZN 
                           => n73);
   U79 : AOI22_X1 port map( A1 => n201, A2 => n80, B1 => A(6), B2 => n195, ZN 
                           => n77);
   U80 : AOI22_X1 port map( A1 => n201, A2 => n84, B1 => A(5), B2 => n195, ZN 
                           => n81);
   U81 : AOI22_X1 port map( A1 => n201, A2 => n88, B1 => A(4), B2 => n195, ZN 
                           => n85);
   U82 : AOI22_X1 port map( A1 => n201, A2 => n92, B1 => A(3), B2 => n195, ZN 
                           => n89);
   U83 : AOI22_X1 port map( A1 => n201, A2 => n68, B1 => n195, B2 => A(9), ZN 
                           => n65);
   U84 : AOI22_X1 port map( A1 => n200, A2 => n100, B1 => A(30), B2 => n194, ZN
                           => n97);
   U85 : AOI22_X1 port map( A1 => n200, A2 => n108, B1 => A(29), B2 => n194, ZN
                           => n105);
   U86 : AOI22_X1 port map( A1 => n200, A2 => n112, B1 => A(28), B2 => n194, ZN
                           => n109);
   U87 : AOI22_X1 port map( A1 => n200, A2 => n116, B1 => A(27), B2 => n194, ZN
                           => n113);
   U88 : AOI22_X1 port map( A1 => n200, A2 => n120, B1 => A(26), B2 => n194, ZN
                           => n117);
   U89 : AOI22_X1 port map( A1 => n200, A2 => n124, B1 => A(25), B2 => n194, ZN
                           => n121);
   U90 : AOI22_X1 port map( A1 => n200, A2 => n128, B1 => A(24), B2 => n194, ZN
                           => n125);
   U91 : AOI22_X1 port map( A1 => n200, A2 => n132, B1 => A(23), B2 => n194, ZN
                           => n129);
   U92 : AOI22_X1 port map( A1 => n200, A2 => n136, B1 => A(22), B2 => n194, ZN
                           => n133);
   U93 : AOI22_X1 port map( A1 => n200, A2 => n140, B1 => A(21), B2 => n194, ZN
                           => n137);
   U94 : AOI22_X1 port map( A1 => n200, A2 => n144, B1 => A(20), B2 => n194, ZN
                           => n141);
   U95 : AOI22_X1 port map( A1 => n199, A2 => n152, B1 => A(19), B2 => n193, ZN
                           => n149);
   U96 : AOI22_X1 port map( A1 => n199, A2 => n156, B1 => A(18), B2 => n193, ZN
                           => n153);
   U97 : AOI22_X1 port map( A1 => n199, A2 => n160, B1 => A(17), B2 => n193, ZN
                           => n157);
   U98 : AOI22_X1 port map( A1 => n199, A2 => n164, B1 => A(16), B2 => n193, ZN
                           => n161);
   U99 : AOI22_X1 port map( A1 => n199, A2 => n168, B1 => A(15), B2 => n193, ZN
                           => n165);
   U100 : AOI22_X1 port map( A1 => n199, A2 => n172, B1 => A(14), B2 => n193, 
                           ZN => n169);
   U101 : AOI22_X1 port map( A1 => n199, A2 => n176, B1 => A(13), B2 => n193, 
                           ZN => n173);
   U102 : AOI22_X1 port map( A1 => n199, A2 => n180, B1 => A(12), B2 => n193, 
                           ZN => n177);
   U103 : AOI22_X1 port map( A1 => n199, A2 => n184, B1 => A(11), B2 => n193, 
                           ZN => n181);
   U104 : AOI22_X1 port map( A1 => n199, A2 => n188, B1 => A(10), B2 => n193, 
                           ZN => n185);
   U105 : AOI22_X1 port map( A1 => n200, A2 => n104, B1 => A(2), B2 => n194, ZN
                           => n101);
   U106 : AOI22_X1 port map( A1 => n199, A2 => n148, B1 => A(1), B2 => n193, ZN
                           => n145);
   U107 : INV_X1 port map( A => A(9), ZN => n68);
   U108 : INV_X1 port map( A => A(31), ZN => n96);
   U109 : INV_X1 port map( A => A(30), ZN => n100);
   U110 : INV_X1 port map( A => A(29), ZN => n108);
   U111 : INV_X1 port map( A => A(28), ZN => n112);
   U112 : INV_X1 port map( A => A(27), ZN => n116);
   U113 : INV_X1 port map( A => A(26), ZN => n120);
   U114 : INV_X1 port map( A => A(25), ZN => n124);
   U115 : INV_X1 port map( A => A(24), ZN => n128);
   U116 : INV_X1 port map( A => A(23), ZN => n132);
   U117 : INV_X1 port map( A => A(22), ZN => n136);
   U118 : INV_X1 port map( A => A(21), ZN => n140);
   U119 : INV_X1 port map( A => A(20), ZN => n144);
   U120 : INV_X1 port map( A => A(19), ZN => n152);
   U121 : INV_X1 port map( A => A(18), ZN => n156);
   U122 : INV_X1 port map( A => A(17), ZN => n160);
   U123 : INV_X1 port map( A => A(16), ZN => n164);
   U124 : INV_X1 port map( A => A(15), ZN => n168);
   U125 : INV_X1 port map( A => A(14), ZN => n172);
   U126 : INV_X1 port map( A => A(13), ZN => n176);
   U127 : INV_X1 port map( A => A(12), ZN => n180);
   U128 : INV_X1 port map( A => A(11), ZN => n184);
   U129 : INV_X1 port map( A => A(10), ZN => n188);
   U130 : INV_X1 port map( A => A(8), ZN => n72);
   U131 : INV_X1 port map( A => A(7), ZN => n76);
   U132 : INV_X1 port map( A => A(6), ZN => n80);
   U133 : INV_X1 port map( A => A(5), ZN => n84);
   U134 : INV_X1 port map( A => A(4), ZN => n88);
   U135 : INV_X1 port map( A => A(3), ZN => n92);
   U136 : INV_X1 port map( A => A(2), ZN => n104);
   U137 : INV_X1 port map( A => A(1), ZN => n148);
   U138 : INV_X1 port map( A => A(0), ZN => n192);
   U139 : INV_X1 port map( A => B(31), ZN => n94);
   U140 : INV_X1 port map( A => B(30), ZN => n98);
   U141 : INV_X1 port map( A => B(29), ZN => n106);
   U142 : INV_X1 port map( A => B(28), ZN => n110);
   U143 : INV_X1 port map( A => B(27), ZN => n114);
   U144 : INV_X1 port map( A => B(26), ZN => n118);
   U145 : INV_X1 port map( A => B(25), ZN => n122);
   U146 : INV_X1 port map( A => B(24), ZN => n126);
   U147 : INV_X1 port map( A => B(23), ZN => n130);
   U148 : INV_X1 port map( A => B(22), ZN => n134);
   U149 : INV_X1 port map( A => B(21), ZN => n138);
   U150 : INV_X1 port map( A => B(20), ZN => n142);
   U151 : INV_X1 port map( A => B(19), ZN => n150);
   U152 : INV_X1 port map( A => B(18), ZN => n154);
   U153 : INV_X1 port map( A => B(17), ZN => n158);
   U154 : INV_X1 port map( A => B(16), ZN => n162);
   U155 : INV_X1 port map( A => B(15), ZN => n166);
   U156 : INV_X1 port map( A => B(14), ZN => n170);
   U157 : INV_X1 port map( A => B(13), ZN => n174);
   U158 : INV_X1 port map( A => B(12), ZN => n178);
   U159 : INV_X1 port map( A => B(11), ZN => n182);
   U160 : INV_X1 port map( A => B(10), ZN => n186);
   U161 : INV_X1 port map( A => B(9), ZN => n66);
   U162 : INV_X1 port map( A => B(8), ZN => n70);
   U163 : INV_X1 port map( A => B(7), ZN => n74);
   U164 : INV_X1 port map( A => B(6), ZN => n78);
   U165 : INV_X1 port map( A => B(5), ZN => n82);
   U166 : INV_X1 port map( A => B(4), ZN => n86);
   U167 : INV_X1 port map( A => B(3), ZN => n90);
   U168 : INV_X1 port map( A => B(2), ZN => n102);
   U169 : INV_X1 port map( A => B(1), ZN => n146);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity booth_mul_N16 is

   port( A, B : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end booth_mul_N16;

architecture SYN_struct of booth_mul_N16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component cla_adder_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_4
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_5
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux_N32_1
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_2
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_3
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_4
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_5
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_6
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_7
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_0
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component shift_mul_N16_S14
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S12
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S10
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S8
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S6
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S4
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S2
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S0
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, muxInE_7_31_port, muxInE_7_30_port, muxInE_7_29_port, 
      muxInE_7_28_port, muxInE_7_27_port, muxInE_7_26_port, muxInE_7_25_port, 
      muxInE_7_24_port, muxInE_7_23_port, muxInE_7_22_port, muxInE_7_21_port, 
      muxInE_7_20_port, muxInE_7_19_port, muxInE_7_18_port, muxInE_7_17_port, 
      muxInE_7_16_port, muxInE_7_15_port, muxInE_7_14_port, muxInE_7_13_port, 
      muxInE_7_12_port, muxInE_7_11_port, muxInE_7_10_port, muxInE_7_9_port, 
      muxInE_7_8_port, muxInE_7_7_port, muxInE_7_6_port, muxInE_7_5_port, 
      muxInE_7_4_port, muxInE_7_3_port, muxInE_7_2_port, muxInE_7_1_port, 
      muxInE_7_0_port, muxInE_6_31_port, muxInE_6_30_port, muxInE_6_29_port, 
      muxInE_6_28_port, muxInE_6_27_port, muxInE_6_26_port, muxInE_6_25_port, 
      muxInE_6_24_port, muxInE_6_23_port, muxInE_6_22_port, muxInE_6_21_port, 
      muxInE_6_20_port, muxInE_6_19_port, muxInE_6_18_port, muxInE_6_17_port, 
      muxInE_6_16_port, muxInE_6_15_port, muxInE_6_14_port, muxInE_6_13_port, 
      muxInE_6_12_port, muxInE_6_11_port, muxInE_6_10_port, muxInE_6_9_port, 
      muxInE_6_8_port, muxInE_6_7_port, muxInE_6_6_port, muxInE_6_5_port, 
      muxInE_6_4_port, muxInE_6_3_port, muxInE_6_2_port, muxInE_6_1_port, 
      muxInE_6_0_port, muxInE_5_31_port, muxInE_5_30_port, muxInE_5_29_port, 
      muxInE_5_28_port, muxInE_5_27_port, muxInE_5_26_port, muxInE_5_25_port, 
      muxInE_5_24_port, muxInE_5_23_port, muxInE_5_22_port, muxInE_5_21_port, 
      muxInE_5_20_port, muxInE_5_19_port, muxInE_5_18_port, muxInE_5_17_port, 
      muxInE_5_16_port, muxInE_5_15_port, muxInE_5_14_port, muxInE_5_13_port, 
      muxInE_5_12_port, muxInE_5_11_port, muxInE_5_10_port, muxInE_5_9_port, 
      muxInE_5_8_port, muxInE_5_7_port, muxInE_5_6_port, muxInE_5_5_port, 
      muxInE_5_4_port, muxInE_5_3_port, muxInE_5_2_port, muxInE_5_1_port, 
      muxInE_5_0_port, muxInE_4_31_port, muxInE_4_30_port, muxInE_4_29_port, 
      muxInE_4_28_port, muxInE_4_27_port, muxInE_4_26_port, muxInE_4_25_port, 
      muxInE_4_24_port, muxInE_4_23_port, muxInE_4_22_port, muxInE_4_21_port, 
      muxInE_4_20_port, muxInE_4_19_port, muxInE_4_18_port, muxInE_4_17_port, 
      muxInE_4_16_port, muxInE_4_15_port, muxInE_4_14_port, muxInE_4_13_port, 
      muxInE_4_12_port, muxInE_4_11_port, muxInE_4_10_port, muxInE_4_9_port, 
      muxInE_4_8_port, muxInE_4_7_port, muxInE_4_6_port, muxInE_4_5_port, 
      muxInE_4_4_port, muxInE_4_3_port, muxInE_4_2_port, muxInE_4_1_port, 
      muxInE_4_0_port, muxInE_3_31_port, muxInE_3_30_port, muxInE_3_29_port, 
      muxInE_3_28_port, muxInE_3_27_port, muxInE_3_26_port, muxInE_3_25_port, 
      muxInE_3_24_port, muxInE_3_23_port, muxInE_3_22_port, muxInE_3_21_port, 
      muxInE_3_20_port, muxInE_3_19_port, muxInE_3_18_port, muxInE_3_17_port, 
      muxInE_3_16_port, muxInE_3_15_port, muxInE_3_14_port, muxInE_3_13_port, 
      muxInE_3_12_port, muxInE_3_11_port, muxInE_3_10_port, muxInE_3_9_port, 
      muxInE_3_8_port, muxInE_3_7_port, muxInE_3_6_port, muxInE_3_5_port, 
      muxInE_3_4_port, muxInE_3_3_port, muxInE_3_2_port, muxInE_3_1_port, 
      muxInE_3_0_port, muxInE_2_31_port, muxInE_2_30_port, muxInE_2_29_port, 
      muxInE_2_28_port, muxInE_2_27_port, muxInE_2_26_port, muxInE_2_25_port, 
      muxInE_2_24_port, muxInE_2_23_port, muxInE_2_22_port, muxInE_2_21_port, 
      muxInE_2_19_port, muxInE_2_18_port, muxInE_2_17_port, muxInE_2_16_port, 
      muxInE_2_15_port, muxInE_2_14_port, muxInE_2_13_port, muxInE_2_12_port, 
      muxInE_2_11_port, muxInE_2_10_port, muxInE_2_9_port, muxInE_2_8_port, 
      muxInE_2_7_port, muxInE_2_6_port, muxInE_2_5_port, muxInE_2_4_port, 
      muxInE_2_3_port, muxInE_2_2_port, muxInE_2_1_port, muxInE_2_0_port, 
      muxInE_1_31_port, muxInE_1_30_port, muxInE_1_29_port, muxInE_1_28_port, 
      muxInE_1_27_port, muxInE_1_26_port, muxInE_1_25_port, muxInE_1_24_port, 
      muxInE_1_23_port, muxInE_1_22_port, muxInE_1_21_port, muxInE_1_20_port, 
      muxInE_1_19_port, muxInE_1_18_port, muxInE_1_17_port, muxInE_1_16_port, 
      muxInE_1_15_port, muxInE_1_14_port, muxInE_1_13_port, muxInE_1_12_port, 
      muxInE_1_11_port, muxInE_1_10_port, muxInE_1_9_port, muxInE_1_8_port, 
      muxInE_1_7_port, muxInE_1_6_port, muxInE_1_5_port, muxInE_1_4_port, 
      muxInE_1_3_port, muxInE_1_2_port, muxInE_1_1_port, muxInE_1_0_port, 
      muxInE_0_31_port, muxInE_0_30_port, muxInE_0_29_port, muxInE_0_28_port, 
      muxInE_0_27_port, muxInE_0_26_port, muxInE_0_24_port, muxInE_0_23_port, 
      muxInE_0_21_port, muxInE_0_20_port, muxInE_0_19_port, muxInE_0_18_port, 
      muxInE_0_16_port, muxInE_0_15_port, muxInE_0_14_port, muxInE_0_13_port, 
      muxInE_0_12_port, muxInE_0_11_port, muxInE_0_10_port, muxInE_0_9_port, 
      muxInE_0_8_port, muxInE_0_7_port, muxInE_0_6_port, muxInE_0_5_port, 
      muxInE_0_4_port, muxInE_0_3_port, muxInE_0_2_port, muxInE_0_1_port, 
      muxInE_0_0_port, muxInD_7_31_port, muxInD_7_30_port, muxInD_7_29_port, 
      muxInD_7_28_port, muxInD_7_27_port, muxInD_7_26_port, muxInD_7_25_port, 
      muxInD_7_24_port, muxInD_7_23_port, muxInD_7_22_port, muxInD_7_21_port, 
      muxInD_7_20_port, muxInD_7_19_port, muxInD_7_18_port, muxInD_7_17_port, 
      muxInD_7_16_port, muxInD_7_15_port, muxInD_7_14_port, muxInD_7_13_port, 
      muxInD_7_12_port, muxInD_7_11_port, muxInD_7_10_port, muxInD_7_9_port, 
      muxInD_7_8_port, muxInD_7_7_port, muxInD_7_6_port, muxInD_7_5_port, 
      muxInD_7_4_port, muxInD_7_3_port, muxInD_7_2_port, muxInD_7_1_port, 
      muxInD_7_0_port, muxInD_6_31_port, muxInD_6_30_port, muxInD_6_29_port, 
      muxInD_6_28_port, muxInD_6_27_port, muxInD_6_26_port, muxInD_6_25_port, 
      muxInD_6_24_port, muxInD_6_23_port, muxInD_6_22_port, muxInD_6_21_port, 
      muxInD_6_20_port, muxInD_6_19_port, muxInD_6_18_port, muxInD_6_17_port, 
      muxInD_6_16_port, muxInD_6_15_port, muxInD_6_14_port, muxInD_6_13_port, 
      muxInD_6_12_port, muxInD_6_11_port, muxInD_6_10_port, muxInD_6_9_port, 
      muxInD_6_8_port, muxInD_6_7_port, muxInD_6_6_port, muxInD_6_5_port, 
      muxInD_6_4_port, muxInD_6_3_port, muxInD_6_2_port, muxInD_6_1_port, 
      muxInD_6_0_port, muxInD_5_31_port, muxInD_5_30_port, muxInD_5_29_port, 
      muxInD_5_28_port, muxInD_5_27_port, muxInD_5_26_port, muxInD_5_25_port, 
      muxInD_5_24_port, muxInD_5_23_port, muxInD_5_22_port, muxInD_5_21_port, 
      muxInD_5_20_port, muxInD_5_19_port, muxInD_5_18_port, muxInD_5_17_port, 
      muxInD_5_16_port, muxInD_5_15_port, muxInD_5_14_port, muxInD_5_13_port, 
      muxInD_5_12_port, muxInD_5_11_port, muxInD_5_10_port, muxInD_5_9_port, 
      muxInD_5_8_port, muxInD_5_7_port, muxInD_5_6_port, muxInD_5_5_port, 
      muxInD_5_4_port, muxInD_5_3_port, muxInD_5_2_port, muxInD_5_1_port, 
      muxInD_5_0_port, muxInD_4_31_port, muxInD_4_30_port, muxInD_4_29_port, 
      muxInD_4_28_port, muxInD_4_27_port, muxInD_4_26_port, muxInD_4_25_port, 
      muxInD_4_24_port, muxInD_4_23_port, muxInD_4_22_port, muxInD_4_21_port, 
      muxInD_4_20_port, muxInD_4_19_port, muxInD_4_18_port, muxInD_4_17_port, 
      muxInD_4_16_port, muxInD_4_15_port, muxInD_4_14_port, muxInD_4_13_port, 
      muxInD_4_12_port, muxInD_4_11_port, muxInD_4_10_port, muxInD_4_9_port, 
      muxInD_4_8_port, muxInD_4_7_port, muxInD_4_6_port, muxInD_4_5_port, 
      muxInD_4_4_port, muxInD_4_3_port, muxInD_4_2_port, muxInD_4_1_port, 
      muxInD_4_0_port, muxInD_3_31_port, muxInD_3_30_port, muxInD_3_29_port, 
      muxInD_3_28_port, muxInD_3_27_port, muxInD_3_26_port, muxInD_3_25_port, 
      muxInD_3_24_port, muxInD_3_23_port, muxInD_3_22_port, muxInD_3_21_port, 
      muxInD_3_20_port, muxInD_3_19_port, muxInD_3_18_port, muxInD_3_17_port, 
      muxInD_3_16_port, muxInD_3_15_port, muxInD_3_14_port, muxInD_3_13_port, 
      muxInD_3_12_port, muxInD_3_11_port, muxInD_3_10_port, muxInD_3_9_port, 
      muxInD_3_8_port, muxInD_3_7_port, muxInD_3_6_port, muxInD_3_5_port, 
      muxInD_3_4_port, muxInD_3_3_port, muxInD_3_2_port, muxInD_3_1_port, 
      muxInD_3_0_port, muxInD_2_31_port, muxInD_2_30_port, muxInD_2_29_port, 
      muxInD_2_28_port, muxInD_2_27_port, muxInD_2_26_port, muxInD_2_25_port, 
      muxInD_2_24_port, muxInD_2_23_port, muxInD_2_22_port, muxInD_2_21_port, 
      muxInD_2_20_port, muxInD_2_19_port, muxInD_2_18_port, muxInD_2_17_port, 
      muxInD_2_16_port, muxInD_2_15_port, muxInD_2_14_port, muxInD_2_13_port, 
      muxInD_2_12_port, muxInD_2_11_port, muxInD_2_10_port, muxInD_2_9_port, 
      muxInD_2_8_port, muxInD_2_7_port, muxInD_2_6_port, muxInD_2_5_port, 
      muxInD_2_4_port, muxInD_2_3_port, muxInD_2_2_port, muxInD_2_1_port, 
      muxInD_2_0_port, muxInD_1_31_port, muxInD_1_30_port, muxInD_1_29_port, 
      muxInD_1_28_port, muxInD_1_27_port, muxInD_1_26_port, muxInD_1_25_port, 
      muxInD_1_24_port, muxInD_1_23_port, muxInD_1_22_port, muxInD_1_21_port, 
      muxInD_1_20_port, muxInD_1_19_port, muxInD_1_18_port, muxInD_1_17_port, 
      muxInD_1_16_port, muxInD_1_15_port, muxInD_1_14_port, muxInD_1_13_port, 
      muxInD_1_12_port, muxInD_1_11_port, muxInD_1_10_port, muxInD_1_9_port, 
      muxInD_1_8_port, muxInD_1_7_port, muxInD_1_6_port, muxInD_1_5_port, 
      muxInD_1_4_port, muxInD_1_3_port, muxInD_1_2_port, muxInD_1_1_port, 
      muxInD_1_0_port, muxInD_0_31_port, muxInD_0_30_port, muxInD_0_29_port, 
      muxInD_0_28_port, muxInD_0_27_port, muxInD_0_26_port, muxInD_0_25_port, 
      muxInD_0_24_port, muxInD_0_23_port, muxInD_0_22_port, muxInD_0_21_port, 
      muxInD_0_20_port, muxInD_0_19_port, muxInD_0_18_port, muxInD_0_17_port, 
      muxInD_0_16_port, muxInD_0_15_port, muxInD_0_14_port, muxInD_0_13_port, 
      muxInD_0_12_port, muxInD_0_11_port, muxInD_0_10_port, muxInD_0_9_port, 
      muxInD_0_8_port, muxInD_0_7_port, muxInD_0_6_port, muxInD_0_5_port, 
      muxInD_0_4_port, muxInD_0_3_port, muxInD_0_2_port, muxInD_0_1_port, 
      muxInD_0_0_port, muxInC_7_31_port, muxInC_7_30_port, muxInC_7_29_port, 
      muxInC_7_28_port, muxInC_7_27_port, muxInC_7_26_port, muxInC_7_25_port, 
      muxInC_7_24_port, muxInC_7_23_port, muxInC_7_22_port, muxInC_7_21_port, 
      muxInC_7_20_port, muxInC_7_19_port, muxInC_7_18_port, muxInC_7_17_port, 
      muxInC_7_16_port, muxInC_7_15_port, muxInC_7_14_port, muxInC_7_13_port, 
      muxInC_7_12_port, muxInC_7_11_port, muxInC_7_10_port, muxInC_7_9_port, 
      muxInC_7_8_port, muxInC_7_7_port, muxInC_7_6_port, muxInC_7_5_port, 
      muxInC_7_4_port, muxInC_7_3_port, muxInC_7_2_port, muxInC_7_1_port, 
      muxInC_7_0_port, muxInC_6_31_port, muxInC_6_30_port, muxInC_6_29_port, 
      muxInC_6_28_port, muxInC_6_27_port, muxInC_6_26_port, muxInC_6_25_port, 
      muxInC_6_24_port, muxInC_6_23_port, muxInC_6_22_port, muxInC_6_21_port, 
      muxInC_6_20_port, muxInC_6_19_port, muxInC_6_18_port, muxInC_6_17_port, 
      muxInC_6_16_port, muxInC_6_15_port, muxInC_6_14_port, muxInC_6_13_port, 
      muxInC_6_12_port, muxInC_6_11_port, muxInC_6_10_port, muxInC_6_9_port, 
      muxInC_6_8_port, muxInC_6_7_port, muxInC_6_6_port, muxInC_6_5_port, 
      muxInC_6_4_port, muxInC_6_3_port, muxInC_6_2_port, muxInC_6_1_port, 
      muxInC_6_0_port, muxInC_5_31_port, muxInC_5_30_port, muxInC_5_29_port, 
      muxInC_5_28_port, muxInC_5_27_port, muxInC_5_26_port, muxInC_5_25_port, 
      muxInC_5_24_port, muxInC_5_23_port, muxInC_5_22_port, muxInC_5_21_port, 
      muxInC_5_20_port, muxInC_5_19_port, muxInC_5_18_port, muxInC_5_17_port, 
      muxInC_5_16_port, muxInC_5_15_port, muxInC_5_14_port, muxInC_5_13_port, 
      muxInC_5_12_port, muxInC_5_11_port, muxInC_5_10_port, muxInC_5_9_port, 
      muxInC_5_8_port, muxInC_5_7_port, muxInC_5_6_port, muxInC_5_5_port, 
      muxInC_5_4_port, muxInC_5_3_port, muxInC_5_2_port, muxInC_5_1_port, 
      muxInC_5_0_port, muxInC_4_31_port, muxInC_4_30_port, muxInC_4_29_port, 
      muxInC_4_28_port, muxInC_4_27_port, muxInC_4_26_port, muxInC_4_25_port, 
      muxInC_4_24_port, muxInC_4_23_port, muxInC_4_22_port, muxInC_4_21_port, 
      muxInC_4_20_port, muxInC_4_19_port, muxInC_4_18_port, muxInC_4_17_port, 
      muxInC_4_16_port, muxInC_4_15_port, muxInC_4_14_port, muxInC_4_13_port, 
      muxInC_4_12_port, muxInC_4_11_port, muxInC_4_10_port, muxInC_4_9_port, 
      muxInC_4_8_port, muxInC_4_7_port, muxInC_4_6_port, muxInC_4_5_port, 
      muxInC_4_4_port, muxInC_4_3_port, muxInC_4_2_port, muxInC_4_1_port, 
      muxInC_4_0_port, muxInC_3_31_port, muxInC_3_30_port, muxInC_3_29_port, 
      muxInC_3_28_port, muxInC_3_27_port, muxInC_3_26_port, muxInC_3_25_port, 
      muxInC_3_24_port, muxInC_3_23_port, muxInC_3_22_port, muxInC_3_21_port, 
      muxInC_3_20_port, muxInC_3_19_port, muxInC_3_18_port, muxInC_3_17_port, 
      muxInC_3_16_port, muxInC_3_15_port, muxInC_3_14_port, muxInC_3_13_port, 
      muxInC_3_12_port, muxInC_3_11_port, muxInC_3_10_port, muxInC_3_9_port, 
      muxInC_3_8_port, muxInC_3_7_port, muxInC_3_6_port, muxInC_3_5_port, 
      muxInC_3_4_port, muxInC_3_3_port, muxInC_3_2_port, muxInC_3_1_port, 
      muxInC_3_0_port, muxInC_2_31_port, muxInC_2_30_port, muxInC_2_29_port, 
      muxInC_2_28_port, muxInC_2_27_port, muxInC_2_26_port, muxInC_2_25_port, 
      muxInC_2_24_port, muxInC_2_23_port, muxInC_2_22_port, muxInC_2_21_port, 
      muxInC_2_20_port, muxInC_2_19_port, muxInC_2_18_port, muxInC_2_17_port, 
      muxInC_2_16_port, muxInC_2_15_port, muxInC_2_14_port, muxInC_2_13_port, 
      muxInC_2_12_port, muxInC_2_11_port, muxInC_2_10_port, muxInC_2_9_port, 
      muxInC_2_8_port, muxInC_2_7_port, muxInC_2_6_port, muxInC_2_5_port, 
      muxInC_2_4_port, muxInC_2_3_port, muxInC_2_2_port, muxInC_2_1_port, 
      muxInC_2_0_port, muxInC_1_31_port, muxInC_1_30_port, muxInC_1_29_port, 
      muxInC_1_28_port, muxInC_1_27_port, muxInC_1_26_port, muxInC_1_25_port, 
      muxInC_1_24_port, muxInC_1_23_port, muxInC_1_22_port, muxInC_1_21_port, 
      muxInC_1_20_port, muxInC_1_18_port, muxInC_1_17_port, muxInC_1_16_port, 
      muxInC_1_15_port, muxInC_1_14_port, muxInC_1_13_port, muxInC_1_12_port, 
      muxInC_1_11_port, muxInC_1_10_port, muxInC_1_9_port, muxInC_1_8_port, 
      muxInC_1_7_port, muxInC_1_6_port, muxInC_1_5_port, muxInC_1_4_port, 
      muxInC_1_3_port, muxInC_1_2_port, muxInC_1_1_port, muxInC_1_0_port, 
      muxInC_0_31_port, muxInC_0_30_port, muxInC_0_29_port, muxInC_0_28_port, 
      muxInC_0_27_port, muxInC_0_26_port, muxInC_0_25_port, muxInC_0_24_port, 
      muxInC_0_23_port, muxInC_0_22_port, muxInC_0_21_port, muxInC_0_20_port, 
      muxInC_0_19_port, muxInC_0_18_port, muxInC_0_17_port, muxInC_0_16_port, 
      muxInC_0_15_port, muxInC_0_14_port, muxInC_0_13_port, muxInC_0_12_port, 
      muxInC_0_11_port, muxInC_0_10_port, muxInC_0_9_port, muxInC_0_8_port, 
      muxInC_0_7_port, muxInC_0_6_port, muxInC_0_5_port, muxInC_0_4_port, 
      muxInC_0_3_port, muxInC_0_2_port, muxInC_0_1_port, muxInC_0_0_port, 
      muxInB_7_31_port, muxInB_7_30_port, muxInB_7_29_port, muxInB_7_28_port, 
      muxInB_7_27_port, muxInB_7_26_port, muxInB_7_25_port, muxInB_7_24_port, 
      muxInB_7_23_port, muxInB_7_22_port, muxInB_7_21_port, muxInB_7_20_port, 
      muxInB_7_19_port, muxInB_7_18_port, muxInB_7_17_port, muxInB_7_16_port, 
      muxInB_7_15_port, muxInB_7_14_port, muxInB_7_13_port, muxInB_7_12_port, 
      muxInB_7_11_port, muxInB_7_10_port, muxInB_7_9_port, muxInB_7_8_port, 
      muxInB_7_7_port, muxInB_7_6_port, muxInB_7_5_port, muxInB_7_4_port, 
      muxInB_7_3_port, muxInB_7_2_port, muxInB_7_1_port, muxInB_7_0_port, 
      muxInB_6_31_port, muxInB_6_30_port, muxInB_6_29_port, muxInB_6_28_port, 
      muxInB_6_27_port, muxInB_6_26_port, muxInB_6_25_port, muxInB_6_24_port, 
      muxInB_6_23_port, muxInB_6_22_port, muxInB_6_21_port, muxInB_6_20_port, 
      muxInB_6_19_port, muxInB_6_18_port, muxInB_6_17_port, muxInB_6_16_port, 
      muxInB_6_15_port, muxInB_6_14_port, muxInB_6_13_port, muxInB_6_12_port, 
      muxInB_6_11_port, muxInB_6_10_port, muxInB_6_9_port, muxInB_6_8_port, 
      muxInB_6_7_port, muxInB_6_6_port, muxInB_6_5_port, muxInB_6_4_port, 
      muxInB_6_3_port, muxInB_6_2_port, muxInB_6_1_port, muxInB_6_0_port, 
      muxInB_5_31_port, muxInB_5_30_port, muxInB_5_29_port, muxInB_5_28_port, 
      muxInB_5_27_port, muxInB_5_26_port, muxInB_5_25_port, muxInB_5_24_port, 
      muxInB_5_23_port, muxInB_5_22_port, muxInB_5_21_port, muxInB_5_20_port, 
      muxInB_5_19_port, muxInB_5_18_port, muxInB_5_17_port, muxInB_5_16_port, 
      muxInB_5_15_port, muxInB_5_14_port, muxInB_5_13_port, muxInB_5_12_port, 
      muxInB_5_11_port, muxInB_5_10_port, muxInB_5_9_port, muxInB_5_8_port, 
      muxInB_5_7_port, muxInB_5_6_port, muxInB_5_5_port, muxInB_5_4_port, 
      muxInB_5_3_port, muxInB_5_2_port, muxInB_5_1_port, muxInB_5_0_port, 
      muxInB_4_31_port, muxInB_4_30_port, muxInB_4_29_port, muxInB_4_28_port, 
      muxInB_4_27_port, muxInB_4_26_port, muxInB_4_25_port, muxInB_4_24_port, 
      muxInB_4_23_port, muxInB_4_22_port, muxInB_4_21_port, muxInB_4_20_port, 
      muxInB_4_19_port, muxInB_4_18_port, muxInB_4_17_port, muxInB_4_16_port, 
      muxInB_4_15_port, muxInB_4_14_port, muxInB_4_13_port, muxInB_4_12_port, 
      muxInB_4_11_port, muxInB_4_10_port, muxInB_4_9_port, muxInB_4_8_port, 
      muxInB_4_7_port, muxInB_4_6_port, muxInB_4_5_port, muxInB_4_4_port, 
      muxInB_4_3_port, muxInB_4_2_port, muxInB_4_1_port, muxInB_4_0_port, 
      muxInB_3_31_port, muxInB_3_30_port, muxInB_3_29_port, muxInB_3_28_port, 
      muxInB_3_27_port, muxInB_3_26_port, muxInB_3_25_port, muxInB_3_24_port, 
      muxInB_3_23_port, muxInB_3_22_port, muxInB_3_21_port, muxInB_3_20_port, 
      muxInB_3_19_port, muxInB_3_18_port, muxInB_3_17_port, muxInB_3_16_port, 
      muxInB_3_15_port, muxInB_3_14_port, muxInB_3_13_port, muxInB_3_12_port, 
      muxInB_3_11_port, muxInB_3_10_port, muxInB_3_9_port, muxInB_3_8_port, 
      muxInB_3_7_port, muxInB_3_6_port, muxInB_3_5_port, muxInB_3_4_port, 
      muxInB_3_3_port, muxInB_3_2_port, muxInB_3_1_port, muxInB_3_0_port, 
      muxInB_2_31_port, muxInB_2_30_port, muxInB_2_29_port, muxInB_2_28_port, 
      muxInB_2_27_port, muxInB_2_26_port, muxInB_2_25_port, muxInB_2_24_port, 
      muxInB_2_23_port, muxInB_2_22_port, muxInB_2_21_port, muxInB_2_20_port, 
      muxInB_2_19_port, muxInB_2_18_port, muxInB_2_17_port, muxInB_2_16_port, 
      muxInB_2_15_port, muxInB_2_14_port, muxInB_2_13_port, muxInB_2_12_port, 
      muxInB_2_11_port, muxInB_2_10_port, muxInB_2_9_port, muxInB_2_8_port, 
      muxInB_2_7_port, muxInB_2_6_port, muxInB_2_5_port, muxInB_2_4_port, 
      muxInB_2_3_port, muxInB_2_2_port, muxInB_2_1_port, muxInB_2_0_port, 
      muxInB_1_31_port, muxInB_1_30_port, muxInB_1_29_port, muxInB_1_28_port, 
      muxInB_1_27_port, muxInB_1_26_port, muxInB_1_25_port, muxInB_1_24_port, 
      muxInB_1_23_port, muxInB_1_22_port, muxInB_1_21_port, muxInB_1_20_port, 
      muxInB_1_19_port, muxInB_1_18_port, muxInB_1_17_port, muxInB_1_16_port, 
      muxInB_1_15_port, muxInB_1_14_port, muxInB_1_13_port, muxInB_1_12_port, 
      muxInB_1_11_port, muxInB_1_10_port, muxInB_1_9_port, muxInB_1_8_port, 
      muxInB_1_7_port, muxInB_1_6_port, muxInB_1_5_port, muxInB_1_4_port, 
      muxInB_1_3_port, muxInB_1_2_port, muxInB_1_1_port, muxInB_1_0_port, 
      muxInB_0_31_port, muxInB_0_30_port, muxInB_0_29_port, muxInB_0_28_port, 
      muxInB_0_27_port, muxInB_0_26_port, muxInB_0_25_port, muxInB_0_24_port, 
      muxInB_0_23_port, muxInB_0_22_port, muxInB_0_21_port, muxInB_0_20_port, 
      muxInB_0_19_port, muxInB_0_18_port, muxInB_0_17_port, muxInB_0_16_port, 
      muxInB_0_15_port, muxInB_0_14_port, muxInB_0_13_port, muxInB_0_12_port, 
      muxInB_0_11_port, muxInB_0_10_port, muxInB_0_9_port, muxInB_0_8_port, 
      muxInB_0_7_port, muxInB_0_6_port, muxInB_0_5_port, muxInB_0_4_port, 
      muxInB_0_3_port, muxInB_0_2_port, muxInB_0_1_port, muxInB_0_0_port, 
      outmux_7_31_port, outmux_7_30_port, outmux_7_29_port, outmux_7_28_port, 
      outmux_7_27_port, outmux_7_26_port, outmux_7_25_port, outmux_7_24_port, 
      outmux_7_23_port, outmux_7_22_port, outmux_7_21_port, outmux_7_20_port, 
      outmux_7_19_port, outmux_7_18_port, outmux_7_17_port, outmux_7_16_port, 
      outmux_7_15_port, outmux_7_14_port, outmux_7_13_port, outmux_7_12_port, 
      outmux_7_11_port, outmux_7_10_port, outmux_7_9_port, outmux_7_8_port, 
      outmux_7_7_port, outmux_7_6_port, outmux_7_5_port, outmux_7_4_port, 
      outmux_7_3_port, outmux_7_2_port, outmux_7_1_port, outmux_7_0_port, 
      outmux_6_31_port, outmux_6_30_port, outmux_6_29_port, outmux_6_28_port, 
      outmux_6_27_port, outmux_6_26_port, outmux_6_25_port, outmux_6_24_port, 
      outmux_6_23_port, outmux_6_22_port, outmux_6_21_port, outmux_6_20_port, 
      outmux_6_19_port, outmux_6_18_port, outmux_6_17_port, outmux_6_16_port, 
      outmux_6_15_port, outmux_6_14_port, outmux_6_13_port, outmux_6_12_port, 
      outmux_6_11_port, outmux_6_10_port, outmux_6_9_port, outmux_6_8_port, 
      outmux_6_7_port, outmux_6_6_port, outmux_6_5_port, outmux_6_4_port, 
      outmux_6_3_port, outmux_6_2_port, outmux_6_1_port, outmux_6_0_port, 
      outmux_5_31_port, outmux_5_30_port, outmux_5_29_port, outmux_5_28_port, 
      outmux_5_27_port, outmux_5_26_port, outmux_5_25_port, outmux_5_24_port, 
      outmux_5_23_port, outmux_5_22_port, outmux_5_21_port, outmux_5_20_port, 
      outmux_5_19_port, outmux_5_18_port, outmux_5_17_port, outmux_5_16_port, 
      outmux_5_15_port, outmux_5_14_port, outmux_5_13_port, outmux_5_12_port, 
      outmux_5_11_port, outmux_5_10_port, outmux_5_9_port, outmux_5_8_port, 
      outmux_5_7_port, outmux_5_6_port, outmux_5_5_port, outmux_5_4_port, 
      outmux_5_3_port, outmux_5_2_port, outmux_5_1_port, outmux_5_0_port, 
      outmux_4_31_port, outmux_4_30_port, outmux_4_29_port, outmux_4_28_port, 
      outmux_4_27_port, outmux_4_26_port, outmux_4_25_port, outmux_4_24_port, 
      outmux_4_23_port, outmux_4_22_port, outmux_4_21_port, outmux_4_20_port, 
      outmux_4_19_port, outmux_4_18_port, outmux_4_17_port, outmux_4_16_port, 
      outmux_4_15_port, outmux_4_14_port, outmux_4_13_port, outmux_4_12_port, 
      outmux_4_11_port, outmux_4_10_port, outmux_4_9_port, outmux_4_8_port, 
      outmux_4_7_port, outmux_4_6_port, outmux_4_5_port, outmux_4_4_port, 
      outmux_4_3_port, outmux_4_2_port, outmux_4_1_port, outmux_4_0_port, 
      outmux_3_31_port, outmux_3_30_port, outmux_3_29_port, outmux_3_28_port, 
      outmux_3_27_port, outmux_3_26_port, outmux_3_25_port, outmux_3_24_port, 
      outmux_3_23_port, outmux_3_22_port, outmux_3_21_port, outmux_3_20_port, 
      outmux_3_19_port, outmux_3_18_port, outmux_3_17_port, outmux_3_16_port, 
      outmux_3_15_port, outmux_3_14_port, outmux_3_13_port, outmux_3_12_port, 
      outmux_3_11_port, outmux_3_10_port, outmux_3_9_port, outmux_3_8_port, 
      outmux_3_7_port, outmux_3_6_port, outmux_3_5_port, outmux_3_4_port, 
      outmux_3_3_port, outmux_3_2_port, outmux_3_1_port, outmux_3_0_port, 
      outmux_2_31_port, outmux_2_30_port, outmux_2_29_port, outmux_2_28_port, 
      outmux_2_27_port, outmux_2_26_port, outmux_2_25_port, outmux_2_24_port, 
      outmux_2_23_port, outmux_2_22_port, outmux_2_21_port, outmux_2_20_port, 
      outmux_2_19_port, outmux_2_18_port, outmux_2_17_port, outmux_2_16_port, 
      outmux_2_15_port, outmux_2_14_port, outmux_2_13_port, outmux_2_12_port, 
      outmux_2_11_port, outmux_2_10_port, outmux_2_9_port, outmux_2_8_port, 
      outmux_2_7_port, outmux_2_6_port, outmux_2_5_port, outmux_2_4_port, 
      outmux_2_3_port, outmux_2_2_port, outmux_2_1_port, outmux_2_0_port, 
      outmux_1_31_port, outmux_1_30_port, outmux_1_29_port, outmux_1_28_port, 
      outmux_1_27_port, outmux_1_26_port, outmux_1_25_port, outmux_1_24_port, 
      outmux_1_23_port, outmux_1_22_port, outmux_1_21_port, outmux_1_20_port, 
      outmux_1_19_port, outmux_1_18_port, outmux_1_17_port, outmux_1_16_port, 
      outmux_1_15_port, outmux_1_14_port, outmux_1_13_port, outmux_1_12_port, 
      outmux_1_11_port, outmux_1_10_port, outmux_1_9_port, outmux_1_8_port, 
      outmux_1_7_port, outmux_1_6_port, outmux_1_5_port, outmux_1_4_port, 
      outmux_1_3_port, outmux_1_2_port, outmux_1_1_port, outmux_1_0_port, 
      outmux_0_31_port, outmux_0_30_port, outmux_0_29_port, outmux_0_28_port, 
      outmux_0_27_port, outmux_0_26_port, outmux_0_25_port, outmux_0_24_port, 
      outmux_0_23_port, outmux_0_22_port, outmux_0_21_port, outmux_0_20_port, 
      outmux_0_19_port, outmux_0_18_port, outmux_0_17_port, outmux_0_16_port, 
      outmux_0_15_port, outmux_0_14_port, outmux_0_13_port, outmux_0_12_port, 
      outmux_0_11_port, outmux_0_10_port, outmux_0_9_port, outmux_0_8_port, 
      outmux_0_7_port, outmux_0_6_port, outmux_0_5_port, outmux_0_4_port, 
      outmux_0_3_port, outmux_0_2_port, outmux_0_1_port, outmux_0_0_port, 
      cout_array_5_31_port, cout_array_5_30_port, cout_array_5_29_port, 
      cout_array_5_28_port, cout_array_5_27_port, cout_array_5_26_port, 
      cout_array_5_25_port, cout_array_5_24_port, cout_array_5_23_port, 
      cout_array_5_22_port, cout_array_5_21_port, cout_array_5_20_port, 
      cout_array_5_19_port, cout_array_5_18_port, cout_array_5_17_port, 
      cout_array_5_16_port, cout_array_5_15_port, cout_array_5_14_port, 
      cout_array_5_13_port, cout_array_5_12_port, cout_array_5_11_port, 
      cout_array_5_10_port, cout_array_5_9_port, cout_array_5_8_port, 
      cout_array_5_7_port, cout_array_5_6_port, cout_array_5_5_port, 
      cout_array_5_4_port, cout_array_5_3_port, cout_array_5_2_port, 
      cout_array_5_1_port, cout_array_5_0_port, cout_array_4_31_port, 
      cout_array_4_30_port, cout_array_4_29_port, cout_array_4_28_port, 
      cout_array_4_27_port, cout_array_4_26_port, cout_array_4_25_port, 
      cout_array_4_24_port, cout_array_4_23_port, cout_array_4_22_port, 
      cout_array_4_21_port, cout_array_4_20_port, cout_array_4_19_port, 
      cout_array_4_18_port, cout_array_4_17_port, cout_array_4_16_port, 
      cout_array_4_15_port, cout_array_4_14_port, cout_array_4_13_port, 
      cout_array_4_12_port, cout_array_4_11_port, cout_array_4_10_port, 
      cout_array_4_9_port, cout_array_4_8_port, cout_array_4_7_port, 
      cout_array_4_6_port, cout_array_4_5_port, cout_array_4_4_port, 
      cout_array_4_3_port, cout_array_4_2_port, cout_array_4_1_port, 
      cout_array_4_0_port, cout_array_3_31_port, cout_array_3_30_port, 
      cout_array_3_29_port, cout_array_3_28_port, cout_array_3_27_port, 
      cout_array_3_26_port, cout_array_3_25_port, cout_array_3_24_port, 
      cout_array_3_23_port, cout_array_3_22_port, cout_array_3_21_port, 
      cout_array_3_20_port, cout_array_3_19_port, cout_array_3_18_port, 
      cout_array_3_17_port, cout_array_3_16_port, cout_array_3_15_port, 
      cout_array_3_14_port, cout_array_3_13_port, cout_array_3_12_port, 
      cout_array_3_11_port, cout_array_3_10_port, cout_array_3_9_port, 
      cout_array_3_8_port, cout_array_3_7_port, cout_array_3_6_port, 
      cout_array_3_5_port, cout_array_3_4_port, cout_array_3_3_port, 
      cout_array_3_2_port, cout_array_3_1_port, cout_array_3_0_port, 
      cout_array_2_31_port, cout_array_2_30_port, cout_array_2_29_port, 
      cout_array_2_28_port, cout_array_2_27_port, cout_array_2_26_port, 
      cout_array_2_25_port, cout_array_2_24_port, cout_array_2_23_port, 
      cout_array_2_22_port, cout_array_2_21_port, cout_array_2_20_port, 
      cout_array_2_19_port, cout_array_2_18_port, cout_array_2_17_port, 
      cout_array_2_16_port, cout_array_2_15_port, cout_array_2_14_port, 
      cout_array_2_13_port, cout_array_2_12_port, cout_array_2_11_port, 
      cout_array_2_10_port, cout_array_2_9_port, cout_array_2_8_port, 
      cout_array_2_7_port, cout_array_2_6_port, cout_array_2_5_port, 
      cout_array_2_4_port, cout_array_2_3_port, cout_array_2_2_port, 
      cout_array_2_1_port, cout_array_2_0_port, cout_array_1_31_port, 
      cout_array_1_30_port, cout_array_1_29_port, cout_array_1_28_port, 
      cout_array_1_27_port, cout_array_1_26_port, cout_array_1_25_port, 
      cout_array_1_24_port, cout_array_1_23_port, cout_array_1_22_port, 
      cout_array_1_21_port, cout_array_1_20_port, cout_array_1_19_port, 
      cout_array_1_18_port, cout_array_1_17_port, cout_array_1_16_port, 
      cout_array_1_15_port, cout_array_1_14_port, cout_array_1_13_port, 
      cout_array_1_12_port, cout_array_1_11_port, cout_array_1_10_port, 
      cout_array_1_9_port, cout_array_1_8_port, cout_array_1_7_port, 
      cout_array_1_6_port, cout_array_1_5_port, cout_array_1_4_port, 
      cout_array_1_3_port, cout_array_1_2_port, cout_array_1_1_port, 
      cout_array_1_0_port, cout_array_0_31_port, cout_array_0_30_port, 
      cout_array_0_29_port, cout_array_0_28_port, cout_array_0_27_port, 
      cout_array_0_26_port, cout_array_0_25_port, cout_array_0_24_port, 
      cout_array_0_23_port, cout_array_0_22_port, cout_array_0_21_port, 
      cout_array_0_20_port, cout_array_0_19_port, cout_array_0_18_port, 
      cout_array_0_17_port, cout_array_0_16_port, cout_array_0_15_port, 
      cout_array_0_14_port, cout_array_0_13_port, cout_array_0_12_port, 
      cout_array_0_11_port, cout_array_0_10_port, cout_array_0_9_port, 
      cout_array_0_8_port, cout_array_0_7_port, cout_array_0_6_port, 
      cout_array_0_5_port, cout_array_0_4_port, cout_array_0_3_port, 
      cout_array_0_2_port, cout_array_0_1_port, cout_array_0_0_port, 
      sum_array_5_31_port, sum_array_5_30_port, sum_array_5_29_port, 
      sum_array_5_28_port, sum_array_5_27_port, sum_array_5_26_port, 
      sum_array_5_25_port, sum_array_5_24_port, sum_array_5_23_port, 
      sum_array_5_22_port, sum_array_5_21_port, sum_array_5_20_port, 
      sum_array_5_19_port, sum_array_5_18_port, sum_array_5_17_port, 
      sum_array_5_16_port, sum_array_5_15_port, sum_array_5_14_port, 
      sum_array_5_13_port, sum_array_5_12_port, sum_array_5_11_port, 
      sum_array_5_10_port, sum_array_5_9_port, sum_array_5_8_port, 
      sum_array_5_7_port, sum_array_5_6_port, sum_array_5_5_port, 
      sum_array_5_4_port, sum_array_5_3_port, sum_array_5_2_port, 
      sum_array_5_1_port, sum_array_5_0_port, sum_array_4_31_port, 
      sum_array_4_30_port, sum_array_4_29_port, sum_array_4_28_port, 
      sum_array_4_27_port, sum_array_4_26_port, sum_array_4_25_port, 
      sum_array_4_24_port, sum_array_4_23_port, sum_array_4_22_port, 
      sum_array_4_21_port, sum_array_4_20_port, sum_array_4_19_port, 
      sum_array_4_18_port, sum_array_4_17_port, sum_array_4_16_port, 
      sum_array_4_15_port, sum_array_4_14_port, sum_array_4_13_port, 
      sum_array_4_12_port, sum_array_4_11_port, sum_array_4_10_port, 
      sum_array_4_9_port, sum_array_4_8_port, sum_array_4_7_port, 
      sum_array_4_6_port, sum_array_4_5_port, sum_array_4_4_port, 
      sum_array_4_3_port, sum_array_4_2_port, sum_array_4_1_port, 
      sum_array_4_0_port, sum_array_3_31_port, sum_array_3_30_port, 
      sum_array_3_29_port, sum_array_3_28_port, sum_array_3_27_port, 
      sum_array_3_26_port, sum_array_3_25_port, sum_array_3_24_port, 
      sum_array_3_23_port, sum_array_3_22_port, sum_array_3_21_port, 
      sum_array_3_20_port, sum_array_3_19_port, sum_array_3_18_port, 
      sum_array_3_17_port, sum_array_3_16_port, sum_array_3_15_port, 
      sum_array_3_14_port, sum_array_3_13_port, sum_array_3_12_port, 
      sum_array_3_11_port, sum_array_3_10_port, sum_array_3_9_port, 
      sum_array_3_8_port, sum_array_3_7_port, sum_array_3_6_port, 
      sum_array_3_5_port, sum_array_3_4_port, sum_array_3_3_port, 
      sum_array_3_2_port, sum_array_3_1_port, sum_array_3_0_port, 
      sum_array_2_31_port, sum_array_2_30_port, sum_array_2_29_port, 
      sum_array_2_28_port, sum_array_2_27_port, sum_array_2_26_port, 
      sum_array_2_25_port, sum_array_2_24_port, sum_array_2_23_port, 
      sum_array_2_22_port, sum_array_2_21_port, sum_array_2_20_port, 
      sum_array_2_19_port, sum_array_2_18_port, sum_array_2_17_port, 
      sum_array_2_16_port, sum_array_2_15_port, sum_array_2_14_port, 
      sum_array_2_13_port, sum_array_2_12_port, sum_array_2_11_port, 
      sum_array_2_10_port, sum_array_2_9_port, sum_array_2_8_port, 
      sum_array_2_7_port, sum_array_2_6_port, sum_array_2_5_port, 
      sum_array_2_4_port, sum_array_2_3_port, sum_array_2_2_port, 
      sum_array_2_1_port, sum_array_2_0_port, sum_array_1_31_port, 
      sum_array_1_30_port, sum_array_1_29_port, sum_array_1_28_port, 
      sum_array_1_27_port, sum_array_1_26_port, sum_array_1_25_port, 
      sum_array_1_24_port, sum_array_1_23_port, sum_array_1_22_port, 
      sum_array_1_21_port, sum_array_1_20_port, sum_array_1_19_port, 
      sum_array_1_18_port, sum_array_1_17_port, sum_array_1_16_port, 
      sum_array_1_15_port, sum_array_1_14_port, sum_array_1_13_port, 
      sum_array_1_12_port, sum_array_1_11_port, sum_array_1_10_port, 
      sum_array_1_9_port, sum_array_1_8_port, sum_array_1_7_port, 
      sum_array_1_6_port, sum_array_1_5_port, sum_array_1_4_port, 
      sum_array_1_3_port, sum_array_1_2_port, sum_array_1_1_port, 
      sum_array_1_0_port, sum_array_0_31_port, sum_array_0_30_port, 
      sum_array_0_29_port, sum_array_0_28_port, sum_array_0_27_port, 
      sum_array_0_26_port, sum_array_0_25_port, sum_array_0_24_port, 
      sum_array_0_23_port, sum_array_0_22_port, sum_array_0_21_port, 
      sum_array_0_20_port, sum_array_0_19_port, sum_array_0_18_port, 
      sum_array_0_17_port, sum_array_0_16_port, sum_array_0_15_port, 
      sum_array_0_14_port, sum_array_0_13_port, sum_array_0_12_port, 
      sum_array_0_11_port, sum_array_0_10_port, sum_array_0_9_port, 
      sum_array_0_8_port, sum_array_0_7_port, sum_array_0_6_port, 
      sum_array_0_5_port, sum_array_0_4_port, sum_array_0_3_port, 
      sum_array_0_2_port, sum_array_0_1_port, sum_array_0_0_port, net6197, n20,
      net51440, net51450, net51451, net51452, n2, n3, n10, n11, n13, n14, n15, 
      n17, n18, n19, n21, n22, n25, n26, n27, n28, net59829, net59830, net59831
      , net59832, net59833, net59834, net59835, net59836, net59837, net59838, 
      net59839, net59840, net59841, net59842, net59843, net59844, net59845, 
      net59846, net59847, net59848, net59849, net59850, net59851, net59852, 
      net59853, net59854, net59855, net59856, net59857, net59858, net59859, 
      net59860, net59861, net59862, net59863, net59864, net59865, net59866, 
      net59867, net59868, net59869, net59870, net59871, net59872, net59873, 
      net59874, net59875, net59876, net59877, net59878, net59879, net59880, 
      net59881, net59882, net59883, net59884, net59885, net59886, net59887, 
      net59888, net59889, net59890, net59891, net59892, net59893, net59894, 
      net59895, net59896, net59897, net59898, net59899, net59900, net59901, 
      net59902, net59903, net59904, net59905, net59906, net59907, net59908, 
      net59909, net59910, net59911, net59912, net59913, net59914, net59915, 
      net59916, net59917, net59918, net59919, net59920, net59921, net59922, 
      net59923, net59924, net59925, net59926, net59927, net59928, net59929, 
      net59930, net59931, net59932, net59933, net59934, net59935, net59936, 
      net59937, net59938, net59939, net59940, net59941, net59942, net59943, 
      net59944, net59945, net59946, net59947, net59948, net59949, net59950, 
      net59951, net59952, net59953, net59954, net59955, net59956, net59957, 
      net59958, net59959, net59960, net59961, net59962, net59963, net59964, 
      net59965, net59966, net59967, net59968, net59969, net59970, net59971, 
      net59972, net59973, net59974, net59975, net59976, net59977, net59978, 
      net59979, net59980, net59981, net59982, net59983, net59984, net59985, 
      net59986, net59987, net59988, net59989, net59990, net59991, net59992, 
      net59993, net59994, net59995, net59996, net59997, net59998, net59999, 
      net60000, net60001, net60002, net60003, net60004, net60005, net60006, 
      net60007, net60008, net60009, net60010, net60011, net60012, net60013, 
      net60014, net60015, net60016, net60017, net60018, net60019, net60020, 
      net60021, net60022, net60023, net60024, net60025, net60026, net60027, 
      net60028, net60029, net60030, net60031, net60032, net60033, net60034, 
      net60035, net60036, net60037, net60038, net60039, net60040, net60041, 
      net60042, net60043, net60044, net60045, net60046, net60047, net60048, 
      net60049, net60050, net60051, net60052, net60053, net60054, net60055, 
      net60056, net60057, net60058, net60059, net60060, net60061, net60062, 
      net60063, net60064, net60065, net60066, net60067, net60068, net60069, 
      net60070, net60071, net60072, net60073, net60074 : std_logic;

begin
   
   X_Logic0_port <= '0';
   SHIFTERS_0 : shift_mul_N16_S0 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_0_31_port, B(30)
                           => muxInB_0_30_port, B(29) => muxInB_0_29_port, 
                           B(28) => muxInB_0_28_port, B(27) => muxInB_0_27_port
                           , B(26) => muxInB_0_26_port, B(25) => 
                           muxInB_0_25_port, B(24) => muxInB_0_24_port, B(23) 
                           => muxInB_0_23_port, B(22) => muxInB_0_22_port, 
                           B(21) => muxInB_0_21_port, B(20) => muxInB_0_20_port
                           , B(19) => muxInB_0_19_port, B(18) => 
                           muxInB_0_18_port, B(17) => muxInB_0_17_port, B(16) 
                           => muxInB_0_16_port, B(15) => muxInB_0_15_port, 
                           B(14) => muxInB_0_14_port, B(13) => muxInB_0_13_port
                           , B(12) => muxInB_0_12_port, B(11) => 
                           muxInB_0_11_port, B(10) => muxInB_0_10_port, B(9) =>
                           muxInB_0_9_port, B(8) => muxInB_0_8_port, B(7) => 
                           muxInB_0_7_port, B(6) => muxInB_0_6_port, B(5) => 
                           muxInB_0_5_port, B(4) => muxInB_0_4_port, B(3) => 
                           muxInB_0_3_port, B(2) => muxInB_0_2_port, B(1) => 
                           muxInB_0_1_port, B(0) => muxInB_0_0_port, C(31) => 
                           muxInC_0_31_port, C(30) => muxInC_0_30_port, C(29) 
                           => muxInC_0_29_port, C(28) => muxInC_0_28_port, 
                           C(27) => muxInC_0_27_port, C(26) => muxInC_0_26_port
                           , C(25) => muxInC_0_25_port, C(24) => 
                           muxInC_0_24_port, C(23) => muxInC_0_23_port, C(22) 
                           => muxInC_0_22_port, C(21) => muxInC_0_21_port, 
                           C(20) => muxInC_0_20_port, C(19) => muxInC_0_19_port
                           , C(18) => muxInC_0_18_port, C(17) => 
                           muxInC_0_17_port, C(16) => muxInC_0_16_port, C(15) 
                           => muxInC_0_15_port, C(14) => muxInC_0_14_port, 
                           C(13) => muxInC_0_13_port, C(12) => muxInC_0_12_port
                           , C(11) => muxInC_0_11_port, C(10) => 
                           muxInC_0_10_port, C(9) => muxInC_0_9_port, C(8) => 
                           muxInC_0_8_port, C(7) => muxInC_0_7_port, C(6) => 
                           muxInC_0_6_port, C(5) => muxInC_0_5_port, C(4) => 
                           muxInC_0_4_port, C(3) => muxInC_0_3_port, C(2) => 
                           muxInC_0_2_port, C(1) => muxInC_0_1_port, C(0) => 
                           muxInC_0_0_port, D(31) => muxInD_0_31_port, D(30) =>
                           muxInD_0_30_port, D(29) => muxInD_0_29_port, D(28) 
                           => muxInD_0_28_port, D(27) => muxInD_0_27_port, 
                           D(26) => muxInD_0_26_port, D(25) => muxInD_0_25_port
                           , D(24) => muxInD_0_24_port, D(23) => 
                           muxInD_0_23_port, D(22) => muxInD_0_22_port, D(21) 
                           => muxInD_0_21_port, D(20) => muxInD_0_20_port, 
                           D(19) => muxInD_0_19_port, D(18) => muxInD_0_18_port
                           , D(17) => muxInD_0_17_port, D(16) => 
                           muxInD_0_16_port, D(15) => muxInD_0_15_port, D(14) 
                           => muxInD_0_14_port, D(13) => muxInD_0_13_port, 
                           D(12) => muxInD_0_12_port, D(11) => muxInD_0_11_port
                           , D(10) => muxInD_0_10_port, D(9) => muxInD_0_9_port
                           , D(8) => muxInD_0_8_port, D(7) => muxInD_0_7_port, 
                           D(6) => muxInD_0_6_port, D(5) => muxInD_0_5_port, 
                           D(4) => muxInD_0_4_port, D(3) => muxInD_0_3_port, 
                           D(2) => muxInD_0_2_port, D(1) => muxInD_0_1_port, 
                           D(0) => net60073, E(31) => muxInE_0_31_port, E(30) 
                           => muxInE_0_30_port, E(29) => muxInE_0_29_port, 
                           E(28) => muxInE_0_28_port, E(27) => muxInE_0_27_port
                           , E(26) => muxInE_0_26_port, E(25) => net51450, 
                           E(24) => muxInE_0_24_port, E(23) => muxInE_0_23_port
                           , E(22) => net51451, E(21) => muxInE_0_21_port, 
                           E(20) => muxInE_0_20_port, E(19) => muxInE_0_19_port
                           , E(18) => muxInE_0_18_port, E(17) => net51452, 
                           E(16) => muxInE_0_16_port, E(15) => muxInE_0_15_port
                           , E(14) => muxInE_0_14_port, E(13) => 
                           muxInE_0_13_port, E(12) => muxInE_0_12_port, E(11) 
                           => muxInE_0_11_port, E(10) => muxInE_0_10_port, E(9)
                           => muxInE_0_9_port, E(8) => muxInE_0_8_port, E(7) =>
                           muxInE_0_7_port, E(6) => muxInE_0_6_port, E(5) => 
                           muxInE_0_5_port, E(4) => muxInE_0_4_port, E(3) => 
                           muxInE_0_3_port, E(2) => muxInE_0_2_port, E(1) => 
                           muxInE_0_1_port, E(0) => net60074);
   SHIFTERS_1 : shift_mul_N16_S2 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_1_31_port, B(30)
                           => muxInB_1_30_port, B(29) => muxInB_1_29_port, 
                           B(28) => muxInB_1_28_port, B(27) => muxInB_1_27_port
                           , B(26) => muxInB_1_26_port, B(25) => 
                           muxInB_1_25_port, B(24) => muxInB_1_24_port, B(23) 
                           => muxInB_1_23_port, B(22) => muxInB_1_22_port, 
                           B(21) => muxInB_1_21_port, B(20) => muxInB_1_20_port
                           , B(19) => muxInB_1_19_port, B(18) => 
                           muxInB_1_18_port, B(17) => muxInB_1_17_port, B(16) 
                           => muxInB_1_16_port, B(15) => muxInB_1_15_port, 
                           B(14) => muxInB_1_14_port, B(13) => muxInB_1_13_port
                           , B(12) => muxInB_1_12_port, B(11) => 
                           muxInB_1_11_port, B(10) => muxInB_1_10_port, B(9) =>
                           muxInB_1_9_port, B(8) => muxInB_1_8_port, B(7) => 
                           muxInB_1_7_port, B(6) => muxInB_1_6_port, B(5) => 
                           muxInB_1_5_port, B(4) => muxInB_1_4_port, B(3) => 
                           muxInB_1_3_port, B(2) => muxInB_1_2_port, B(1) => 
                           net60063, B(0) => net60064, C(31) => 
                           muxInC_1_31_port, C(30) => muxInC_1_30_port, C(29) 
                           => muxInC_1_29_port, C(28) => muxInC_1_28_port, 
                           C(27) => muxInC_1_27_port, C(26) => muxInC_1_26_port
                           , C(25) => muxInC_1_25_port, C(24) => 
                           muxInC_1_24_port, C(23) => muxInC_1_23_port, C(22) 
                           => muxInC_1_22_port, C(21) => muxInC_1_21_port, 
                           C(20) => muxInC_1_20_port, C(19) => net51440, C(18) 
                           => muxInC_1_18_port, C(17) => muxInC_1_17_port, 
                           C(16) => muxInC_1_16_port, C(15) => muxInC_1_15_port
                           , C(14) => muxInC_1_14_port, C(13) => 
                           muxInC_1_13_port, C(12) => muxInC_1_12_port, C(11) 
                           => muxInC_1_11_port, C(10) => muxInC_1_10_port, C(9)
                           => muxInC_1_9_port, C(8) => muxInC_1_8_port, C(7) =>
                           muxInC_1_7_port, C(6) => muxInC_1_6_port, C(5) => 
                           muxInC_1_5_port, C(4) => muxInC_1_4_port, C(3) => 
                           muxInC_1_3_port, C(2) => muxInC_1_2_port, C(1) => 
                           net60065, C(0) => net60066, D(31) => 
                           muxInD_1_31_port, D(30) => muxInD_1_30_port, D(29) 
                           => muxInD_1_29_port, D(28) => muxInD_1_28_port, 
                           D(27) => muxInD_1_27_port, D(26) => muxInD_1_26_port
                           , D(25) => muxInD_1_25_port, D(24) => 
                           muxInD_1_24_port, D(23) => muxInD_1_23_port, D(22) 
                           => muxInD_1_22_port, D(21) => muxInD_1_21_port, 
                           D(20) => muxInD_1_20_port, D(19) => muxInD_1_19_port
                           , D(18) => muxInD_1_18_port, D(17) => 
                           muxInD_1_17_port, D(16) => muxInD_1_16_port, D(15) 
                           => muxInD_1_15_port, D(14) => muxInD_1_14_port, 
                           D(13) => muxInD_1_13_port, D(12) => muxInD_1_12_port
                           , D(11) => muxInD_1_11_port, D(10) => 
                           muxInD_1_10_port, D(9) => muxInD_1_9_port, D(8) => 
                           muxInD_1_8_port, D(7) => muxInD_1_7_port, D(6) => 
                           muxInD_1_6_port, D(5) => muxInD_1_5_port, D(4) => 
                           muxInD_1_4_port, D(3) => muxInD_1_3_port, D(2) => 
                           net60067, D(1) => net60068, D(0) => net60069, E(31) 
                           => muxInE_1_31_port, E(30) => muxInE_1_30_port, 
                           E(29) => muxInE_1_29_port, E(28) => muxInE_1_28_port
                           , E(27) => muxInE_1_27_port, E(26) => 
                           muxInE_1_26_port, E(25) => muxInE_1_25_port, E(24) 
                           => muxInE_1_24_port, E(23) => muxInE_1_23_port, 
                           E(22) => muxInE_1_22_port, E(21) => muxInE_1_21_port
                           , E(20) => muxInE_1_20_port, E(19) => 
                           muxInE_1_19_port, E(18) => muxInE_1_18_port, E(17) 
                           => muxInE_1_17_port, E(16) => muxInE_1_16_port, 
                           E(15) => muxInE_1_15_port, E(14) => muxInE_1_14_port
                           , E(13) => muxInE_1_13_port, E(12) => 
                           muxInE_1_12_port, E(11) => muxInE_1_11_port, E(10) 
                           => muxInE_1_10_port, E(9) => muxInE_1_9_port, E(8) 
                           => muxInE_1_8_port, E(7) => muxInE_1_7_port, E(6) =>
                           muxInE_1_6_port, E(5) => muxInE_1_5_port, E(4) => 
                           muxInE_1_4_port, E(3) => muxInE_1_3_port, E(2) => 
                           net60070, E(1) => net60071, E(0) => net60072);
   SHIFTERS_2 : shift_mul_N16_S4 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_2_31_port, B(30)
                           => muxInB_2_30_port, B(29) => muxInB_2_29_port, 
                           B(28) => muxInB_2_28_port, B(27) => muxInB_2_27_port
                           , B(26) => muxInB_2_26_port, B(25) => 
                           muxInB_2_25_port, B(24) => muxInB_2_24_port, B(23) 
                           => muxInB_2_23_port, B(22) => muxInB_2_22_port, 
                           B(21) => muxInB_2_21_port, B(20) => muxInB_2_20_port
                           , B(19) => muxInB_2_19_port, B(18) => 
                           muxInB_2_18_port, B(17) => muxInB_2_17_port, B(16) 
                           => muxInB_2_16_port, B(15) => muxInB_2_15_port, 
                           B(14) => muxInB_2_14_port, B(13) => muxInB_2_13_port
                           , B(12) => muxInB_2_12_port, B(11) => 
                           muxInB_2_11_port, B(10) => muxInB_2_10_port, B(9) =>
                           muxInB_2_9_port, B(8) => muxInB_2_8_port, B(7) => 
                           muxInB_2_7_port, B(6) => muxInB_2_6_port, B(5) => 
                           muxInB_2_5_port, B(4) => muxInB_2_4_port, B(3) => 
                           net60045, B(2) => net60046, B(1) => net60047, B(0) 
                           => net60048, C(31) => muxInC_2_31_port, C(30) => 
                           muxInC_2_30_port, C(29) => muxInC_2_29_port, C(28) 
                           => muxInC_2_28_port, C(27) => muxInC_2_27_port, 
                           C(26) => muxInC_2_26_port, C(25) => muxInC_2_25_port
                           , C(24) => muxInC_2_24_port, C(23) => 
                           muxInC_2_23_port, C(22) => muxInC_2_22_port, C(21) 
                           => muxInC_2_21_port, C(20) => muxInC_2_20_port, 
                           C(19) => muxInC_2_19_port, C(18) => muxInC_2_18_port
                           , C(17) => muxInC_2_17_port, C(16) => 
                           muxInC_2_16_port, C(15) => muxInC_2_15_port, C(14) 
                           => muxInC_2_14_port, C(13) => muxInC_2_13_port, 
                           C(12) => muxInC_2_12_port, C(11) => muxInC_2_11_port
                           , C(10) => muxInC_2_10_port, C(9) => muxInC_2_9_port
                           , C(8) => muxInC_2_8_port, C(7) => muxInC_2_7_port, 
                           C(6) => muxInC_2_6_port, C(5) => muxInC_2_5_port, 
                           C(4) => muxInC_2_4_port, C(3) => net60049, C(2) => 
                           net60050, C(1) => net60051, C(0) => net60052, D(31) 
                           => muxInD_2_31_port, D(30) => muxInD_2_30_port, 
                           D(29) => muxInD_2_29_port, D(28) => muxInD_2_28_port
                           , D(27) => muxInD_2_27_port, D(26) => 
                           muxInD_2_26_port, D(25) => muxInD_2_25_port, D(24) 
                           => muxInD_2_24_port, D(23) => muxInD_2_23_port, 
                           D(22) => muxInD_2_22_port, D(21) => muxInD_2_21_port
                           , D(20) => muxInD_2_20_port, D(19) => 
                           muxInD_2_19_port, D(18) => muxInD_2_18_port, D(17) 
                           => muxInD_2_17_port, D(16) => muxInD_2_16_port, 
                           D(15) => muxInD_2_15_port, D(14) => muxInD_2_14_port
                           , D(13) => muxInD_2_13_port, D(12) => 
                           muxInD_2_12_port, D(11) => muxInD_2_11_port, D(10) 
                           => muxInD_2_10_port, D(9) => muxInD_2_9_port, D(8) 
                           => muxInD_2_8_port, D(7) => muxInD_2_7_port, D(6) =>
                           muxInD_2_6_port, D(5) => muxInD_2_5_port, D(4) => 
                           net60053, D(3) => net60054, D(2) => net60055, D(1) 
                           => net60056, D(0) => net60057, E(31) => 
                           muxInE_2_31_port, E(30) => muxInE_2_30_port, E(29) 
                           => muxInE_2_29_port, E(28) => muxInE_2_28_port, 
                           E(27) => muxInE_2_27_port, E(26) => muxInE_2_26_port
                           , E(25) => muxInE_2_25_port, E(24) => 
                           muxInE_2_24_port, E(23) => muxInE_2_23_port, E(22) 
                           => muxInE_2_22_port, E(21) => muxInE_2_21_port, 
                           E(20) => n20, E(19) => muxInE_2_19_port, E(18) => 
                           muxInE_2_18_port, E(17) => muxInE_2_17_port, E(16) 
                           => muxInE_2_16_port, E(15) => muxInE_2_15_port, 
                           E(14) => muxInE_2_14_port, E(13) => muxInE_2_13_port
                           , E(12) => muxInE_2_12_port, E(11) => 
                           muxInE_2_11_port, E(10) => muxInE_2_10_port, E(9) =>
                           muxInE_2_9_port, E(8) => muxInE_2_8_port, E(7) => 
                           muxInE_2_7_port, E(6) => muxInE_2_6_port, E(5) => 
                           muxInE_2_5_port, E(4) => net60058, E(3) => net60059,
                           E(2) => net60060, E(1) => net60061, E(0) => net60062
                           );
   SHIFTERS_3 : shift_mul_N16_S6 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n3, B(31) => muxInB_3_31_port, B(30)
                           => muxInB_3_30_port, B(29) => muxInB_3_29_port, 
                           B(28) => muxInB_3_28_port, B(27) => muxInB_3_27_port
                           , B(26) => muxInB_3_26_port, B(25) => 
                           muxInB_3_25_port, B(24) => muxInB_3_24_port, B(23) 
                           => muxInB_3_23_port, B(22) => muxInB_3_22_port, 
                           B(21) => muxInB_3_21_port, B(20) => muxInB_3_20_port
                           , B(19) => muxInB_3_19_port, B(18) => 
                           muxInB_3_18_port, B(17) => muxInB_3_17_port, B(16) 
                           => muxInB_3_16_port, B(15) => muxInB_3_15_port, 
                           B(14) => muxInB_3_14_port, B(13) => muxInB_3_13_port
                           , B(12) => muxInB_3_12_port, B(11) => 
                           muxInB_3_11_port, B(10) => muxInB_3_10_port, B(9) =>
                           muxInB_3_9_port, B(8) => muxInB_3_8_port, B(7) => 
                           muxInB_3_7_port, B(6) => muxInB_3_6_port, B(5) => 
                           net60019, B(4) => net60020, B(3) => net60021, B(2) 
                           => net60022, B(1) => net60023, B(0) => net60024, 
                           C(31) => muxInC_3_31_port, C(30) => muxInC_3_30_port
                           , C(29) => muxInC_3_29_port, C(28) => 
                           muxInC_3_28_port, C(27) => muxInC_3_27_port, C(26) 
                           => muxInC_3_26_port, C(25) => muxInC_3_25_port, 
                           C(24) => muxInC_3_24_port, C(23) => muxInC_3_23_port
                           , C(22) => muxInC_3_22_port, C(21) => 
                           muxInC_3_21_port, C(20) => muxInC_3_20_port, C(19) 
                           => muxInC_3_19_port, C(18) => muxInC_3_18_port, 
                           C(17) => muxInC_3_17_port, C(16) => muxInC_3_16_port
                           , C(15) => muxInC_3_15_port, C(14) => 
                           muxInC_3_14_port, C(13) => muxInC_3_13_port, C(12) 
                           => muxInC_3_12_port, C(11) => muxInC_3_11_port, 
                           C(10) => muxInC_3_10_port, C(9) => muxInC_3_9_port, 
                           C(8) => muxInC_3_8_port, C(7) => muxInC_3_7_port, 
                           C(6) => muxInC_3_6_port, C(5) => net60025, C(4) => 
                           net60026, C(3) => net60027, C(2) => net60028, C(1) 
                           => net60029, C(0) => net60030, D(31) => 
                           muxInD_3_31_port, D(30) => muxInD_3_30_port, D(29) 
                           => muxInD_3_29_port, D(28) => muxInD_3_28_port, 
                           D(27) => muxInD_3_27_port, D(26) => muxInD_3_26_port
                           , D(25) => muxInD_3_25_port, D(24) => 
                           muxInD_3_24_port, D(23) => muxInD_3_23_port, D(22) 
                           => muxInD_3_22_port, D(21) => muxInD_3_21_port, 
                           D(20) => muxInD_3_20_port, D(19) => muxInD_3_19_port
                           , D(18) => muxInD_3_18_port, D(17) => 
                           muxInD_3_17_port, D(16) => muxInD_3_16_port, D(15) 
                           => muxInD_3_15_port, D(14) => muxInD_3_14_port, 
                           D(13) => muxInD_3_13_port, D(12) => muxInD_3_12_port
                           , D(11) => muxInD_3_11_port, D(10) => 
                           muxInD_3_10_port, D(9) => muxInD_3_9_port, D(8) => 
                           muxInD_3_8_port, D(7) => muxInD_3_7_port, D(6) => 
                           net60031, D(5) => net60032, D(4) => net60033, D(3) 
                           => net60034, D(2) => net60035, D(1) => net60036, 
                           D(0) => net60037, E(31) => muxInE_3_31_port, E(30) 
                           => muxInE_3_30_port, E(29) => muxInE_3_29_port, 
                           E(28) => muxInE_3_28_port, E(27) => muxInE_3_27_port
                           , E(26) => muxInE_3_26_port, E(25) => 
                           muxInE_3_25_port, E(24) => muxInE_3_24_port, E(23) 
                           => muxInE_3_23_port, E(22) => muxInE_3_22_port, 
                           E(21) => muxInE_3_21_port, E(20) => muxInE_3_20_port
                           , E(19) => muxInE_3_19_port, E(18) => 
                           muxInE_3_18_port, E(17) => muxInE_3_17_port, E(16) 
                           => muxInE_3_16_port, E(15) => muxInE_3_15_port, 
                           E(14) => muxInE_3_14_port, E(13) => muxInE_3_13_port
                           , E(12) => muxInE_3_12_port, E(11) => 
                           muxInE_3_11_port, E(10) => muxInE_3_10_port, E(9) =>
                           muxInE_3_9_port, E(8) => muxInE_3_8_port, E(7) => 
                           muxInE_3_7_port, E(6) => net60038, E(5) => net60039,
                           E(4) => net60040, E(3) => net60041, E(2) => net60042
                           , E(1) => net60043, E(0) => net60044);
   SHIFTERS_4 : shift_mul_N16_S8 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_4_31_port, B(30)
                           => muxInB_4_30_port, B(29) => muxInB_4_29_port, 
                           B(28) => muxInB_4_28_port, B(27) => muxInB_4_27_port
                           , B(26) => muxInB_4_26_port, B(25) => 
                           muxInB_4_25_port, B(24) => muxInB_4_24_port, B(23) 
                           => muxInB_4_23_port, B(22) => muxInB_4_22_port, 
                           B(21) => muxInB_4_21_port, B(20) => muxInB_4_20_port
                           , B(19) => muxInB_4_19_port, B(18) => 
                           muxInB_4_18_port, B(17) => muxInB_4_17_port, B(16) 
                           => muxInB_4_16_port, B(15) => muxInB_4_15_port, 
                           B(14) => muxInB_4_14_port, B(13) => muxInB_4_13_port
                           , B(12) => muxInB_4_12_port, B(11) => 
                           muxInB_4_11_port, B(10) => muxInB_4_10_port, B(9) =>
                           muxInB_4_9_port, B(8) => muxInB_4_8_port, B(7) => 
                           net59985, B(6) => net59986, B(5) => net59987, B(4) 
                           => net59988, B(3) => net59989, B(2) => net59990, 
                           B(1) => net59991, B(0) => net59992, C(31) => 
                           muxInC_4_31_port, C(30) => muxInC_4_30_port, C(29) 
                           => muxInC_4_29_port, C(28) => muxInC_4_28_port, 
                           C(27) => muxInC_4_27_port, C(26) => muxInC_4_26_port
                           , C(25) => muxInC_4_25_port, C(24) => 
                           muxInC_4_24_port, C(23) => muxInC_4_23_port, C(22) 
                           => muxInC_4_22_port, C(21) => muxInC_4_21_port, 
                           C(20) => muxInC_4_20_port, C(19) => muxInC_4_19_port
                           , C(18) => muxInC_4_18_port, C(17) => 
                           muxInC_4_17_port, C(16) => muxInC_4_16_port, C(15) 
                           => muxInC_4_15_port, C(14) => muxInC_4_14_port, 
                           C(13) => muxInC_4_13_port, C(12) => muxInC_4_12_port
                           , C(11) => muxInC_4_11_port, C(10) => 
                           muxInC_4_10_port, C(9) => muxInC_4_9_port, C(8) => 
                           muxInC_4_8_port, C(7) => net59993, C(6) => net59994,
                           C(5) => net59995, C(4) => net59996, C(3) => net59997
                           , C(2) => net59998, C(1) => net59999, C(0) => 
                           net60000, D(31) => muxInD_4_31_port, D(30) => 
                           muxInD_4_30_port, D(29) => muxInD_4_29_port, D(28) 
                           => muxInD_4_28_port, D(27) => muxInD_4_27_port, 
                           D(26) => muxInD_4_26_port, D(25) => muxInD_4_25_port
                           , D(24) => muxInD_4_24_port, D(23) => 
                           muxInD_4_23_port, D(22) => muxInD_4_22_port, D(21) 
                           => muxInD_4_21_port, D(20) => muxInD_4_20_port, 
                           D(19) => muxInD_4_19_port, D(18) => muxInD_4_18_port
                           , D(17) => muxInD_4_17_port, D(16) => 
                           muxInD_4_16_port, D(15) => muxInD_4_15_port, D(14) 
                           => muxInD_4_14_port, D(13) => muxInD_4_13_port, 
                           D(12) => muxInD_4_12_port, D(11) => muxInD_4_11_port
                           , D(10) => muxInD_4_10_port, D(9) => muxInD_4_9_port
                           , D(8) => net60001, D(7) => net60002, D(6) => 
                           net60003, D(5) => net60004, D(4) => net60005, D(3) 
                           => net60006, D(2) => net60007, D(1) => net60008, 
                           D(0) => net60009, E(31) => muxInE_4_31_port, E(30) 
                           => muxInE_4_30_port, E(29) => muxInE_4_29_port, 
                           E(28) => muxInE_4_28_port, E(27) => muxInE_4_27_port
                           , E(26) => muxInE_4_26_port, E(25) => 
                           muxInE_4_25_port, E(24) => muxInE_4_24_port, E(23) 
                           => muxInE_4_23_port, E(22) => muxInE_4_22_port, 
                           E(21) => muxInE_4_21_port, E(20) => muxInE_4_20_port
                           , E(19) => muxInE_4_19_port, E(18) => 
                           muxInE_4_18_port, E(17) => muxInE_4_17_port, E(16) 
                           => muxInE_4_16_port, E(15) => muxInE_4_15_port, 
                           E(14) => muxInE_4_14_port, E(13) => muxInE_4_13_port
                           , E(12) => muxInE_4_12_port, E(11) => 
                           muxInE_4_11_port, E(10) => muxInE_4_10_port, E(9) =>
                           muxInE_4_9_port, E(8) => net60010, E(7) => net60011,
                           E(6) => net60012, E(5) => net60013, E(4) => net60014
                           , E(3) => net60015, E(2) => net60016, E(1) => 
                           net60017, E(0) => net60018);
   SHIFTERS_5 : shift_mul_N16_S10 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n3, B(31) => muxInB_5_31_port, 
                           B(30) => muxInB_5_30_port, B(29) => muxInB_5_29_port
                           , B(28) => muxInB_5_28_port, B(27) => 
                           muxInB_5_27_port, B(26) => muxInB_5_26_port, B(25) 
                           => muxInB_5_25_port, B(24) => muxInB_5_24_port, 
                           B(23) => muxInB_5_23_port, B(22) => muxInB_5_22_port
                           , B(21) => muxInB_5_21_port, B(20) => 
                           muxInB_5_20_port, B(19) => muxInB_5_19_port, B(18) 
                           => muxInB_5_18_port, B(17) => muxInB_5_17_port, 
                           B(16) => muxInB_5_16_port, B(15) => muxInB_5_15_port
                           , B(14) => muxInB_5_14_port, B(13) => 
                           muxInB_5_13_port, B(12) => muxInB_5_12_port, B(11) 
                           => muxInB_5_11_port, B(10) => muxInB_5_10_port, B(9)
                           => net59943, B(8) => net59944, B(7) => net59945, 
                           B(6) => net59946, B(5) => net59947, B(4) => net59948
                           , B(3) => net59949, B(2) => net59950, B(1) => 
                           net59951, B(0) => net59952, C(31) => 
                           muxInC_5_31_port, C(30) => muxInC_5_30_port, C(29) 
                           => muxInC_5_29_port, C(28) => muxInC_5_28_port, 
                           C(27) => muxInC_5_27_port, C(26) => muxInC_5_26_port
                           , C(25) => muxInC_5_25_port, C(24) => 
                           muxInC_5_24_port, C(23) => muxInC_5_23_port, C(22) 
                           => muxInC_5_22_port, C(21) => muxInC_5_21_port, 
                           C(20) => muxInC_5_20_port, C(19) => muxInC_5_19_port
                           , C(18) => muxInC_5_18_port, C(17) => 
                           muxInC_5_17_port, C(16) => muxInC_5_16_port, C(15) 
                           => muxInC_5_15_port, C(14) => muxInC_5_14_port, 
                           C(13) => muxInC_5_13_port, C(12) => muxInC_5_12_port
                           , C(11) => muxInC_5_11_port, C(10) => 
                           muxInC_5_10_port, C(9) => net59953, C(8) => net59954
                           , C(7) => net59955, C(6) => net59956, C(5) => 
                           net59957, C(4) => net59958, C(3) => net59959, C(2) 
                           => net59960, C(1) => net59961, C(0) => net59962, 
                           D(31) => muxInD_5_31_port, D(30) => muxInD_5_30_port
                           , D(29) => muxInD_5_29_port, D(28) => 
                           muxInD_5_28_port, D(27) => muxInD_5_27_port, D(26) 
                           => muxInD_5_26_port, D(25) => muxInD_5_25_port, 
                           D(24) => muxInD_5_24_port, D(23) => muxInD_5_23_port
                           , D(22) => muxInD_5_22_port, D(21) => 
                           muxInD_5_21_port, D(20) => muxInD_5_20_port, D(19) 
                           => muxInD_5_19_port, D(18) => muxInD_5_18_port, 
                           D(17) => muxInD_5_17_port, D(16) => muxInD_5_16_port
                           , D(15) => muxInD_5_15_port, D(14) => 
                           muxInD_5_14_port, D(13) => muxInD_5_13_port, D(12) 
                           => muxInD_5_12_port, D(11) => muxInD_5_11_port, 
                           D(10) => net59963, D(9) => net59964, D(8) => 
                           net59965, D(7) => net59966, D(6) => net59967, D(5) 
                           => net59968, D(4) => net59969, D(3) => net59970, 
                           D(2) => net59971, D(1) => net59972, D(0) => net59973
                           , E(31) => muxInE_5_31_port, E(30) => 
                           muxInE_5_30_port, E(29) => muxInE_5_29_port, E(28) 
                           => muxInE_5_28_port, E(27) => muxInE_5_27_port, 
                           E(26) => muxInE_5_26_port, E(25) => muxInE_5_25_port
                           , E(24) => muxInE_5_24_port, E(23) => 
                           muxInE_5_23_port, E(22) => muxInE_5_22_port, E(21) 
                           => muxInE_5_21_port, E(20) => muxInE_5_20_port, 
                           E(19) => muxInE_5_19_port, E(18) => muxInE_5_18_port
                           , E(17) => muxInE_5_17_port, E(16) => 
                           muxInE_5_16_port, E(15) => muxInE_5_15_port, E(14) 
                           => muxInE_5_14_port, E(13) => muxInE_5_13_port, 
                           E(12) => muxInE_5_12_port, E(11) => muxInE_5_11_port
                           , E(10) => net59974, E(9) => net59975, E(8) => 
                           net59976, E(7) => net59977, E(6) => net59978, E(5) 
                           => net59979, E(4) => net59980, E(3) => net59981, 
                           E(2) => net59982, E(1) => net59983, E(0) => net59984
                           );
   SHIFTERS_6 : shift_mul_N16_S12 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n3, B(31) => muxInB_6_31_port, 
                           B(30) => muxInB_6_30_port, B(29) => muxInB_6_29_port
                           , B(28) => muxInB_6_28_port, B(27) => 
                           muxInB_6_27_port, B(26) => muxInB_6_26_port, B(25) 
                           => muxInB_6_25_port, B(24) => muxInB_6_24_port, 
                           B(23) => muxInB_6_23_port, B(22) => muxInB_6_22_port
                           , B(21) => muxInB_6_21_port, B(20) => 
                           muxInB_6_20_port, B(19) => muxInB_6_19_port, B(18) 
                           => muxInB_6_18_port, B(17) => muxInB_6_17_port, 
                           B(16) => muxInB_6_16_port, B(15) => muxInB_6_15_port
                           , B(14) => muxInB_6_14_port, B(13) => 
                           muxInB_6_13_port, B(12) => muxInB_6_12_port, B(11) 
                           => net59893, B(10) => net59894, B(9) => net59895, 
                           B(8) => net59896, B(7) => net59897, B(6) => net59898
                           , B(5) => net59899, B(4) => net59900, B(3) => 
                           net59901, B(2) => net59902, B(1) => net59903, B(0) 
                           => net59904, C(31) => muxInC_6_31_port, C(30) => 
                           muxInC_6_30_port, C(29) => muxInC_6_29_port, C(28) 
                           => muxInC_6_28_port, C(27) => muxInC_6_27_port, 
                           C(26) => muxInC_6_26_port, C(25) => muxInC_6_25_port
                           , C(24) => muxInC_6_24_port, C(23) => 
                           muxInC_6_23_port, C(22) => muxInC_6_22_port, C(21) 
                           => muxInC_6_21_port, C(20) => muxInC_6_20_port, 
                           C(19) => muxInC_6_19_port, C(18) => muxInC_6_18_port
                           , C(17) => muxInC_6_17_port, C(16) => 
                           muxInC_6_16_port, C(15) => muxInC_6_15_port, C(14) 
                           => muxInC_6_14_port, C(13) => muxInC_6_13_port, 
                           C(12) => muxInC_6_12_port, C(11) => net59905, C(10) 
                           => net59906, C(9) => net59907, C(8) => net59908, 
                           C(7) => net59909, C(6) => net59910, C(5) => net59911
                           , C(4) => net59912, C(3) => net59913, C(2) => 
                           net59914, C(1) => net59915, C(0) => net59916, D(31) 
                           => muxInD_6_31_port, D(30) => muxInD_6_30_port, 
                           D(29) => muxInD_6_29_port, D(28) => muxInD_6_28_port
                           , D(27) => muxInD_6_27_port, D(26) => 
                           muxInD_6_26_port, D(25) => muxInD_6_25_port, D(24) 
                           => muxInD_6_24_port, D(23) => muxInD_6_23_port, 
                           D(22) => muxInD_6_22_port, D(21) => muxInD_6_21_port
                           , D(20) => muxInD_6_20_port, D(19) => 
                           muxInD_6_19_port, D(18) => muxInD_6_18_port, D(17) 
                           => muxInD_6_17_port, D(16) => muxInD_6_16_port, 
                           D(15) => muxInD_6_15_port, D(14) => muxInD_6_14_port
                           , D(13) => muxInD_6_13_port, D(12) => net59917, 
                           D(11) => net59918, D(10) => net59919, D(9) => 
                           net59920, D(8) => net59921, D(7) => net59922, D(6) 
                           => net59923, D(5) => net59924, D(4) => net59925, 
                           D(3) => net59926, D(2) => net59927, D(1) => net59928
                           , D(0) => net59929, E(31) => muxInE_6_31_port, E(30)
                           => muxInE_6_30_port, E(29) => muxInE_6_29_port, 
                           E(28) => muxInE_6_28_port, E(27) => muxInE_6_27_port
                           , E(26) => muxInE_6_26_port, E(25) => 
                           muxInE_6_25_port, E(24) => muxInE_6_24_port, E(23) 
                           => muxInE_6_23_port, E(22) => muxInE_6_22_port, 
                           E(21) => muxInE_6_21_port, E(20) => muxInE_6_20_port
                           , E(19) => muxInE_6_19_port, E(18) => 
                           muxInE_6_18_port, E(17) => muxInE_6_17_port, E(16) 
                           => muxInE_6_16_port, E(15) => muxInE_6_15_port, 
                           E(14) => muxInE_6_14_port, E(13) => muxInE_6_13_port
                           , E(12) => net59930, E(11) => net59931, E(10) => 
                           net59932, E(9) => net59933, E(8) => net59934, E(7) 
                           => net59935, E(6) => net59936, E(5) => net59937, 
                           E(4) => net59938, E(3) => net59939, E(2) => net59940
                           , E(1) => net59941, E(0) => net59942);
   SHIFTERS_7 : shift_mul_N16_S14 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n2, B(31) => muxInB_7_31_port, 
                           B(30) => muxInB_7_30_port, B(29) => muxInB_7_29_port
                           , B(28) => muxInB_7_28_port, B(27) => 
                           muxInB_7_27_port, B(26) => muxInB_7_26_port, B(25) 
                           => muxInB_7_25_port, B(24) => muxInB_7_24_port, 
                           B(23) => muxInB_7_23_port, B(22) => muxInB_7_22_port
                           , B(21) => muxInB_7_21_port, B(20) => 
                           muxInB_7_20_port, B(19) => muxInB_7_19_port, B(18) 
                           => muxInB_7_18_port, B(17) => muxInB_7_17_port, 
                           B(16) => muxInB_7_16_port, B(15) => muxInB_7_15_port
                           , B(14) => muxInB_7_14_port, B(13) => net59835, 
                           B(12) => net59836, B(11) => net59837, B(10) => 
                           net59838, B(9) => net59839, B(8) => net59840, B(7) 
                           => net59841, B(6) => net59842, B(5) => net59843, 
                           B(4) => net59844, B(3) => net59845, B(2) => net59846
                           , B(1) => net59847, B(0) => net59848, C(31) => 
                           muxInC_7_31_port, C(30) => muxInC_7_30_port, C(29) 
                           => muxInC_7_29_port, C(28) => muxInC_7_28_port, 
                           C(27) => muxInC_7_27_port, C(26) => muxInC_7_26_port
                           , C(25) => muxInC_7_25_port, C(24) => 
                           muxInC_7_24_port, C(23) => muxInC_7_23_port, C(22) 
                           => muxInC_7_22_port, C(21) => muxInC_7_21_port, 
                           C(20) => muxInC_7_20_port, C(19) => muxInC_7_19_port
                           , C(18) => muxInC_7_18_port, C(17) => 
                           muxInC_7_17_port, C(16) => muxInC_7_16_port, C(15) 
                           => muxInC_7_15_port, C(14) => muxInC_7_14_port, 
                           C(13) => net59849, C(12) => net59850, C(11) => 
                           net59851, C(10) => net59852, C(9) => net59853, C(8) 
                           => net59854, C(7) => net59855, C(6) => net59856, 
                           C(5) => net59857, C(4) => net59858, C(3) => net59859
                           , C(2) => net59860, C(1) => net59861, C(0) => 
                           net59862, D(31) => muxInD_7_31_port, D(30) => 
                           muxInD_7_30_port, D(29) => muxInD_7_29_port, D(28) 
                           => muxInD_7_28_port, D(27) => muxInD_7_27_port, 
                           D(26) => muxInD_7_26_port, D(25) => muxInD_7_25_port
                           , D(24) => muxInD_7_24_port, D(23) => 
                           muxInD_7_23_port, D(22) => muxInD_7_22_port, D(21) 
                           => muxInD_7_21_port, D(20) => muxInD_7_20_port, 
                           D(19) => muxInD_7_19_port, D(18) => muxInD_7_18_port
                           , D(17) => muxInD_7_17_port, D(16) => 
                           muxInD_7_16_port, D(15) => muxInD_7_15_port, D(14) 
                           => net59863, D(13) => net59864, D(12) => net59865, 
                           D(11) => net59866, D(10) => net59867, D(9) => 
                           net59868, D(8) => net59869, D(7) => net59870, D(6) 
                           => net59871, D(5) => net59872, D(4) => net59873, 
                           D(3) => net59874, D(2) => net59875, D(1) => net59876
                           , D(0) => net59877, E(31) => muxInE_7_31_port, E(30)
                           => muxInE_7_30_port, E(29) => muxInE_7_29_port, 
                           E(28) => muxInE_7_28_port, E(27) => muxInE_7_27_port
                           , E(26) => muxInE_7_26_port, E(25) => 
                           muxInE_7_25_port, E(24) => muxInE_7_24_port, E(23) 
                           => muxInE_7_23_port, E(22) => muxInE_7_22_port, 
                           E(21) => muxInE_7_21_port, E(20) => muxInE_7_20_port
                           , E(19) => muxInE_7_19_port, E(18) => 
                           muxInE_7_18_port, E(17) => muxInE_7_17_port, E(16) 
                           => muxInE_7_16_port, E(15) => muxInE_7_15_port, 
                           E(14) => net59878, E(13) => net59879, E(12) => 
                           net59880, E(11) => net59881, E(10) => net59882, E(9)
                           => net59883, E(8) => net59884, E(7) => net59885, 
                           E(6) => net59886, E(5) => net59887, E(4) => net59888
                           , E(3) => net59889, E(2) => net59890, E(1) => 
                           net59891, E(0) => net59892);
   MUXGEN_0 : mux_N32_0 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_0_31_port, B(30) => 
                           muxInB_0_30_port, B(29) => muxInB_0_29_port, B(28) 
                           => muxInB_0_28_port, B(27) => muxInB_0_27_port, 
                           B(26) => muxInB_0_26_port, B(25) => muxInB_0_25_port
                           , B(24) => muxInB_0_24_port, B(23) => 
                           muxInB_0_23_port, B(22) => muxInB_0_22_port, B(21) 
                           => muxInB_0_21_port, B(20) => muxInB_0_20_port, 
                           B(19) => muxInB_0_19_port, B(18) => muxInB_0_18_port
                           , B(17) => muxInB_0_17_port, B(16) => 
                           muxInB_0_16_port, B(15) => muxInB_0_15_port, B(14) 
                           => muxInB_0_14_port, B(13) => muxInB_0_13_port, 
                           B(12) => muxInB_0_12_port, B(11) => muxInB_0_11_port
                           , B(10) => muxInB_0_10_port, B(9) => muxInB_0_9_port
                           , B(8) => muxInB_0_8_port, B(7) => muxInB_0_7_port, 
                           B(6) => muxInB_0_6_port, B(5) => muxInB_0_5_port, 
                           B(4) => muxInB_0_4_port, B(3) => muxInB_0_3_port, 
                           B(2) => muxInB_0_2_port, B(1) => muxInB_0_1_port, 
                           B(0) => muxInB_0_0_port, C(31) => muxInC_0_31_port, 
                           C(30) => muxInC_0_30_port, C(29) => muxInC_0_29_port
                           , C(28) => muxInC_0_28_port, C(27) => 
                           muxInC_0_20_port, C(26) => muxInC_0_26_port, C(25) 
                           => muxInC_0_25_port, C(24) => muxInC_0_24_port, 
                           C(23) => muxInC_0_23_port, C(22) => muxInC_0_22_port
                           , C(21) => muxInC_0_21_port, C(20) => 
                           muxInC_0_20_port, C(19) => muxInC_0_19_port, C(18) 
                           => muxInC_0_18_port, C(17) => muxInC_0_17_port, 
                           C(16) => muxInC_0_16_port, C(15) => muxInC_0_15_port
                           , C(14) => muxInC_0_14_port, C(13) => 
                           muxInC_0_13_port, C(12) => muxInC_0_12_port, C(11) 
                           => muxInC_0_11_port, C(10) => muxInC_0_10_port, C(9)
                           => muxInC_0_9_port, C(8) => muxInC_0_8_port, C(7) =>
                           muxInC_0_7_port, C(6) => muxInC_0_6_port, C(5) => 
                           muxInC_0_5_port, C(4) => muxInC_0_4_port, C(3) => 
                           muxInC_0_3_port, C(2) => muxInC_0_2_port, C(1) => 
                           muxInC_0_1_port, C(0) => muxInC_0_0_port, D(31) => 
                           muxInD_0_31_port, D(30) => muxInD_0_30_port, D(29) 
                           => muxInD_0_29_port, D(28) => muxInD_0_28_port, 
                           D(27) => muxInD_0_27_port, D(26) => muxInD_0_26_port
                           , D(25) => muxInD_0_25_port, D(24) => 
                           muxInD_0_24_port, D(23) => muxInD_0_23_port, D(22) 
                           => muxInD_0_22_port, D(21) => muxInD_0_21_port, 
                           D(20) => muxInD_0_20_port, D(19) => muxInD_0_19_port
                           , D(18) => muxInD_0_18_port, D(17) => 
                           muxInD_0_17_port, D(16) => muxInD_0_16_port, D(15) 
                           => muxInD_0_15_port, D(14) => muxInD_0_14_port, 
                           D(13) => muxInD_0_13_port, D(12) => muxInD_0_12_port
                           , D(11) => muxInD_0_11_port, D(10) => 
                           muxInD_0_10_port, D(9) => muxInD_0_9_port, D(8) => 
                           muxInD_0_8_port, D(7) => muxInD_0_7_port, D(6) => 
                           muxInD_0_6_port, D(5) => muxInD_0_5_port, D(4) => 
                           muxInD_0_4_port, D(3) => muxInD_0_3_port, D(2) => 
                           muxInD_0_2_port, D(1) => muxInD_0_1_port, D(0) => 
                           muxInD_0_0_port, E(31) => muxInE_0_31_port, E(30) =>
                           muxInE_0_30_port, E(29) => muxInE_0_29_port, E(28) 
                           => muxInE_0_28_port, E(27) => muxInE_0_27_port, 
                           E(26) => muxInE_0_26_port, E(25) => muxInC_0_20_port
                           , E(24) => muxInE_0_24_port, E(23) => 
                           muxInE_0_23_port, E(22) => muxInC_0_27_port, E(21) 
                           => muxInE_0_21_port, E(20) => muxInE_0_20_port, 
                           E(19) => muxInE_0_19_port, E(18) => muxInE_0_18_port
                           , E(17) => muxInC_0_29_port, E(16) => 
                           muxInE_0_16_port, E(15) => muxInE_0_15_port, E(14) 
                           => muxInE_0_14_port, E(13) => muxInE_0_13_port, 
                           E(12) => muxInE_0_12_port, E(11) => muxInE_0_11_port
                           , E(10) => muxInE_0_10_port, E(9) => muxInE_0_9_port
                           , E(8) => muxInE_0_8_port, E(7) => muxInE_0_7_port, 
                           E(6) => muxInE_0_6_port, E(5) => muxInE_0_5_port, 
                           E(4) => muxInE_0_4_port, E(3) => muxInE_0_3_port, 
                           E(2) => muxInE_0_2_port, E(1) => muxInE_0_1_port, 
                           E(0) => muxInE_0_0_port, Sel(2) => B(1), Sel(1) => 
                           B(0), Sel(0) => X_Logic0_port, O(31) => 
                           outmux_0_31_port, O(30) => outmux_0_30_port, O(29) 
                           => outmux_0_29_port, O(28) => outmux_0_28_port, 
                           O(27) => outmux_0_27_port, O(26) => outmux_0_26_port
                           , O(25) => outmux_0_25_port, O(24) => 
                           outmux_0_24_port, O(23) => outmux_0_23_port, O(22) 
                           => outmux_0_22_port, O(21) => outmux_0_21_port, 
                           O(20) => outmux_0_20_port, O(19) => outmux_0_19_port
                           , O(18) => outmux_0_18_port, O(17) => 
                           outmux_0_17_port, O(16) => outmux_0_16_port, O(15) 
                           => outmux_0_15_port, O(14) => outmux_0_14_port, 
                           O(13) => outmux_0_13_port, O(12) => outmux_0_12_port
                           , O(11) => outmux_0_11_port, O(10) => 
                           outmux_0_10_port, O(9) => outmux_0_9_port, O(8) => 
                           outmux_0_8_port, O(7) => outmux_0_7_port, O(6) => 
                           outmux_0_6_port, O(5) => outmux_0_5_port, O(4) => 
                           outmux_0_4_port, O(3) => outmux_0_3_port, O(2) => 
                           outmux_0_2_port, O(1) => outmux_0_1_port, O(0) => 
                           outmux_0_0_port);
   MUXGEN_1 : mux_N32_7 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_1_31_port, B(30) => 
                           muxInB_1_30_port, B(29) => muxInB_1_29_port, B(28) 
                           => muxInB_1_28_port, B(27) => muxInB_1_27_port, 
                           B(26) => muxInB_1_26_port, B(25) => muxInB_1_25_port
                           , B(24) => muxInB_1_24_port, B(23) => 
                           muxInB_1_23_port, B(22) => muxInB_1_22_port, B(21) 
                           => muxInB_1_21_port, B(20) => muxInB_1_20_port, 
                           B(19) => muxInB_1_19_port, B(18) => muxInB_1_18_port
                           , B(17) => muxInB_1_17_port, B(16) => 
                           muxInB_1_16_port, B(15) => muxInB_1_15_port, B(14) 
                           => muxInB_1_14_port, B(13) => muxInB_1_13_port, 
                           B(12) => muxInB_1_12_port, B(11) => muxInB_1_11_port
                           , B(10) => muxInB_1_10_port, B(9) => muxInB_1_9_port
                           , B(8) => muxInB_1_8_port, B(7) => muxInB_1_7_port, 
                           B(6) => muxInB_1_6_port, B(5) => muxInB_1_5_port, 
                           B(4) => muxInB_1_4_port, B(3) => muxInB_1_3_port, 
                           B(2) => muxInB_1_2_port, B(1) => muxInB_1_1_port, 
                           B(0) => muxInB_1_0_port, C(31) => muxInC_1_31_port, 
                           C(30) => muxInC_1_30_port, C(29) => muxInC_1_29_port
                           , C(28) => muxInC_1_28_port, C(27) => 
                           muxInC_1_27_port, C(26) => muxInC_1_26_port, C(25) 
                           => muxInC_1_25_port, C(24) => muxInC_1_24_port, 
                           C(23) => muxInE_1_23_port, C(22) => muxInC_1_22_port
                           , C(21) => muxInC_1_21_port, C(20) => 
                           muxInC_1_20_port, C(19) => muxInC_1_23_port, C(18) 
                           => muxInC_1_18_port, C(17) => muxInC_1_17_port, 
                           C(16) => muxInC_1_16_port, C(15) => muxInC_1_15_port
                           , C(14) => muxInC_1_14_port, C(13) => 
                           muxInC_1_13_port, C(12) => muxInC_1_12_port, C(11) 
                           => muxInC_1_11_port, C(10) => muxInC_1_10_port, C(9)
                           => muxInC_1_9_port, C(8) => muxInC_1_8_port, C(7) =>
                           muxInC_1_7_port, C(6) => muxInC_1_6_port, C(5) => 
                           muxInC_1_5_port, C(4) => muxInC_1_4_port, C(3) => 
                           muxInC_1_3_port, C(2) => muxInC_1_2_port, C(1) => 
                           muxInC_1_1_port, C(0) => muxInC_1_0_port, D(31) => 
                           muxInD_1_31_port, D(30) => muxInD_1_30_port, D(29) 
                           => muxInD_1_29_port, D(28) => muxInD_1_28_port, 
                           D(27) => muxInD_1_27_port, D(26) => muxInD_1_26_port
                           , D(25) => muxInD_1_25_port, D(24) => 
                           muxInD_1_24_port, D(23) => muxInD_1_23_port, D(22) 
                           => muxInD_1_22_port, D(21) => muxInD_1_21_port, 
                           D(20) => muxInD_1_20_port, D(19) => muxInD_1_19_port
                           , D(18) => muxInD_1_18_port, D(17) => 
                           muxInD_1_17_port, D(16) => muxInD_1_16_port, D(15) 
                           => muxInD_1_15_port, D(14) => muxInD_1_14_port, 
                           D(13) => muxInD_1_13_port, D(12) => muxInD_1_12_port
                           , D(11) => muxInD_1_11_port, D(10) => 
                           muxInD_1_10_port, D(9) => muxInD_1_9_port, D(8) => 
                           muxInD_1_8_port, D(7) => muxInD_1_7_port, D(6) => 
                           muxInD_1_6_port, D(5) => muxInD_1_5_port, D(4) => 
                           muxInD_1_4_port, D(3) => muxInD_1_3_port, D(2) => 
                           muxInD_1_2_port, D(1) => muxInD_1_1_port, D(0) => 
                           muxInD_1_0_port, E(31) => muxInE_1_31_port, E(30) =>
                           muxInE_1_30_port, E(29) => muxInE_1_29_port, E(28) 
                           => muxInE_1_28_port, E(27) => muxInE_1_27_port, 
                           E(26) => muxInE_1_26_port, E(25) => muxInE_1_25_port
                           , E(24) => muxInE_1_24_port, E(23) => 
                           muxInE_1_23_port, E(22) => muxInE_1_22_port, E(21) 
                           => muxInE_1_21_port, E(20) => muxInE_1_20_port, 
                           E(19) => muxInE_1_19_port, E(18) => muxInE_1_18_port
                           , E(17) => muxInE_1_17_port, E(16) => 
                           muxInE_1_16_port, E(15) => muxInE_1_15_port, E(14) 
                           => muxInE_1_14_port, E(13) => muxInE_1_13_port, 
                           E(12) => muxInE_1_12_port, E(11) => muxInE_1_11_port
                           , E(10) => muxInE_1_10_port, E(9) => muxInE_1_9_port
                           , E(8) => muxInE_1_8_port, E(7) => muxInE_1_7_port, 
                           E(6) => muxInE_1_6_port, E(5) => muxInE_1_5_port, 
                           E(4) => muxInE_1_4_port, E(3) => muxInE_1_3_port, 
                           E(2) => muxInE_1_2_port, E(1) => muxInE_1_1_port, 
                           E(0) => muxInE_1_0_port, Sel(2) => B(3), Sel(1) => 
                           B(2), Sel(0) => B(1), O(31) => outmux_1_31_port, 
                           O(30) => outmux_1_30_port, O(29) => outmux_1_29_port
                           , O(28) => outmux_1_28_port, O(27) => 
                           outmux_1_27_port, O(26) => outmux_1_26_port, O(25) 
                           => outmux_1_25_port, O(24) => outmux_1_24_port, 
                           O(23) => outmux_1_23_port, O(22) => outmux_1_22_port
                           , O(21) => outmux_1_21_port, O(20) => 
                           outmux_1_20_port, O(19) => outmux_1_19_port, O(18) 
                           => outmux_1_18_port, O(17) => outmux_1_17_port, 
                           O(16) => outmux_1_16_port, O(15) => outmux_1_15_port
                           , O(14) => outmux_1_14_port, O(13) => 
                           outmux_1_13_port, O(12) => outmux_1_12_port, O(11) 
                           => outmux_1_11_port, O(10) => outmux_1_10_port, O(9)
                           => outmux_1_9_port, O(8) => outmux_1_8_port, O(7) =>
                           outmux_1_7_port, O(6) => outmux_1_6_port, O(5) => 
                           outmux_1_5_port, O(4) => outmux_1_4_port, O(3) => 
                           outmux_1_3_port, O(2) => outmux_1_2_port, O(1) => 
                           outmux_1_1_port, O(0) => outmux_1_0_port);
   MUXGEN_2 : mux_N32_6 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_2_31_port, B(30) => 
                           muxInB_2_30_port, B(29) => muxInB_2_29_port, B(28) 
                           => muxInB_2_28_port, B(27) => muxInB_2_27_port, 
                           B(26) => muxInB_2_26_port, B(25) => muxInB_2_25_port
                           , B(24) => muxInB_2_24_port, B(23) => 
                           muxInB_2_23_port, B(22) => muxInB_2_22_port, B(21) 
                           => muxInB_2_21_port, B(20) => muxInB_2_20_port, 
                           B(19) => muxInB_2_19_port, B(18) => muxInB_2_18_port
                           , B(17) => muxInB_2_17_port, B(16) => 
                           muxInB_2_16_port, B(15) => muxInB_2_15_port, B(14) 
                           => muxInB_2_14_port, B(13) => muxInB_2_13_port, 
                           B(12) => muxInB_2_12_port, B(11) => muxInB_2_11_port
                           , B(10) => muxInB_2_10_port, B(9) => muxInB_2_9_port
                           , B(8) => muxInB_2_8_port, B(7) => muxInB_2_7_port, 
                           B(6) => muxInB_2_6_port, B(5) => muxInB_2_5_port, 
                           B(4) => muxInB_2_4_port, B(3) => muxInB_2_3_port, 
                           B(2) => muxInB_2_2_port, B(1) => muxInB_2_1_port, 
                           B(0) => muxInB_2_0_port, C(31) => muxInC_2_31_port, 
                           C(30) => muxInC_2_30_port, C(29) => muxInC_2_29_port
                           , C(28) => muxInC_2_28_port, C(27) => 
                           muxInC_2_27_port, C(26) => muxInC_2_26_port, C(25) 
                           => muxInC_2_25_port, C(24) => muxInC_2_24_port, 
                           C(23) => muxInC_2_23_port, C(22) => muxInC_2_22_port
                           , C(21) => muxInC_2_21_port, C(20) => 
                           muxInC_2_20_port, C(19) => n20, C(18) => 
                           muxInC_2_18_port, C(17) => muxInC_2_17_port, C(16) 
                           => muxInC_2_16_port, C(15) => muxInC_2_15_port, 
                           C(14) => muxInC_2_14_port, C(13) => muxInC_2_13_port
                           , C(12) => muxInC_2_12_port, C(11) => 
                           muxInC_2_11_port, C(10) => muxInC_2_10_port, C(9) =>
                           muxInC_2_9_port, C(8) => muxInC_2_8_port, C(7) => 
                           muxInC_2_7_port, C(6) => muxInC_2_6_port, C(5) => 
                           muxInC_2_5_port, C(4) => muxInC_2_4_port, C(3) => 
                           muxInC_2_3_port, C(2) => muxInC_2_2_port, C(1) => 
                           muxInC_2_1_port, C(0) => muxInC_2_0_port, D(31) => 
                           muxInD_2_31_port, D(30) => muxInD_2_30_port, D(29) 
                           => muxInD_2_29_port, D(28) => muxInD_2_28_port, 
                           D(27) => muxInD_2_27_port, D(26) => muxInD_2_26_port
                           , D(25) => muxInD_2_25_port, D(24) => 
                           muxInD_2_24_port, D(23) => muxInD_2_23_port, D(22) 
                           => muxInD_2_22_port, D(21) => muxInD_2_21_port, 
                           D(20) => muxInD_2_20_port, D(19) => muxInD_2_19_port
                           , D(18) => muxInD_2_18_port, D(17) => 
                           muxInD_2_17_port, D(16) => muxInD_2_16_port, D(15) 
                           => muxInD_2_15_port, D(14) => muxInD_2_14_port, 
                           D(13) => muxInD_2_13_port, D(12) => muxInD_2_12_port
                           , D(11) => muxInD_2_11_port, D(10) => 
                           muxInD_2_10_port, D(9) => muxInD_2_9_port, D(8) => 
                           muxInD_2_8_port, D(7) => muxInD_2_7_port, D(6) => 
                           muxInD_2_6_port, D(5) => muxInD_2_5_port, D(4) => 
                           muxInD_2_4_port, D(3) => muxInD_2_3_port, D(2) => 
                           muxInD_2_2_port, D(1) => muxInD_2_1_port, D(0) => 
                           muxInD_2_0_port, E(31) => muxInE_2_31_port, E(30) =>
                           muxInE_2_30_port, E(29) => muxInE_2_29_port, E(28) 
                           => muxInE_2_28_port, E(27) => muxInE_2_27_port, 
                           E(26) => muxInE_2_26_port, E(25) => muxInE_2_25_port
                           , E(24) => muxInE_2_24_port, E(23) => 
                           muxInE_2_23_port, E(22) => muxInE_2_22_port, E(21) 
                           => muxInE_2_21_port, E(20) => muxInC_2_19_port, 
                           E(19) => muxInE_2_19_port, E(18) => muxInE_2_18_port
                           , E(17) => muxInE_2_17_port, E(16) => 
                           muxInE_2_16_port, E(15) => muxInE_2_15_port, E(14) 
                           => muxInE_2_14_port, E(13) => muxInE_2_13_port, 
                           E(12) => muxInE_2_12_port, E(11) => muxInE_2_11_port
                           , E(10) => muxInE_2_10_port, E(9) => muxInE_2_9_port
                           , E(8) => muxInE_2_8_port, E(7) => muxInE_2_7_port, 
                           E(6) => muxInE_2_6_port, E(5) => muxInE_2_5_port, 
                           E(4) => muxInE_2_4_port, E(3) => muxInE_2_3_port, 
                           E(2) => muxInE_2_2_port, E(1) => muxInE_2_1_port, 
                           E(0) => muxInE_2_0_port, Sel(2) => B(5), Sel(1) => 
                           B(4), Sel(0) => B(3), O(31) => outmux_2_31_port, 
                           O(30) => outmux_2_30_port, O(29) => outmux_2_29_port
                           , O(28) => outmux_2_28_port, O(27) => 
                           outmux_2_27_port, O(26) => outmux_2_26_port, O(25) 
                           => outmux_2_25_port, O(24) => outmux_2_24_port, 
                           O(23) => outmux_2_23_port, O(22) => outmux_2_22_port
                           , O(21) => outmux_2_21_port, O(20) => 
                           outmux_2_20_port, O(19) => outmux_2_19_port, O(18) 
                           => outmux_2_18_port, O(17) => outmux_2_17_port, 
                           O(16) => outmux_2_16_port, O(15) => outmux_2_15_port
                           , O(14) => outmux_2_14_port, O(13) => 
                           outmux_2_13_port, O(12) => outmux_2_12_port, O(11) 
                           => outmux_2_11_port, O(10) => outmux_2_10_port, O(9)
                           => outmux_2_9_port, O(8) => outmux_2_8_port, O(7) =>
                           outmux_2_7_port, O(6) => outmux_2_6_port, O(5) => 
                           outmux_2_5_port, O(4) => outmux_2_4_port, O(3) => 
                           outmux_2_3_port, O(2) => outmux_2_2_port, O(1) => 
                           outmux_2_1_port, O(0) => outmux_2_0_port);
   MUXGEN_3 : mux_N32_5 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_3_31_port, B(30) => 
                           muxInB_3_30_port, B(29) => muxInB_3_29_port, B(28) 
                           => muxInB_3_28_port, B(27) => muxInB_3_27_port, 
                           B(26) => muxInB_3_26_port, B(25) => muxInB_3_25_port
                           , B(24) => muxInB_3_24_port, B(23) => 
                           muxInB_3_23_port, B(22) => muxInB_3_22_port, B(21) 
                           => muxInB_3_21_port, B(20) => muxInB_3_20_port, 
                           B(19) => muxInB_3_19_port, B(18) => muxInB_3_18_port
                           , B(17) => muxInB_3_17_port, B(16) => 
                           muxInB_3_16_port, B(15) => muxInB_3_15_port, B(14) 
                           => muxInB_3_14_port, B(13) => muxInB_3_13_port, 
                           B(12) => muxInB_3_12_port, B(11) => muxInB_3_11_port
                           , B(10) => muxInB_3_10_port, B(9) => muxInB_3_9_port
                           , B(8) => muxInB_3_8_port, B(7) => muxInB_3_7_port, 
                           B(6) => muxInB_3_6_port, B(5) => muxInB_3_5_port, 
                           B(4) => muxInB_3_4_port, B(3) => muxInB_3_3_port, 
                           B(2) => muxInB_3_2_port, B(1) => muxInB_3_1_port, 
                           B(0) => muxInB_3_0_port, C(31) => muxInC_3_31_port, 
                           C(30) => muxInC_3_30_port, C(29) => muxInC_3_29_port
                           , C(28) => muxInC_3_28_port, C(27) => 
                           muxInC_3_27_port, C(26) => muxInC_3_26_port, C(25) 
                           => muxInC_3_25_port, C(24) => muxInC_3_24_port, 
                           C(23) => muxInC_3_23_port, C(22) => muxInC_3_22_port
                           , C(21) => muxInC_3_21_port, C(20) => 
                           muxInC_3_20_port, C(19) => muxInC_3_19_port, C(18) 
                           => muxInC_3_18_port, C(17) => muxInC_3_17_port, 
                           C(16) => muxInC_3_16_port, C(15) => muxInC_3_15_port
                           , C(14) => muxInC_3_14_port, C(13) => 
                           muxInC_3_13_port, C(12) => muxInC_3_12_port, C(11) 
                           => muxInC_3_11_port, C(10) => muxInC_3_10_port, C(9)
                           => muxInC_3_9_port, C(8) => muxInC_3_8_port, C(7) =>
                           muxInC_3_7_port, C(6) => muxInC_3_6_port, C(5) => 
                           muxInC_3_5_port, C(4) => muxInC_3_4_port, C(3) => 
                           muxInC_3_3_port, C(2) => muxInC_3_2_port, C(1) => 
                           muxInC_3_1_port, C(0) => muxInC_3_0_port, D(31) => 
                           muxInD_3_31_port, D(30) => muxInD_3_30_port, D(29) 
                           => muxInD_3_29_port, D(28) => muxInD_3_28_port, 
                           D(27) => muxInD_3_27_port, D(26) => muxInD_3_26_port
                           , D(25) => muxInD_3_25_port, D(24) => 
                           muxInD_3_24_port, D(23) => muxInD_3_23_port, D(22) 
                           => muxInD_3_22_port, D(21) => muxInD_3_21_port, 
                           D(20) => muxInD_3_20_port, D(19) => muxInD_3_19_port
                           , D(18) => muxInD_3_18_port, D(17) => 
                           muxInD_3_17_port, D(16) => muxInD_3_16_port, D(15) 
                           => muxInD_3_15_port, D(14) => muxInD_3_14_port, 
                           D(13) => muxInD_3_13_port, D(12) => muxInD_3_12_port
                           , D(11) => muxInD_3_11_port, D(10) => 
                           muxInD_3_10_port, D(9) => muxInD_3_9_port, D(8) => 
                           muxInD_3_8_port, D(7) => muxInD_3_7_port, D(6) => 
                           muxInD_3_6_port, D(5) => muxInD_3_5_port, D(4) => 
                           muxInD_3_4_port, D(3) => muxInD_3_3_port, D(2) => 
                           muxInD_3_2_port, D(1) => muxInD_3_1_port, D(0) => 
                           muxInD_3_0_port, E(31) => muxInE_3_31_port, E(30) =>
                           muxInE_3_30_port, E(29) => muxInE_3_29_port, E(28) 
                           => muxInE_3_28_port, E(27) => muxInE_3_27_port, 
                           E(26) => muxInE_3_26_port, E(25) => muxInE_3_25_port
                           , E(24) => muxInE_3_24_port, E(23) => 
                           muxInE_3_23_port, E(22) => muxInE_3_22_port, E(21) 
                           => muxInE_3_21_port, E(20) => muxInE_3_20_port, 
                           E(19) => muxInE_3_19_port, E(18) => muxInE_3_18_port
                           , E(17) => muxInE_3_17_port, E(16) => 
                           muxInE_3_16_port, E(15) => muxInE_3_15_port, E(14) 
                           => muxInE_3_14_port, E(13) => muxInE_3_13_port, 
                           E(12) => muxInE_3_12_port, E(11) => muxInE_3_11_port
                           , E(10) => muxInE_3_10_port, E(9) => muxInE_3_9_port
                           , E(8) => muxInE_3_8_port, E(7) => muxInE_3_7_port, 
                           E(6) => muxInE_3_6_port, E(5) => muxInE_3_5_port, 
                           E(4) => muxInE_3_4_port, E(3) => muxInE_3_3_port, 
                           E(2) => muxInE_3_2_port, E(1) => muxInE_3_1_port, 
                           E(0) => muxInE_3_0_port, Sel(2) => B(7), Sel(1) => 
                           B(6), Sel(0) => B(5), O(31) => outmux_3_31_port, 
                           O(30) => outmux_3_30_port, O(29) => outmux_3_29_port
                           , O(28) => outmux_3_28_port, O(27) => 
                           outmux_3_27_port, O(26) => outmux_3_26_port, O(25) 
                           => outmux_3_25_port, O(24) => outmux_3_24_port, 
                           O(23) => outmux_3_23_port, O(22) => outmux_3_22_port
                           , O(21) => outmux_3_21_port, O(20) => 
                           outmux_3_20_port, O(19) => outmux_3_19_port, O(18) 
                           => outmux_3_18_port, O(17) => outmux_3_17_port, 
                           O(16) => outmux_3_16_port, O(15) => outmux_3_15_port
                           , O(14) => outmux_3_14_port, O(13) => 
                           outmux_3_13_port, O(12) => outmux_3_12_port, O(11) 
                           => outmux_3_11_port, O(10) => outmux_3_10_port, O(9)
                           => outmux_3_9_port, O(8) => outmux_3_8_port, O(7) =>
                           outmux_3_7_port, O(6) => outmux_3_6_port, O(5) => 
                           outmux_3_5_port, O(4) => outmux_3_4_port, O(3) => 
                           outmux_3_3_port, O(2) => outmux_3_2_port, O(1) => 
                           outmux_3_1_port, O(0) => outmux_3_0_port);
   MUXGEN_4 : mux_N32_4 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_4_31_port, B(30) => 
                           muxInB_4_30_port, B(29) => muxInB_4_29_port, B(28) 
                           => muxInB_4_28_port, B(27) => muxInB_4_27_port, 
                           B(26) => muxInB_4_26_port, B(25) => muxInB_4_25_port
                           , B(24) => muxInB_4_24_port, B(23) => 
                           muxInB_4_23_port, B(22) => muxInB_4_22_port, B(21) 
                           => muxInB_4_21_port, B(20) => muxInB_4_20_port, 
                           B(19) => muxInB_4_19_port, B(18) => muxInB_4_18_port
                           , B(17) => muxInB_4_17_port, B(16) => 
                           muxInB_4_16_port, B(15) => muxInB_4_15_port, B(14) 
                           => muxInB_4_14_port, B(13) => muxInB_4_13_port, 
                           B(12) => muxInB_4_12_port, B(11) => muxInB_4_11_port
                           , B(10) => muxInB_4_10_port, B(9) => muxInB_4_9_port
                           , B(8) => muxInB_4_8_port, B(7) => muxInB_4_7_port, 
                           B(6) => muxInB_4_6_port, B(5) => muxInB_4_5_port, 
                           B(4) => muxInB_4_4_port, B(3) => muxInB_4_3_port, 
                           B(2) => muxInB_4_2_port, B(1) => muxInB_4_1_port, 
                           B(0) => muxInB_4_0_port, C(31) => muxInC_4_31_port, 
                           C(30) => muxInC_4_30_port, C(29) => muxInC_4_29_port
                           , C(28) => muxInC_4_28_port, C(27) => 
                           muxInC_4_27_port, C(26) => muxInC_4_26_port, C(25) 
                           => muxInC_4_25_port, C(24) => muxInC_4_24_port, 
                           C(23) => muxInC_4_23_port, C(22) => muxInC_4_22_port
                           , C(21) => muxInC_4_21_port, C(20) => 
                           muxInC_4_20_port, C(19) => muxInC_4_19_port, C(18) 
                           => muxInC_4_18_port, C(17) => muxInC_4_17_port, 
                           C(16) => muxInC_4_16_port, C(15) => muxInC_4_15_port
                           , C(14) => muxInC_4_14_port, C(13) => 
                           muxInC_4_13_port, C(12) => muxInC_4_12_port, C(11) 
                           => muxInC_4_11_port, C(10) => muxInC_4_10_port, C(9)
                           => muxInC_4_9_port, C(8) => muxInC_4_8_port, C(7) =>
                           muxInC_4_7_port, C(6) => muxInC_4_6_port, C(5) => 
                           muxInC_4_5_port, C(4) => muxInC_4_4_port, C(3) => 
                           muxInC_4_3_port, C(2) => muxInC_4_2_port, C(1) => 
                           muxInC_4_1_port, C(0) => muxInC_4_0_port, D(31) => 
                           muxInD_4_31_port, D(30) => muxInD_4_30_port, D(29) 
                           => muxInD_4_29_port, D(28) => muxInD_4_28_port, 
                           D(27) => muxInD_4_27_port, D(26) => muxInD_4_26_port
                           , D(25) => muxInD_4_25_port, D(24) => 
                           muxInD_4_24_port, D(23) => muxInD_4_23_port, D(22) 
                           => muxInD_4_22_port, D(21) => muxInD_4_21_port, 
                           D(20) => muxInD_4_20_port, D(19) => muxInD_4_19_port
                           , D(18) => muxInD_4_18_port, D(17) => 
                           muxInD_4_17_port, D(16) => muxInD_4_16_port, D(15) 
                           => muxInD_4_15_port, D(14) => muxInD_4_14_port, 
                           D(13) => muxInD_4_13_port, D(12) => muxInD_4_12_port
                           , D(11) => muxInD_4_11_port, D(10) => 
                           muxInD_4_10_port, D(9) => muxInD_4_9_port, D(8) => 
                           muxInD_4_8_port, D(7) => muxInD_4_7_port, D(6) => 
                           muxInD_4_6_port, D(5) => muxInD_4_5_port, D(4) => 
                           muxInD_4_4_port, D(3) => muxInD_4_3_port, D(2) => 
                           muxInD_4_2_port, D(1) => muxInD_4_1_port, D(0) => 
                           muxInD_4_0_port, E(31) => muxInE_4_31_port, E(30) =>
                           muxInE_4_30_port, E(29) => muxInE_4_29_port, E(28) 
                           => muxInE_4_28_port, E(27) => muxInE_4_27_port, 
                           E(26) => muxInE_4_26_port, E(25) => muxInE_4_25_port
                           , E(24) => muxInE_4_24_port, E(23) => 
                           muxInE_4_23_port, E(22) => muxInE_4_22_port, E(21) 
                           => muxInE_4_21_port, E(20) => muxInE_4_20_port, 
                           E(19) => muxInE_4_19_port, E(18) => muxInE_4_18_port
                           , E(17) => muxInE_4_17_port, E(16) => 
                           muxInE_4_16_port, E(15) => muxInE_4_15_port, E(14) 
                           => muxInE_4_14_port, E(13) => muxInE_4_13_port, 
                           E(12) => muxInE_4_12_port, E(11) => muxInE_4_11_port
                           , E(10) => muxInE_4_10_port, E(9) => muxInE_4_9_port
                           , E(8) => muxInE_4_8_port, E(7) => muxInE_4_7_port, 
                           E(6) => muxInE_4_6_port, E(5) => muxInE_4_5_port, 
                           E(4) => muxInE_4_4_port, E(3) => muxInE_4_3_port, 
                           E(2) => muxInE_4_2_port, E(1) => muxInE_4_1_port, 
                           E(0) => muxInE_4_0_port, Sel(2) => B(9), Sel(1) => 
                           B(8), Sel(0) => B(7), O(31) => outmux_4_31_port, 
                           O(30) => outmux_4_30_port, O(29) => outmux_4_29_port
                           , O(28) => outmux_4_28_port, O(27) => 
                           outmux_4_27_port, O(26) => outmux_4_26_port, O(25) 
                           => outmux_4_25_port, O(24) => outmux_4_24_port, 
                           O(23) => outmux_4_23_port, O(22) => outmux_4_22_port
                           , O(21) => outmux_4_21_port, O(20) => 
                           outmux_4_20_port, O(19) => outmux_4_19_port, O(18) 
                           => outmux_4_18_port, O(17) => outmux_4_17_port, 
                           O(16) => outmux_4_16_port, O(15) => outmux_4_15_port
                           , O(14) => outmux_4_14_port, O(13) => 
                           outmux_4_13_port, O(12) => outmux_4_12_port, O(11) 
                           => outmux_4_11_port, O(10) => outmux_4_10_port, O(9)
                           => outmux_4_9_port, O(8) => outmux_4_8_port, O(7) =>
                           outmux_4_7_port, O(6) => outmux_4_6_port, O(5) => 
                           outmux_4_5_port, O(4) => outmux_4_4_port, O(3) => 
                           outmux_4_3_port, O(2) => outmux_4_2_port, O(1) => 
                           outmux_4_1_port, O(0) => outmux_4_0_port);
   MUXGEN_5 : mux_N32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_5_31_port, B(30) => 
                           muxInB_5_30_port, B(29) => muxInB_5_29_port, B(28) 
                           => muxInB_5_28_port, B(27) => muxInB_5_27_port, 
                           B(26) => muxInB_5_26_port, B(25) => muxInB_5_25_port
                           , B(24) => muxInB_5_24_port, B(23) => 
                           muxInB_5_23_port, B(22) => muxInB_5_22_port, B(21) 
                           => muxInB_5_21_port, B(20) => muxInB_5_20_port, 
                           B(19) => muxInB_5_19_port, B(18) => muxInB_5_18_port
                           , B(17) => muxInB_5_17_port, B(16) => 
                           muxInB_5_16_port, B(15) => muxInB_5_15_port, B(14) 
                           => muxInB_5_14_port, B(13) => muxInB_5_13_port, 
                           B(12) => muxInB_5_12_port, B(11) => muxInB_5_11_port
                           , B(10) => muxInB_5_10_port, B(9) => muxInB_5_9_port
                           , B(8) => muxInB_5_8_port, B(7) => muxInB_5_7_port, 
                           B(6) => muxInB_5_6_port, B(5) => muxInB_5_5_port, 
                           B(4) => muxInB_5_4_port, B(3) => muxInB_5_3_port, 
                           B(2) => muxInB_5_2_port, B(1) => muxInB_5_1_port, 
                           B(0) => muxInB_5_0_port, C(31) => muxInC_5_31_port, 
                           C(30) => muxInC_5_30_port, C(29) => muxInC_5_29_port
                           , C(28) => muxInC_5_28_port, C(27) => 
                           muxInC_5_27_port, C(26) => muxInC_5_26_port, C(25) 
                           => muxInC_5_25_port, C(24) => muxInC_5_24_port, 
                           C(23) => muxInC_5_23_port, C(22) => muxInC_5_22_port
                           , C(21) => muxInC_5_21_port, C(20) => 
                           muxInC_5_20_port, C(19) => muxInC_5_19_port, C(18) 
                           => muxInC_5_18_port, C(17) => muxInC_5_17_port, 
                           C(16) => muxInC_5_16_port, C(15) => muxInC_5_15_port
                           , C(14) => muxInC_5_14_port, C(13) => 
                           muxInC_5_13_port, C(12) => muxInC_5_12_port, C(11) 
                           => muxInC_5_11_port, C(10) => muxInC_5_10_port, C(9)
                           => muxInC_5_9_port, C(8) => muxInC_5_8_port, C(7) =>
                           muxInC_5_7_port, C(6) => muxInC_5_6_port, C(5) => 
                           muxInC_5_5_port, C(4) => muxInC_5_4_port, C(3) => 
                           muxInC_5_3_port, C(2) => muxInC_5_2_port, C(1) => 
                           muxInC_5_1_port, C(0) => muxInC_5_0_port, D(31) => 
                           muxInD_5_31_port, D(30) => muxInD_5_30_port, D(29) 
                           => muxInD_5_29_port, D(28) => muxInD_5_28_port, 
                           D(27) => muxInD_5_27_port, D(26) => muxInD_5_26_port
                           , D(25) => muxInD_5_25_port, D(24) => 
                           muxInD_5_24_port, D(23) => muxInD_5_23_port, D(22) 
                           => muxInD_5_22_port, D(21) => muxInD_5_21_port, 
                           D(20) => muxInD_5_20_port, D(19) => muxInD_5_19_port
                           , D(18) => muxInD_5_18_port, D(17) => 
                           muxInD_5_17_port, D(16) => muxInD_5_16_port, D(15) 
                           => muxInD_5_15_port, D(14) => muxInD_5_14_port, 
                           D(13) => muxInD_5_13_port, D(12) => muxInD_5_12_port
                           , D(11) => muxInD_5_11_port, D(10) => 
                           muxInD_5_10_port, D(9) => muxInD_5_9_port, D(8) => 
                           muxInD_5_8_port, D(7) => muxInD_5_7_port, D(6) => 
                           muxInD_5_6_port, D(5) => muxInD_5_5_port, D(4) => 
                           muxInD_5_4_port, D(3) => muxInD_5_3_port, D(2) => 
                           muxInD_5_2_port, D(1) => muxInD_5_1_port, D(0) => 
                           muxInD_5_0_port, E(31) => muxInE_5_31_port, E(30) =>
                           muxInE_5_30_port, E(29) => muxInE_5_29_port, E(28) 
                           => muxInE_5_28_port, E(27) => muxInE_5_27_port, 
                           E(26) => muxInE_5_26_port, E(25) => muxInE_5_25_port
                           , E(24) => muxInE_5_24_port, E(23) => 
                           muxInE_5_23_port, E(22) => muxInE_5_22_port, E(21) 
                           => muxInE_5_21_port, E(20) => muxInE_5_20_port, 
                           E(19) => muxInE_5_19_port, E(18) => muxInE_5_18_port
                           , E(17) => muxInE_5_17_port, E(16) => 
                           muxInE_5_16_port, E(15) => muxInE_5_15_port, E(14) 
                           => muxInE_5_14_port, E(13) => muxInE_5_13_port, 
                           E(12) => muxInE_5_12_port, E(11) => muxInE_5_11_port
                           , E(10) => muxInE_5_10_port, E(9) => muxInE_5_9_port
                           , E(8) => muxInE_5_8_port, E(7) => muxInE_5_7_port, 
                           E(6) => muxInE_5_6_port, E(5) => muxInE_5_5_port, 
                           E(4) => muxInE_5_4_port, E(3) => muxInE_5_3_port, 
                           E(2) => muxInE_5_2_port, E(1) => muxInE_5_1_port, 
                           E(0) => muxInE_5_0_port, Sel(2) => B(11), Sel(1) => 
                           B(10), Sel(0) => B(9), O(31) => outmux_5_31_port, 
                           O(30) => outmux_5_30_port, O(29) => outmux_5_29_port
                           , O(28) => outmux_5_28_port, O(27) => 
                           outmux_5_27_port, O(26) => outmux_5_26_port, O(25) 
                           => outmux_5_25_port, O(24) => outmux_5_24_port, 
                           O(23) => outmux_5_23_port, O(22) => outmux_5_22_port
                           , O(21) => outmux_5_21_port, O(20) => 
                           outmux_5_20_port, O(19) => outmux_5_19_port, O(18) 
                           => outmux_5_18_port, O(17) => outmux_5_17_port, 
                           O(16) => outmux_5_16_port, O(15) => outmux_5_15_port
                           , O(14) => outmux_5_14_port, O(13) => 
                           outmux_5_13_port, O(12) => outmux_5_12_port, O(11) 
                           => outmux_5_11_port, O(10) => outmux_5_10_port, O(9)
                           => outmux_5_9_port, O(8) => outmux_5_8_port, O(7) =>
                           outmux_5_7_port, O(6) => outmux_5_6_port, O(5) => 
                           outmux_5_5_port, O(4) => outmux_5_4_port, O(3) => 
                           outmux_5_3_port, O(2) => outmux_5_2_port, O(1) => 
                           outmux_5_1_port, O(0) => outmux_5_0_port);
   MUXGEN_6 : mux_N32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_6_31_port, B(30) => 
                           muxInB_6_30_port, B(29) => muxInB_6_29_port, B(28) 
                           => muxInB_6_28_port, B(27) => muxInB_6_27_port, 
                           B(26) => muxInB_6_26_port, B(25) => muxInB_6_25_port
                           , B(24) => muxInB_6_24_port, B(23) => 
                           muxInB_6_23_port, B(22) => muxInB_6_22_port, B(21) 
                           => muxInB_6_21_port, B(20) => muxInB_6_20_port, 
                           B(19) => muxInB_6_19_port, B(18) => muxInB_6_18_port
                           , B(17) => muxInB_6_17_port, B(16) => 
                           muxInB_6_16_port, B(15) => muxInB_6_15_port, B(14) 
                           => muxInB_6_14_port, B(13) => muxInB_6_13_port, 
                           B(12) => muxInB_6_12_port, B(11) => muxInB_6_11_port
                           , B(10) => muxInB_6_10_port, B(9) => muxInB_6_9_port
                           , B(8) => muxInB_6_8_port, B(7) => muxInB_6_7_port, 
                           B(6) => muxInB_6_6_port, B(5) => muxInB_6_5_port, 
                           B(4) => muxInB_6_4_port, B(3) => muxInB_6_3_port, 
                           B(2) => muxInB_6_2_port, B(1) => muxInB_6_1_port, 
                           B(0) => muxInB_6_0_port, C(31) => muxInC_6_31_port, 
                           C(30) => muxInC_6_30_port, C(29) => muxInC_6_29_port
                           , C(28) => muxInC_6_28_port, C(27) => 
                           muxInC_6_27_port, C(26) => muxInC_6_26_port, C(25) 
                           => muxInC_6_25_port, C(24) => muxInC_6_24_port, 
                           C(23) => muxInC_6_23_port, C(22) => muxInC_6_22_port
                           , C(21) => muxInC_6_21_port, C(20) => 
                           muxInC_6_20_port, C(19) => muxInC_6_19_port, C(18) 
                           => muxInC_6_18_port, C(17) => muxInC_6_17_port, 
                           C(16) => muxInC_6_16_port, C(15) => muxInC_6_15_port
                           , C(14) => muxInC_6_14_port, C(13) => 
                           muxInC_6_13_port, C(12) => muxInC_6_12_port, C(11) 
                           => muxInC_6_11_port, C(10) => muxInC_6_10_port, C(9)
                           => muxInC_6_9_port, C(8) => muxInC_6_8_port, C(7) =>
                           muxInC_6_7_port, C(6) => muxInC_6_6_port, C(5) => 
                           muxInC_6_5_port, C(4) => muxInC_6_4_port, C(3) => 
                           muxInC_6_3_port, C(2) => muxInC_6_2_port, C(1) => 
                           muxInC_6_1_port, C(0) => muxInC_6_0_port, D(31) => 
                           muxInD_6_31_port, D(30) => muxInD_6_30_port, D(29) 
                           => muxInD_6_29_port, D(28) => muxInD_6_28_port, 
                           D(27) => muxInD_6_27_port, D(26) => muxInD_6_26_port
                           , D(25) => muxInD_6_25_port, D(24) => 
                           muxInD_6_24_port, D(23) => muxInD_6_23_port, D(22) 
                           => muxInD_6_22_port, D(21) => muxInD_6_21_port, 
                           D(20) => muxInD_6_20_port, D(19) => muxInD_6_19_port
                           , D(18) => muxInD_6_18_port, D(17) => 
                           muxInD_6_17_port, D(16) => muxInD_6_16_port, D(15) 
                           => muxInD_6_15_port, D(14) => muxInD_6_14_port, 
                           D(13) => muxInD_6_13_port, D(12) => muxInD_6_12_port
                           , D(11) => muxInD_6_11_port, D(10) => 
                           muxInD_6_10_port, D(9) => muxInD_6_9_port, D(8) => 
                           muxInD_6_8_port, D(7) => muxInD_6_7_port, D(6) => 
                           muxInD_6_6_port, D(5) => muxInD_6_5_port, D(4) => 
                           muxInD_6_4_port, D(3) => muxInD_6_3_port, D(2) => 
                           muxInD_6_2_port, D(1) => muxInD_6_1_port, D(0) => 
                           muxInD_6_0_port, E(31) => muxInE_6_31_port, E(30) =>
                           muxInE_6_30_port, E(29) => muxInE_6_29_port, E(28) 
                           => muxInE_6_28_port, E(27) => muxInE_6_27_port, 
                           E(26) => muxInE_6_26_port, E(25) => muxInE_6_25_port
                           , E(24) => muxInE_6_24_port, E(23) => 
                           muxInE_6_23_port, E(22) => muxInE_6_22_port, E(21) 
                           => muxInE_6_21_port, E(20) => muxInE_6_20_port, 
                           E(19) => muxInE_6_19_port, E(18) => muxInE_6_18_port
                           , E(17) => muxInE_6_17_port, E(16) => 
                           muxInE_6_16_port, E(15) => muxInE_6_15_port, E(14) 
                           => muxInE_6_14_port, E(13) => muxInE_6_13_port, 
                           E(12) => muxInE_6_12_port, E(11) => muxInE_6_11_port
                           , E(10) => muxInE_6_10_port, E(9) => muxInE_6_9_port
                           , E(8) => muxInE_6_8_port, E(7) => muxInE_6_7_port, 
                           E(6) => muxInE_6_6_port, E(5) => muxInE_6_5_port, 
                           E(4) => muxInE_6_4_port, E(3) => muxInE_6_3_port, 
                           E(2) => muxInE_6_2_port, E(1) => muxInE_6_1_port, 
                           E(0) => muxInE_6_0_port, Sel(2) => B(13), Sel(1) => 
                           B(12), Sel(0) => B(11), O(31) => outmux_6_31_port, 
                           O(30) => outmux_6_30_port, O(29) => outmux_6_29_port
                           , O(28) => outmux_6_28_port, O(27) => 
                           outmux_6_27_port, O(26) => outmux_6_26_port, O(25) 
                           => outmux_6_25_port, O(24) => outmux_6_24_port, 
                           O(23) => outmux_6_23_port, O(22) => outmux_6_22_port
                           , O(21) => outmux_6_21_port, O(20) => 
                           outmux_6_20_port, O(19) => outmux_6_19_port, O(18) 
                           => outmux_6_18_port, O(17) => outmux_6_17_port, 
                           O(16) => outmux_6_16_port, O(15) => outmux_6_15_port
                           , O(14) => outmux_6_14_port, O(13) => 
                           outmux_6_13_port, O(12) => outmux_6_12_port, O(11) 
                           => outmux_6_11_port, O(10) => outmux_6_10_port, O(9)
                           => outmux_6_9_port, O(8) => outmux_6_8_port, O(7) =>
                           outmux_6_7_port, O(6) => outmux_6_6_port, O(5) => 
                           outmux_6_5_port, O(4) => outmux_6_4_port, O(3) => 
                           outmux_6_3_port, O(2) => outmux_6_2_port, O(1) => 
                           outmux_6_1_port, O(0) => outmux_6_0_port);
   MUXGEN_7 : mux_N32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_7_31_port, B(30) => 
                           muxInB_7_30_port, B(29) => muxInB_7_29_port, B(28) 
                           => muxInB_7_28_port, B(27) => muxInB_7_27_port, 
                           B(26) => muxInB_7_26_port, B(25) => muxInB_7_25_port
                           , B(24) => muxInB_7_24_port, B(23) => 
                           muxInB_7_23_port, B(22) => muxInB_7_22_port, B(21) 
                           => muxInB_7_21_port, B(20) => muxInB_7_20_port, 
                           B(19) => muxInB_7_19_port, B(18) => muxInB_7_18_port
                           , B(17) => muxInB_7_17_port, B(16) => 
                           muxInB_7_16_port, B(15) => muxInB_7_15_port, B(14) 
                           => muxInB_7_14_port, B(13) => muxInB_7_13_port, 
                           B(12) => muxInB_7_12_port, B(11) => muxInB_7_11_port
                           , B(10) => muxInB_7_10_port, B(9) => muxInB_7_9_port
                           , B(8) => muxInB_7_8_port, B(7) => muxInB_7_7_port, 
                           B(6) => muxInB_7_6_port, B(5) => muxInB_7_5_port, 
                           B(4) => muxInB_7_4_port, B(3) => muxInB_7_3_port, 
                           B(2) => muxInB_7_2_port, B(1) => muxInB_7_1_port, 
                           B(0) => muxInB_7_0_port, C(31) => muxInC_7_31_port, 
                           C(30) => muxInC_7_30_port, C(29) => muxInC_7_29_port
                           , C(28) => muxInC_7_28_port, C(27) => 
                           muxInC_7_27_port, C(26) => muxInC_7_26_port, C(25) 
                           => muxInC_7_25_port, C(24) => muxInC_7_24_port, 
                           C(23) => muxInC_7_23_port, C(22) => muxInC_7_22_port
                           , C(21) => muxInC_7_21_port, C(20) => 
                           muxInC_7_20_port, C(19) => muxInC_7_19_port, C(18) 
                           => muxInC_7_18_port, C(17) => muxInC_7_17_port, 
                           C(16) => muxInC_7_16_port, C(15) => muxInC_7_15_port
                           , C(14) => muxInC_7_14_port, C(13) => 
                           muxInC_7_13_port, C(12) => muxInC_7_12_port, C(11) 
                           => muxInC_7_11_port, C(10) => muxInC_7_10_port, C(9)
                           => muxInC_7_9_port, C(8) => muxInC_7_8_port, C(7) =>
                           muxInC_7_7_port, C(6) => muxInC_7_6_port, C(5) => 
                           muxInC_7_5_port, C(4) => muxInC_7_4_port, C(3) => 
                           muxInC_7_3_port, C(2) => muxInC_7_2_port, C(1) => 
                           muxInC_7_1_port, C(0) => muxInC_7_0_port, D(31) => 
                           muxInD_7_31_port, D(30) => muxInD_7_30_port, D(29) 
                           => muxInD_7_29_port, D(28) => muxInD_7_28_port, 
                           D(27) => muxInD_7_27_port, D(26) => muxInD_7_26_port
                           , D(25) => muxInD_7_25_port, D(24) => 
                           muxInD_7_24_port, D(23) => muxInD_7_23_port, D(22) 
                           => muxInD_7_22_port, D(21) => muxInD_7_21_port, 
                           D(20) => muxInD_7_20_port, D(19) => muxInD_7_19_port
                           , D(18) => muxInD_7_18_port, D(17) => 
                           muxInD_7_17_port, D(16) => muxInD_7_16_port, D(15) 
                           => muxInD_7_15_port, D(14) => muxInD_7_14_port, 
                           D(13) => muxInD_7_13_port, D(12) => muxInD_7_12_port
                           , D(11) => muxInD_7_11_port, D(10) => 
                           muxInD_7_10_port, D(9) => muxInD_7_9_port, D(8) => 
                           muxInD_7_8_port, D(7) => muxInD_7_7_port, D(6) => 
                           muxInD_7_6_port, D(5) => muxInD_7_5_port, D(4) => 
                           muxInD_7_4_port, D(3) => muxInD_7_3_port, D(2) => 
                           muxInD_7_2_port, D(1) => muxInD_7_1_port, D(0) => 
                           muxInD_7_0_port, E(31) => muxInE_7_31_port, E(30) =>
                           muxInE_7_30_port, E(29) => muxInE_7_29_port, E(28) 
                           => muxInE_7_28_port, E(27) => muxInE_7_27_port, 
                           E(26) => muxInE_7_26_port, E(25) => muxInE_7_25_port
                           , E(24) => muxInE_7_24_port, E(23) => 
                           muxInE_7_23_port, E(22) => muxInE_7_22_port, E(21) 
                           => muxInE_7_21_port, E(20) => muxInE_7_20_port, 
                           E(19) => muxInE_7_19_port, E(18) => muxInE_7_18_port
                           , E(17) => muxInE_7_17_port, E(16) => 
                           muxInE_7_16_port, E(15) => muxInE_7_15_port, E(14) 
                           => muxInE_7_14_port, E(13) => muxInE_7_13_port, 
                           E(12) => muxInE_7_12_port, E(11) => muxInE_7_11_port
                           , E(10) => muxInE_7_10_port, E(9) => muxInE_7_9_port
                           , E(8) => muxInE_7_8_port, E(7) => muxInE_7_7_port, 
                           E(6) => muxInE_7_6_port, E(5) => muxInE_7_5_port, 
                           E(4) => muxInE_7_4_port, E(3) => muxInE_7_3_port, 
                           E(2) => muxInE_7_2_port, E(1) => muxInE_7_1_port, 
                           E(0) => muxInE_7_0_port, Sel(2) => B(15), Sel(1) => 
                           B(14), Sel(0) => B(13), O(31) => outmux_7_31_port, 
                           O(30) => outmux_7_30_port, O(29) => outmux_7_29_port
                           , O(28) => outmux_7_28_port, O(27) => 
                           outmux_7_27_port, O(26) => outmux_7_26_port, O(25) 
                           => outmux_7_25_port, O(24) => outmux_7_24_port, 
                           O(23) => outmux_7_23_port, O(22) => outmux_7_22_port
                           , O(21) => outmux_7_21_port, O(20) => 
                           outmux_7_20_port, O(19) => outmux_7_19_port, O(18) 
                           => outmux_7_18_port, O(17) => outmux_7_17_port, 
                           O(16) => outmux_7_16_port, O(15) => outmux_7_15_port
                           , O(14) => outmux_7_14_port, O(13) => 
                           outmux_7_13_port, O(12) => outmux_7_12_port, O(11) 
                           => outmux_7_11_port, O(10) => outmux_7_10_port, O(9)
                           => outmux_7_9_port, O(8) => outmux_7_8_port, O(7) =>
                           outmux_7_7_port, O(6) => outmux_7_6_port, O(5) => 
                           outmux_7_5_port, O(4) => outmux_7_4_port, O(3) => 
                           outmux_7_3_port, O(2) => outmux_7_2_port, O(1) => 
                           outmux_7_1_port, O(0) => outmux_7_0_port);
   Add1IL : CSA_Nbits32_0 port map( A(31) => outmux_0_31_port, A(30) => 
                           outmux_0_30_port, A(29) => outmux_0_29_port, A(28) 
                           => outmux_0_28_port, A(27) => outmux_0_27_port, 
                           A(26) => outmux_0_26_port, A(25) => outmux_0_25_port
                           , A(24) => outmux_0_24_port, A(23) => 
                           outmux_0_23_port, A(22) => outmux_0_22_port, A(21) 
                           => outmux_0_21_port, A(20) => outmux_0_20_port, 
                           A(19) => outmux_0_19_port, A(18) => outmux_0_18_port
                           , A(17) => outmux_0_17_port, A(16) => 
                           outmux_0_16_port, A(15) => outmux_0_15_port, A(14) 
                           => outmux_0_14_port, A(13) => outmux_0_13_port, 
                           A(12) => outmux_0_12_port, A(11) => outmux_0_11_port
                           , A(10) => outmux_0_10_port, A(9) => outmux_0_9_port
                           , A(8) => outmux_0_8_port, A(7) => outmux_0_7_port, 
                           A(6) => outmux_0_6_port, A(5) => outmux_0_5_port, 
                           A(4) => outmux_0_4_port, A(3) => outmux_0_3_port, 
                           A(2) => outmux_0_2_port, A(1) => outmux_0_1_port, 
                           A(0) => outmux_0_0_port, B(31) => outmux_1_31_port, 
                           B(30) => outmux_1_30_port, B(29) => outmux_1_29_port
                           , B(28) => outmux_1_28_port, B(27) => 
                           outmux_1_27_port, B(26) => outmux_1_26_port, B(25) 
                           => outmux_1_25_port, B(24) => outmux_1_24_port, 
                           B(23) => outmux_1_23_port, B(22) => outmux_1_22_port
                           , B(21) => outmux_1_21_port, B(20) => 
                           outmux_1_20_port, B(19) => outmux_1_19_port, B(18) 
                           => outmux_1_18_port, B(17) => outmux_1_17_port, 
                           B(16) => outmux_1_16_port, B(15) => outmux_1_15_port
                           , B(14) => outmux_1_14_port, B(13) => 
                           outmux_1_13_port, B(12) => outmux_1_12_port, B(11) 
                           => outmux_1_11_port, B(10) => outmux_1_10_port, B(9)
                           => outmux_1_9_port, B(8) => outmux_1_8_port, B(7) =>
                           outmux_1_7_port, B(6) => outmux_1_6_port, B(5) => 
                           outmux_1_5_port, B(4) => outmux_1_4_port, B(3) => 
                           outmux_1_3_port, B(2) => outmux_1_2_port, B(1) => 
                           outmux_1_1_port, B(0) => outmux_1_0_port, C(31) => 
                           outmux_2_31_port, C(30) => outmux_2_30_port, C(29) 
                           => outmux_2_29_port, C(28) => outmux_2_28_port, 
                           C(27) => outmux_2_27_port, C(26) => outmux_2_26_port
                           , C(25) => outmux_2_25_port, C(24) => 
                           outmux_2_24_port, C(23) => outmux_2_23_port, C(22) 
                           => outmux_2_22_port, C(21) => outmux_2_21_port, 
                           C(20) => outmux_2_20_port, C(19) => outmux_2_19_port
                           , C(18) => outmux_2_18_port, C(17) => 
                           outmux_2_17_port, C(16) => outmux_2_16_port, C(15) 
                           => outmux_2_15_port, C(14) => outmux_2_14_port, 
                           C(13) => outmux_2_13_port, C(12) => outmux_2_12_port
                           , C(11) => outmux_2_11_port, C(10) => 
                           outmux_2_10_port, C(9) => outmux_2_9_port, C(8) => 
                           outmux_2_8_port, C(7) => outmux_2_7_port, C(6) => 
                           outmux_2_6_port, C(5) => outmux_2_5_port, C(4) => 
                           outmux_2_4_port, C(3) => outmux_2_3_port, C(2) => 
                           outmux_2_2_port, C(1) => outmux_2_1_port, C(0) => 
                           outmux_2_0_port, S(31) => sum_array_0_31_port, S(30)
                           => sum_array_0_30_port, S(29) => sum_array_0_29_port
                           , S(28) => sum_array_0_28_port, S(27) => 
                           sum_array_0_27_port, S(26) => sum_array_0_26_port, 
                           S(25) => sum_array_0_25_port, S(24) => 
                           sum_array_0_24_port, S(23) => sum_array_0_23_port, 
                           S(22) => sum_array_0_22_port, S(21) => 
                           sum_array_0_21_port, S(20) => sum_array_0_20_port, 
                           S(19) => sum_array_0_19_port, S(18) => 
                           sum_array_0_18_port, S(17) => sum_array_0_17_port, 
                           S(16) => sum_array_0_16_port, S(15) => 
                           sum_array_0_15_port, S(14) => sum_array_0_14_port, 
                           S(13) => sum_array_0_13_port, S(12) => 
                           sum_array_0_12_port, S(11) => sum_array_0_11_port, 
                           S(10) => sum_array_0_10_port, S(9) => 
                           sum_array_0_9_port, S(8) => sum_array_0_8_port, S(7)
                           => sum_array_0_7_port, S(6) => sum_array_0_6_port, 
                           S(5) => sum_array_0_5_port, S(4) => 
                           sum_array_0_4_port, S(3) => sum_array_0_3_port, S(2)
                           => sum_array_0_2_port, S(1) => sum_array_0_1_port, 
                           S(0) => sum_array_0_0_port, Cout(31) => 
                           cout_array_0_31_port, Cout(30) => 
                           cout_array_0_30_port, Cout(29) => 
                           cout_array_0_29_port, Cout(28) => 
                           cout_array_0_28_port, Cout(27) => 
                           cout_array_0_27_port, Cout(26) => 
                           cout_array_0_26_port, Cout(25) => 
                           cout_array_0_25_port, Cout(24) => 
                           cout_array_0_24_port, Cout(23) => 
                           cout_array_0_23_port, Cout(22) => 
                           cout_array_0_22_port, Cout(21) => 
                           cout_array_0_21_port, Cout(20) => 
                           cout_array_0_20_port, Cout(19) => 
                           cout_array_0_19_port, Cout(18) => 
                           cout_array_0_18_port, Cout(17) => 
                           cout_array_0_17_port, Cout(16) => 
                           cout_array_0_16_port, Cout(15) => 
                           cout_array_0_15_port, Cout(14) => 
                           cout_array_0_14_port, Cout(13) => 
                           cout_array_0_13_port, Cout(12) => 
                           cout_array_0_12_port, Cout(11) => 
                           cout_array_0_11_port, Cout(10) => 
                           cout_array_0_10_port, Cout(9) => cout_array_0_9_port
                           , Cout(8) => cout_array_0_8_port, Cout(7) => 
                           cout_array_0_7_port, Cout(6) => cout_array_0_6_port,
                           Cout(5) => cout_array_0_5_port, Cout(4) => 
                           cout_array_0_4_port, Cout(3) => cout_array_0_3_port,
                           Cout(2) => cout_array_0_2_port, Cout(1) => 
                           cout_array_0_1_port, Cout(0) => net59834);
   Add2IL : CSA_Nbits32_5 port map( A(31) => outmux_3_31_port, A(30) => 
                           outmux_3_30_port, A(29) => outmux_3_29_port, A(28) 
                           => outmux_3_28_port, A(27) => outmux_3_27_port, 
                           A(26) => outmux_3_26_port, A(25) => outmux_3_25_port
                           , A(24) => outmux_3_24_port, A(23) => 
                           outmux_3_23_port, A(22) => outmux_3_22_port, A(21) 
                           => outmux_3_21_port, A(20) => outmux_3_20_port, 
                           A(19) => outmux_3_19_port, A(18) => outmux_3_18_port
                           , A(17) => outmux_3_17_port, A(16) => 
                           outmux_3_16_port, A(15) => outmux_3_15_port, A(14) 
                           => outmux_3_14_port, A(13) => outmux_3_13_port, 
                           A(12) => outmux_3_12_port, A(11) => outmux_3_11_port
                           , A(10) => outmux_3_10_port, A(9) => outmux_3_9_port
                           , A(8) => outmux_3_8_port, A(7) => outmux_3_7_port, 
                           A(6) => outmux_3_6_port, A(5) => outmux_3_5_port, 
                           A(4) => outmux_3_4_port, A(3) => outmux_3_3_port, 
                           A(2) => outmux_3_2_port, A(1) => outmux_3_1_port, 
                           A(0) => outmux_3_0_port, B(31) => outmux_4_31_port, 
                           B(30) => outmux_4_30_port, B(29) => outmux_4_29_port
                           , B(28) => outmux_4_28_port, B(27) => 
                           outmux_4_27_port, B(26) => outmux_4_26_port, B(25) 
                           => outmux_4_25_port, B(24) => outmux_4_24_port, 
                           B(23) => outmux_4_23_port, B(22) => outmux_4_22_port
                           , B(21) => outmux_4_21_port, B(20) => 
                           outmux_4_20_port, B(19) => outmux_4_19_port, B(18) 
                           => outmux_4_18_port, B(17) => outmux_4_17_port, 
                           B(16) => outmux_4_16_port, B(15) => outmux_4_15_port
                           , B(14) => outmux_4_14_port, B(13) => 
                           outmux_4_13_port, B(12) => outmux_4_12_port, B(11) 
                           => outmux_4_11_port, B(10) => outmux_4_10_port, B(9)
                           => outmux_4_9_port, B(8) => outmux_4_8_port, B(7) =>
                           outmux_4_7_port, B(6) => outmux_4_6_port, B(5) => 
                           outmux_4_5_port, B(4) => outmux_4_4_port, B(3) => 
                           outmux_4_3_port, B(2) => outmux_4_2_port, B(1) => 
                           outmux_4_1_port, B(0) => outmux_4_0_port, C(31) => 
                           outmux_5_31_port, C(30) => outmux_5_30_port, C(29) 
                           => outmux_5_29_port, C(28) => outmux_5_28_port, 
                           C(27) => outmux_5_27_port, C(26) => outmux_5_26_port
                           , C(25) => outmux_5_25_port, C(24) => 
                           outmux_5_24_port, C(23) => outmux_5_23_port, C(22) 
                           => outmux_5_22_port, C(21) => outmux_5_21_port, 
                           C(20) => outmux_5_20_port, C(19) => outmux_5_19_port
                           , C(18) => outmux_5_18_port, C(17) => 
                           outmux_5_17_port, C(16) => outmux_5_16_port, C(15) 
                           => outmux_5_15_port, C(14) => outmux_5_14_port, 
                           C(13) => outmux_5_13_port, C(12) => outmux_5_12_port
                           , C(11) => outmux_5_11_port, C(10) => 
                           outmux_5_10_port, C(9) => outmux_5_9_port, C(8) => 
                           outmux_5_8_port, C(7) => outmux_5_7_port, C(6) => 
                           outmux_5_6_port, C(5) => outmux_5_5_port, C(4) => 
                           outmux_5_4_port, C(3) => outmux_5_3_port, C(2) => 
                           outmux_5_2_port, C(1) => outmux_5_1_port, C(0) => 
                           outmux_5_0_port, S(31) => sum_array_1_31_port, S(30)
                           => sum_array_1_30_port, S(29) => sum_array_1_29_port
                           , S(28) => sum_array_1_28_port, S(27) => 
                           sum_array_1_27_port, S(26) => sum_array_1_26_port, 
                           S(25) => sum_array_1_25_port, S(24) => 
                           sum_array_1_24_port, S(23) => sum_array_1_23_port, 
                           S(22) => sum_array_1_22_port, S(21) => 
                           sum_array_1_21_port, S(20) => sum_array_1_20_port, 
                           S(19) => sum_array_1_19_port, S(18) => 
                           sum_array_1_18_port, S(17) => sum_array_1_17_port, 
                           S(16) => sum_array_1_16_port, S(15) => 
                           sum_array_1_15_port, S(14) => sum_array_1_14_port, 
                           S(13) => sum_array_1_13_port, S(12) => 
                           sum_array_1_12_port, S(11) => sum_array_1_11_port, 
                           S(10) => sum_array_1_10_port, S(9) => 
                           sum_array_1_9_port, S(8) => sum_array_1_8_port, S(7)
                           => sum_array_1_7_port, S(6) => sum_array_1_6_port, 
                           S(5) => sum_array_1_5_port, S(4) => 
                           sum_array_1_4_port, S(3) => sum_array_1_3_port, S(2)
                           => sum_array_1_2_port, S(1) => sum_array_1_1_port, 
                           S(0) => sum_array_1_0_port, Cout(31) => 
                           cout_array_1_31_port, Cout(30) => 
                           cout_array_1_30_port, Cout(29) => 
                           cout_array_1_29_port, Cout(28) => 
                           cout_array_1_28_port, Cout(27) => 
                           cout_array_1_27_port, Cout(26) => 
                           cout_array_1_26_port, Cout(25) => 
                           cout_array_1_25_port, Cout(24) => 
                           cout_array_1_24_port, Cout(23) => 
                           cout_array_1_23_port, Cout(22) => 
                           cout_array_1_22_port, Cout(21) => 
                           cout_array_1_21_port, Cout(20) => 
                           cout_array_1_20_port, Cout(19) => 
                           cout_array_1_19_port, Cout(18) => 
                           cout_array_1_18_port, Cout(17) => 
                           cout_array_1_17_port, Cout(16) => 
                           cout_array_1_16_port, Cout(15) => 
                           cout_array_1_15_port, Cout(14) => 
                           cout_array_1_14_port, Cout(13) => 
                           cout_array_1_13_port, Cout(12) => 
                           cout_array_1_12_port, Cout(11) => 
                           cout_array_1_11_port, Cout(10) => 
                           cout_array_1_10_port, Cout(9) => cout_array_1_9_port
                           , Cout(8) => cout_array_1_8_port, Cout(7) => 
                           cout_array_1_7_port, Cout(6) => cout_array_1_6_port,
                           Cout(5) => cout_array_1_5_port, Cout(4) => 
                           cout_array_1_4_port, Cout(3) => cout_array_1_3_port,
                           Cout(2) => cout_array_1_2_port, Cout(1) => 
                           cout_array_1_1_port, Cout(0) => net59833);
   Add1IIL : CSA_Nbits32_4 port map( A(31) => sum_array_0_31_port, A(30) => 
                           sum_array_0_30_port, A(29) => sum_array_0_29_port, 
                           A(28) => sum_array_0_28_port, A(27) => 
                           sum_array_0_27_port, A(26) => sum_array_0_26_port, 
                           A(25) => sum_array_0_25_port, A(24) => 
                           sum_array_0_24_port, A(23) => sum_array_0_23_port, 
                           A(22) => sum_array_0_22_port, A(21) => 
                           sum_array_0_21_port, A(20) => sum_array_0_20_port, 
                           A(19) => sum_array_0_19_port, A(18) => 
                           sum_array_0_18_port, A(17) => sum_array_0_17_port, 
                           A(16) => sum_array_0_16_port, A(15) => 
                           sum_array_0_15_port, A(14) => sum_array_0_14_port, 
                           A(13) => sum_array_0_13_port, A(12) => 
                           sum_array_0_12_port, A(11) => sum_array_0_11_port, 
                           A(10) => sum_array_0_10_port, A(9) => 
                           sum_array_0_9_port, A(8) => sum_array_0_8_port, A(7)
                           => sum_array_0_7_port, A(6) => sum_array_0_6_port, 
                           A(5) => sum_array_0_5_port, A(4) => 
                           sum_array_0_4_port, A(3) => sum_array_0_3_port, A(2)
                           => sum_array_0_2_port, A(1) => sum_array_0_1_port, 
                           A(0) => sum_array_0_0_port, B(31) => 
                           cout_array_0_31_port, B(30) => cout_array_0_30_port,
                           B(29) => cout_array_0_29_port, B(28) => 
                           cout_array_0_28_port, B(27) => cout_array_0_27_port,
                           B(26) => cout_array_0_26_port, B(25) => 
                           cout_array_0_25_port, B(24) => cout_array_0_24_port,
                           B(23) => cout_array_0_23_port, B(22) => 
                           cout_array_0_22_port, B(21) => cout_array_0_21_port,
                           B(20) => cout_array_0_20_port, B(19) => 
                           cout_array_0_19_port, B(18) => cout_array_0_18_port,
                           B(17) => cout_array_0_17_port, B(16) => 
                           cout_array_0_16_port, B(15) => cout_array_0_15_port,
                           B(14) => cout_array_0_14_port, B(13) => 
                           cout_array_0_13_port, B(12) => cout_array_0_12_port,
                           B(11) => cout_array_0_11_port, B(10) => 
                           cout_array_0_10_port, B(9) => cout_array_0_9_port, 
                           B(8) => cout_array_0_8_port, B(7) => 
                           cout_array_0_7_port, B(6) => cout_array_0_6_port, 
                           B(5) => cout_array_0_5_port, B(4) => 
                           cout_array_0_4_port, B(3) => cout_array_0_3_port, 
                           B(2) => cout_array_0_2_port, B(1) => 
                           cout_array_0_1_port, B(0) => cout_array_0_0_port, 
                           C(31) => sum_array_1_31_port, C(30) => 
                           sum_array_1_30_port, C(29) => sum_array_1_29_port, 
                           C(28) => sum_array_1_28_port, C(27) => 
                           sum_array_1_27_port, C(26) => sum_array_1_26_port, 
                           C(25) => sum_array_1_25_port, C(24) => 
                           sum_array_1_24_port, C(23) => sum_array_1_23_port, 
                           C(22) => sum_array_1_22_port, C(21) => 
                           sum_array_1_21_port, C(20) => sum_array_1_20_port, 
                           C(19) => sum_array_1_19_port, C(18) => 
                           sum_array_1_18_port, C(17) => sum_array_1_17_port, 
                           C(16) => sum_array_1_16_port, C(15) => 
                           sum_array_1_15_port, C(14) => sum_array_1_14_port, 
                           C(13) => sum_array_1_13_port, C(12) => 
                           sum_array_1_12_port, C(11) => sum_array_1_11_port, 
                           C(10) => sum_array_1_10_port, C(9) => 
                           sum_array_1_9_port, C(8) => sum_array_1_8_port, C(7)
                           => sum_array_1_7_port, C(6) => sum_array_1_6_port, 
                           C(5) => sum_array_1_5_port, C(4) => 
                           sum_array_1_4_port, C(3) => sum_array_1_3_port, C(2)
                           => sum_array_1_2_port, C(1) => sum_array_1_1_port, 
                           C(0) => sum_array_1_0_port, S(31) => 
                           sum_array_2_31_port, S(30) => sum_array_2_30_port, 
                           S(29) => sum_array_2_29_port, S(28) => 
                           sum_array_2_28_port, S(27) => sum_array_2_27_port, 
                           S(26) => sum_array_2_26_port, S(25) => 
                           sum_array_2_25_port, S(24) => sum_array_2_24_port, 
                           S(23) => sum_array_2_23_port, S(22) => 
                           sum_array_2_22_port, S(21) => sum_array_2_21_port, 
                           S(20) => sum_array_2_20_port, S(19) => 
                           sum_array_2_19_port, S(18) => sum_array_2_18_port, 
                           S(17) => sum_array_2_17_port, S(16) => 
                           sum_array_2_16_port, S(15) => sum_array_2_15_port, 
                           S(14) => sum_array_2_14_port, S(13) => 
                           sum_array_2_13_port, S(12) => sum_array_2_12_port, 
                           S(11) => sum_array_2_11_port, S(10) => 
                           sum_array_2_10_port, S(9) => sum_array_2_9_port, 
                           S(8) => sum_array_2_8_port, S(7) => 
                           sum_array_2_7_port, S(6) => sum_array_2_6_port, S(5)
                           => sum_array_2_5_port, S(4) => sum_array_2_4_port, 
                           S(3) => sum_array_2_3_port, S(2) => 
                           sum_array_2_2_port, S(1) => sum_array_2_1_port, S(0)
                           => sum_array_2_0_port, Cout(31) => 
                           cout_array_2_31_port, Cout(30) => 
                           cout_array_2_30_port, Cout(29) => 
                           cout_array_2_29_port, Cout(28) => 
                           cout_array_2_28_port, Cout(27) => 
                           cout_array_2_27_port, Cout(26) => 
                           cout_array_2_26_port, Cout(25) => 
                           cout_array_2_25_port, Cout(24) => 
                           cout_array_2_24_port, Cout(23) => 
                           cout_array_2_23_port, Cout(22) => 
                           cout_array_2_22_port, Cout(21) => 
                           cout_array_2_21_port, Cout(20) => 
                           cout_array_2_20_port, Cout(19) => 
                           cout_array_2_19_port, Cout(18) => 
                           cout_array_2_18_port, Cout(17) => 
                           cout_array_2_17_port, Cout(16) => 
                           cout_array_2_16_port, Cout(15) => 
                           cout_array_2_15_port, Cout(14) => 
                           cout_array_2_14_port, Cout(13) => 
                           cout_array_2_13_port, Cout(12) => 
                           cout_array_2_12_port, Cout(11) => 
                           cout_array_2_11_port, Cout(10) => 
                           cout_array_2_10_port, Cout(9) => cout_array_2_9_port
                           , Cout(8) => cout_array_2_8_port, Cout(7) => 
                           cout_array_2_7_port, Cout(6) => cout_array_2_6_port,
                           Cout(5) => cout_array_2_5_port, Cout(4) => 
                           cout_array_2_4_port, Cout(3) => cout_array_2_3_port,
                           Cout(2) => cout_array_2_2_port, Cout(1) => 
                           cout_array_2_1_port, Cout(0) => net59832);
   Add2IIL : CSA_Nbits32_3 port map( A(31) => cout_array_1_31_port, A(30) => 
                           cout_array_1_30_port, A(29) => cout_array_1_29_port,
                           A(28) => cout_array_1_28_port, A(27) => 
                           cout_array_1_27_port, A(26) => cout_array_1_26_port,
                           A(25) => cout_array_1_25_port, A(24) => 
                           cout_array_1_24_port, A(23) => cout_array_1_23_port,
                           A(22) => cout_array_1_22_port, A(21) => 
                           cout_array_1_21_port, A(20) => cout_array_1_20_port,
                           A(19) => cout_array_1_19_port, A(18) => 
                           cout_array_1_18_port, A(17) => cout_array_1_17_port,
                           A(16) => cout_array_1_16_port, A(15) => 
                           cout_array_1_15_port, A(14) => cout_array_1_14_port,
                           A(13) => cout_array_1_13_port, A(12) => 
                           cout_array_1_12_port, A(11) => cout_array_1_11_port,
                           A(10) => cout_array_1_10_port, A(9) => 
                           cout_array_1_9_port, A(8) => cout_array_1_8_port, 
                           A(7) => cout_array_1_7_port, A(6) => 
                           cout_array_1_6_port, A(5) => cout_array_1_5_port, 
                           A(4) => cout_array_1_4_port, A(3) => 
                           cout_array_1_3_port, A(2) => cout_array_1_2_port, 
                           A(1) => cout_array_1_1_port, A(0) => 
                           cout_array_1_0_port, B(31) => outmux_6_31_port, 
                           B(30) => outmux_6_30_port, B(29) => outmux_6_29_port
                           , B(28) => outmux_6_28_port, B(27) => 
                           outmux_6_27_port, B(26) => outmux_6_26_port, B(25) 
                           => outmux_6_25_port, B(24) => outmux_6_24_port, 
                           B(23) => outmux_6_23_port, B(22) => outmux_6_22_port
                           , B(21) => outmux_6_21_port, B(20) => 
                           outmux_6_20_port, B(19) => outmux_6_19_port, B(18) 
                           => outmux_6_18_port, B(17) => outmux_6_17_port, 
                           B(16) => outmux_6_16_port, B(15) => outmux_6_15_port
                           , B(14) => outmux_6_14_port, B(13) => 
                           outmux_6_13_port, B(12) => outmux_6_12_port, B(11) 
                           => outmux_6_11_port, B(10) => outmux_6_10_port, B(9)
                           => outmux_6_9_port, B(8) => outmux_6_8_port, B(7) =>
                           outmux_6_7_port, B(6) => outmux_6_6_port, B(5) => 
                           outmux_6_5_port, B(4) => outmux_6_4_port, B(3) => 
                           outmux_6_3_port, B(2) => outmux_6_2_port, B(1) => 
                           outmux_6_1_port, B(0) => outmux_6_0_port, C(31) => 
                           outmux_7_31_port, C(30) => outmux_7_30_port, C(29) 
                           => outmux_7_29_port, C(28) => outmux_7_28_port, 
                           C(27) => outmux_7_27_port, C(26) => outmux_7_26_port
                           , C(25) => outmux_7_25_port, C(24) => 
                           outmux_7_24_port, C(23) => outmux_7_23_port, C(22) 
                           => outmux_7_22_port, C(21) => outmux_7_21_port, 
                           C(20) => outmux_7_20_port, C(19) => outmux_7_19_port
                           , C(18) => outmux_7_18_port, C(17) => 
                           outmux_7_17_port, C(16) => outmux_7_16_port, C(15) 
                           => outmux_7_15_port, C(14) => outmux_7_14_port, 
                           C(13) => outmux_7_13_port, C(12) => outmux_7_12_port
                           , C(11) => outmux_7_11_port, C(10) => 
                           outmux_7_10_port, C(9) => outmux_7_9_port, C(8) => 
                           outmux_7_8_port, C(7) => outmux_7_7_port, C(6) => 
                           outmux_7_6_port, C(5) => outmux_7_5_port, C(4) => 
                           outmux_7_4_port, C(3) => outmux_7_3_port, C(2) => 
                           outmux_7_2_port, C(1) => outmux_7_1_port, C(0) => 
                           outmux_7_0_port, S(31) => sum_array_3_31_port, S(30)
                           => sum_array_3_30_port, S(29) => sum_array_3_29_port
                           , S(28) => sum_array_3_28_port, S(27) => 
                           sum_array_3_27_port, S(26) => sum_array_3_26_port, 
                           S(25) => sum_array_3_25_port, S(24) => 
                           sum_array_3_24_port, S(23) => sum_array_3_23_port, 
                           S(22) => sum_array_3_22_port, S(21) => 
                           sum_array_3_21_port, S(20) => sum_array_3_20_port, 
                           S(19) => sum_array_3_19_port, S(18) => 
                           sum_array_3_18_port, S(17) => sum_array_3_17_port, 
                           S(16) => sum_array_3_16_port, S(15) => 
                           sum_array_3_15_port, S(14) => sum_array_3_14_port, 
                           S(13) => sum_array_3_13_port, S(12) => 
                           sum_array_3_12_port, S(11) => sum_array_3_11_port, 
                           S(10) => sum_array_3_10_port, S(9) => 
                           sum_array_3_9_port, S(8) => sum_array_3_8_port, S(7)
                           => sum_array_3_7_port, S(6) => sum_array_3_6_port, 
                           S(5) => sum_array_3_5_port, S(4) => 
                           sum_array_3_4_port, S(3) => sum_array_3_3_port, S(2)
                           => sum_array_3_2_port, S(1) => sum_array_3_1_port, 
                           S(0) => sum_array_3_0_port, Cout(31) => 
                           cout_array_3_31_port, Cout(30) => 
                           cout_array_3_30_port, Cout(29) => 
                           cout_array_3_29_port, Cout(28) => 
                           cout_array_3_28_port, Cout(27) => 
                           cout_array_3_27_port, Cout(26) => 
                           cout_array_3_26_port, Cout(25) => 
                           cout_array_3_25_port, Cout(24) => 
                           cout_array_3_24_port, Cout(23) => 
                           cout_array_3_23_port, Cout(22) => 
                           cout_array_3_22_port, Cout(21) => 
                           cout_array_3_21_port, Cout(20) => 
                           cout_array_3_20_port, Cout(19) => 
                           cout_array_3_19_port, Cout(18) => 
                           cout_array_3_18_port, Cout(17) => 
                           cout_array_3_17_port, Cout(16) => 
                           cout_array_3_16_port, Cout(15) => 
                           cout_array_3_15_port, Cout(14) => 
                           cout_array_3_14_port, Cout(13) => 
                           cout_array_3_13_port, Cout(12) => 
                           cout_array_3_12_port, Cout(11) => 
                           cout_array_3_11_port, Cout(10) => 
                           cout_array_3_10_port, Cout(9) => cout_array_3_9_port
                           , Cout(8) => cout_array_3_8_port, Cout(7) => 
                           cout_array_3_7_port, Cout(6) => cout_array_3_6_port,
                           Cout(5) => cout_array_3_5_port, Cout(4) => 
                           cout_array_3_4_port, Cout(3) => cout_array_3_3_port,
                           Cout(2) => cout_array_3_2_port, Cout(1) => 
                           cout_array_3_1_port, Cout(0) => net59831);
   Add1IIIL : CSA_Nbits32_2 port map( A(31) => sum_array_2_31_port, A(30) => 
                           sum_array_2_30_port, A(29) => sum_array_2_29_port, 
                           A(28) => sum_array_2_28_port, A(27) => 
                           sum_array_2_27_port, A(26) => sum_array_2_26_port, 
                           A(25) => sum_array_2_25_port, A(24) => 
                           sum_array_2_24_port, A(23) => sum_array_2_23_port, 
                           A(22) => sum_array_2_22_port, A(21) => 
                           sum_array_2_21_port, A(20) => sum_array_2_20_port, 
                           A(19) => sum_array_2_19_port, A(18) => 
                           sum_array_2_18_port, A(17) => sum_array_2_17_port, 
                           A(16) => sum_array_2_16_port, A(15) => 
                           sum_array_2_15_port, A(14) => sum_array_2_14_port, 
                           A(13) => sum_array_2_13_port, A(12) => 
                           sum_array_2_12_port, A(11) => sum_array_2_11_port, 
                           A(10) => sum_array_2_10_port, A(9) => 
                           sum_array_2_9_port, A(8) => sum_array_2_8_port, A(7)
                           => sum_array_2_7_port, A(6) => sum_array_2_6_port, 
                           A(5) => sum_array_2_5_port, A(4) => 
                           sum_array_2_4_port, A(3) => sum_array_2_3_port, A(2)
                           => sum_array_2_2_port, A(1) => sum_array_2_1_port, 
                           A(0) => sum_array_2_0_port, B(31) => 
                           cout_array_2_31_port, B(30) => cout_array_2_30_port,
                           B(29) => cout_array_2_29_port, B(28) => 
                           cout_array_2_28_port, B(27) => cout_array_2_27_port,
                           B(26) => cout_array_2_26_port, B(25) => 
                           cout_array_2_25_port, B(24) => cout_array_2_24_port,
                           B(23) => cout_array_2_23_port, B(22) => 
                           cout_array_2_22_port, B(21) => cout_array_2_21_port,
                           B(20) => cout_array_2_20_port, B(19) => 
                           cout_array_2_19_port, B(18) => cout_array_2_18_port,
                           B(17) => cout_array_2_17_port, B(16) => 
                           cout_array_2_16_port, B(15) => cout_array_2_15_port,
                           B(14) => cout_array_2_14_port, B(13) => 
                           cout_array_2_13_port, B(12) => cout_array_2_12_port,
                           B(11) => cout_array_2_11_port, B(10) => 
                           cout_array_2_10_port, B(9) => cout_array_2_9_port, 
                           B(8) => cout_array_2_8_port, B(7) => 
                           cout_array_2_7_port, B(6) => cout_array_2_6_port, 
                           B(5) => cout_array_2_5_port, B(4) => 
                           cout_array_2_4_port, B(3) => cout_array_2_3_port, 
                           B(2) => cout_array_2_2_port, B(1) => 
                           cout_array_2_1_port, B(0) => cout_array_2_0_port, 
                           C(31) => sum_array_3_31_port, C(30) => 
                           sum_array_3_30_port, C(29) => sum_array_3_29_port, 
                           C(28) => sum_array_3_28_port, C(27) => 
                           sum_array_3_27_port, C(26) => sum_array_3_26_port, 
                           C(25) => sum_array_3_25_port, C(24) => 
                           sum_array_3_24_port, C(23) => sum_array_3_23_port, 
                           C(22) => sum_array_3_22_port, C(21) => 
                           sum_array_3_21_port, C(20) => sum_array_3_20_port, 
                           C(19) => sum_array_3_19_port, C(18) => 
                           sum_array_3_18_port, C(17) => sum_array_3_17_port, 
                           C(16) => sum_array_3_16_port, C(15) => 
                           sum_array_3_15_port, C(14) => sum_array_3_14_port, 
                           C(13) => sum_array_3_13_port, C(12) => 
                           sum_array_3_12_port, C(11) => sum_array_3_11_port, 
                           C(10) => sum_array_3_10_port, C(9) => 
                           sum_array_3_9_port, C(8) => sum_array_3_8_port, C(7)
                           => sum_array_3_7_port, C(6) => sum_array_3_6_port, 
                           C(5) => sum_array_3_5_port, C(4) => 
                           sum_array_3_4_port, C(3) => sum_array_3_3_port, C(2)
                           => sum_array_3_2_port, C(1) => sum_array_3_1_port, 
                           C(0) => sum_array_3_0_port, S(31) => 
                           sum_array_4_31_port, S(30) => sum_array_4_30_port, 
                           S(29) => sum_array_4_29_port, S(28) => 
                           sum_array_4_28_port, S(27) => sum_array_4_27_port, 
                           S(26) => sum_array_4_26_port, S(25) => 
                           sum_array_4_25_port, S(24) => sum_array_4_24_port, 
                           S(23) => sum_array_4_23_port, S(22) => 
                           sum_array_4_22_port, S(21) => sum_array_4_21_port, 
                           S(20) => sum_array_4_20_port, S(19) => 
                           sum_array_4_19_port, S(18) => sum_array_4_18_port, 
                           S(17) => sum_array_4_17_port, S(16) => 
                           sum_array_4_16_port, S(15) => sum_array_4_15_port, 
                           S(14) => sum_array_4_14_port, S(13) => 
                           sum_array_4_13_port, S(12) => sum_array_4_12_port, 
                           S(11) => sum_array_4_11_port, S(10) => 
                           sum_array_4_10_port, S(9) => sum_array_4_9_port, 
                           S(8) => sum_array_4_8_port, S(7) => 
                           sum_array_4_7_port, S(6) => sum_array_4_6_port, S(5)
                           => sum_array_4_5_port, S(4) => sum_array_4_4_port, 
                           S(3) => sum_array_4_3_port, S(2) => 
                           sum_array_4_2_port, S(1) => sum_array_4_1_port, S(0)
                           => sum_array_4_0_port, Cout(31) => 
                           cout_array_4_31_port, Cout(30) => 
                           cout_array_4_30_port, Cout(29) => 
                           cout_array_4_29_port, Cout(28) => 
                           cout_array_4_28_port, Cout(27) => 
                           cout_array_4_27_port, Cout(26) => 
                           cout_array_4_26_port, Cout(25) => 
                           cout_array_4_25_port, Cout(24) => 
                           cout_array_4_24_port, Cout(23) => 
                           cout_array_4_23_port, Cout(22) => 
                           cout_array_4_22_port, Cout(21) => 
                           cout_array_4_21_port, Cout(20) => 
                           cout_array_4_20_port, Cout(19) => 
                           cout_array_4_19_port, Cout(18) => 
                           cout_array_4_18_port, Cout(17) => 
                           cout_array_4_17_port, Cout(16) => 
                           cout_array_4_16_port, Cout(15) => 
                           cout_array_4_15_port, Cout(14) => 
                           cout_array_4_14_port, Cout(13) => 
                           cout_array_4_13_port, Cout(12) => 
                           cout_array_4_12_port, Cout(11) => 
                           cout_array_4_11_port, Cout(10) => 
                           cout_array_4_10_port, Cout(9) => cout_array_4_9_port
                           , Cout(8) => cout_array_4_8_port, Cout(7) => 
                           cout_array_4_7_port, Cout(6) => cout_array_4_6_port,
                           Cout(5) => cout_array_4_5_port, Cout(4) => 
                           cout_array_4_4_port, Cout(3) => cout_array_4_3_port,
                           Cout(2) => cout_array_4_2_port, Cout(1) => 
                           cout_array_4_1_port, Cout(0) => net59830);
   AddRCA : CSA_Nbits32_1 port map( A(31) => sum_array_4_31_port, A(30) => 
                           sum_array_4_30_port, A(29) => sum_array_4_29_port, 
                           A(28) => sum_array_4_28_port, A(27) => 
                           sum_array_4_27_port, A(26) => sum_array_4_26_port, 
                           A(25) => sum_array_4_25_port, A(24) => 
                           sum_array_4_24_port, A(23) => sum_array_4_23_port, 
                           A(22) => sum_array_4_22_port, A(21) => 
                           sum_array_4_21_port, A(20) => sum_array_4_20_port, 
                           A(19) => sum_array_4_19_port, A(18) => 
                           sum_array_4_18_port, A(17) => sum_array_4_17_port, 
                           A(16) => sum_array_4_16_port, A(15) => 
                           sum_array_4_15_port, A(14) => sum_array_4_14_port, 
                           A(13) => sum_array_4_13_port, A(12) => 
                           sum_array_4_12_port, A(11) => sum_array_4_11_port, 
                           A(10) => sum_array_4_10_port, A(9) => 
                           sum_array_4_9_port, A(8) => sum_array_4_8_port, A(7)
                           => sum_array_4_7_port, A(6) => sum_array_4_6_port, 
                           A(5) => sum_array_4_5_port, A(4) => 
                           sum_array_4_4_port, A(3) => sum_array_4_3_port, A(2)
                           => sum_array_4_2_port, A(1) => sum_array_4_1_port, 
                           A(0) => sum_array_4_0_port, B(31) => 
                           cout_array_4_31_port, B(30) => cout_array_4_30_port,
                           B(29) => cout_array_4_29_port, B(28) => 
                           cout_array_4_28_port, B(27) => cout_array_4_27_port,
                           B(26) => cout_array_4_26_port, B(25) => 
                           cout_array_4_25_port, B(24) => cout_array_4_24_port,
                           B(23) => cout_array_4_23_port, B(22) => 
                           cout_array_4_22_port, B(21) => cout_array_4_21_port,
                           B(20) => cout_array_4_20_port, B(19) => 
                           cout_array_4_19_port, B(18) => cout_array_4_18_port,
                           B(17) => cout_array_4_17_port, B(16) => 
                           cout_array_4_16_port, B(15) => cout_array_4_15_port,
                           B(14) => cout_array_4_14_port, B(13) => 
                           cout_array_4_13_port, B(12) => cout_array_4_12_port,
                           B(11) => cout_array_4_11_port, B(10) => 
                           cout_array_4_10_port, B(9) => cout_array_4_9_port, 
                           B(8) => cout_array_4_8_port, B(7) => 
                           cout_array_4_7_port, B(6) => cout_array_4_6_port, 
                           B(5) => cout_array_4_5_port, B(4) => 
                           cout_array_4_4_port, B(3) => cout_array_4_3_port, 
                           B(2) => cout_array_4_2_port, B(1) => 
                           cout_array_4_1_port, B(0) => cout_array_4_0_port, 
                           C(31) => cout_array_3_31_port, C(30) => 
                           cout_array_3_30_port, C(29) => cout_array_3_29_port,
                           C(28) => cout_array_3_28_port, C(27) => 
                           cout_array_3_27_port, C(26) => cout_array_3_26_port,
                           C(25) => cout_array_3_25_port, C(24) => 
                           cout_array_3_24_port, C(23) => cout_array_3_23_port,
                           C(22) => cout_array_3_22_port, C(21) => 
                           cout_array_3_21_port, C(20) => cout_array_3_20_port,
                           C(19) => cout_array_3_19_port, C(18) => 
                           cout_array_3_18_port, C(17) => cout_array_3_17_port,
                           C(16) => cout_array_3_16_port, C(15) => 
                           cout_array_3_15_port, C(14) => cout_array_3_14_port,
                           C(13) => cout_array_3_13_port, C(12) => 
                           cout_array_3_12_port, C(11) => cout_array_3_11_port,
                           C(10) => cout_array_3_10_port, C(9) => 
                           cout_array_3_9_port, C(8) => cout_array_3_8_port, 
                           C(7) => cout_array_3_7_port, C(6) => 
                           cout_array_3_6_port, C(5) => cout_array_3_5_port, 
                           C(4) => cout_array_3_4_port, C(3) => 
                           cout_array_3_3_port, C(2) => cout_array_3_2_port, 
                           C(1) => cout_array_3_1_port, C(0) => 
                           cout_array_3_0_port, S(31) => sum_array_5_31_port, 
                           S(30) => sum_array_5_30_port, S(29) => 
                           sum_array_5_29_port, S(28) => sum_array_5_28_port, 
                           S(27) => sum_array_5_27_port, S(26) => 
                           sum_array_5_26_port, S(25) => sum_array_5_25_port, 
                           S(24) => sum_array_5_24_port, S(23) => 
                           sum_array_5_23_port, S(22) => sum_array_5_22_port, 
                           S(21) => sum_array_5_21_port, S(20) => 
                           sum_array_5_20_port, S(19) => sum_array_5_19_port, 
                           S(18) => sum_array_5_18_port, S(17) => 
                           sum_array_5_17_port, S(16) => sum_array_5_16_port, 
                           S(15) => sum_array_5_15_port, S(14) => 
                           sum_array_5_14_port, S(13) => sum_array_5_13_port, 
                           S(12) => sum_array_5_12_port, S(11) => 
                           sum_array_5_11_port, S(10) => sum_array_5_10_port, 
                           S(9) => sum_array_5_9_port, S(8) => 
                           sum_array_5_8_port, S(7) => sum_array_5_7_port, S(6)
                           => sum_array_5_6_port, S(5) => sum_array_5_5_port, 
                           S(4) => sum_array_5_4_port, S(3) => 
                           sum_array_5_3_port, S(2) => sum_array_5_2_port, S(1)
                           => sum_array_5_1_port, S(0) => sum_array_5_0_port, 
                           Cout(31) => cout_array_5_31_port, Cout(30) => 
                           cout_array_5_30_port, Cout(29) => 
                           cout_array_5_29_port, Cout(28) => 
                           cout_array_5_28_port, Cout(27) => 
                           cout_array_5_27_port, Cout(26) => 
                           cout_array_5_26_port, Cout(25) => 
                           cout_array_5_25_port, Cout(24) => 
                           cout_array_5_24_port, Cout(23) => 
                           cout_array_5_23_port, Cout(22) => 
                           cout_array_5_22_port, Cout(21) => 
                           cout_array_5_21_port, Cout(20) => 
                           cout_array_5_20_port, Cout(19) => 
                           cout_array_5_19_port, Cout(18) => 
                           cout_array_5_18_port, Cout(17) => 
                           cout_array_5_17_port, Cout(16) => 
                           cout_array_5_16_port, Cout(15) => 
                           cout_array_5_15_port, Cout(14) => 
                           cout_array_5_14_port, Cout(13) => 
                           cout_array_5_13_port, Cout(12) => 
                           cout_array_5_12_port, Cout(11) => 
                           cout_array_5_11_port, Cout(10) => 
                           cout_array_5_10_port, Cout(9) => cout_array_5_9_port
                           , Cout(8) => cout_array_5_8_port, Cout(7) => 
                           cout_array_5_7_port, Cout(6) => cout_array_5_6_port,
                           Cout(5) => cout_array_5_5_port, Cout(4) => 
                           cout_array_5_4_port, Cout(3) => cout_array_5_3_port,
                           Cout(2) => cout_array_5_2_port, Cout(1) => 
                           cout_array_5_1_port, Cout(0) => net59829);
   P4adder : cla_adder_N32_1 port map( A(31) => sum_array_5_31_port, A(30) => 
                           sum_array_5_30_port, A(29) => sum_array_5_29_port, 
                           A(28) => sum_array_5_28_port, A(27) => 
                           sum_array_5_27_port, A(26) => sum_array_5_26_port, 
                           A(25) => sum_array_5_25_port, A(24) => 
                           sum_array_5_24_port, A(23) => sum_array_5_23_port, 
                           A(22) => sum_array_5_22_port, A(21) => 
                           sum_array_5_21_port, A(20) => sum_array_5_20_port, 
                           A(19) => sum_array_5_19_port, A(18) => 
                           sum_array_5_18_port, A(17) => sum_array_5_17_port, 
                           A(16) => sum_array_5_16_port, A(15) => 
                           sum_array_5_15_port, A(14) => sum_array_5_14_port, 
                           A(13) => sum_array_5_13_port, A(12) => 
                           sum_array_5_12_port, A(11) => sum_array_5_11_port, 
                           A(10) => sum_array_5_10_port, A(9) => 
                           sum_array_5_9_port, A(8) => sum_array_5_8_port, A(7)
                           => sum_array_5_7_port, A(6) => sum_array_5_6_port, 
                           A(5) => sum_array_5_5_port, A(4) => 
                           sum_array_5_4_port, A(3) => sum_array_5_3_port, A(2)
                           => sum_array_5_2_port, A(1) => sum_array_5_1_port, 
                           A(0) => sum_array_5_0_port, B(31) => 
                           cout_array_5_31_port, B(30) => cout_array_5_30_port,
                           B(29) => cout_array_5_29_port, B(28) => 
                           cout_array_5_28_port, B(27) => cout_array_5_27_port,
                           B(26) => cout_array_5_26_port, B(25) => 
                           cout_array_5_25_port, B(24) => cout_array_5_24_port,
                           B(23) => cout_array_5_23_port, B(22) => 
                           cout_array_5_22_port, B(21) => cout_array_5_21_port,
                           B(20) => cout_array_5_20_port, B(19) => 
                           cout_array_5_19_port, B(18) => cout_array_5_18_port,
                           B(17) => cout_array_5_17_port, B(16) => 
                           cout_array_5_16_port, B(15) => cout_array_5_15_port,
                           B(14) => cout_array_5_14_port, B(13) => 
                           cout_array_5_13_port, B(12) => cout_array_5_12_port,
                           B(11) => cout_array_5_11_port, B(10) => 
                           cout_array_5_10_port, B(9) => cout_array_5_9_port, 
                           B(8) => cout_array_5_8_port, B(7) => 
                           cout_array_5_7_port, B(6) => cout_array_5_6_port, 
                           B(5) => cout_array_5_5_port, B(4) => 
                           cout_array_5_4_port, B(3) => cout_array_5_3_port, 
                           B(2) => cout_array_5_2_port, B(1) => 
                           cout_array_5_1_port, B(0) => cout_array_5_0_port, Ci
                           => X_Logic0_port, Cout => net6197, Sum(31) => Y(31),
                           Sum(30) => Y(30), Sum(29) => Y(29), Sum(28) => Y(28)
                           , Sum(27) => Y(27), Sum(26) => Y(26), Sum(25) => 
                           Y(25), Sum(24) => Y(24), Sum(23) => Y(23), Sum(22) 
                           => Y(22), Sum(21) => Y(21), Sum(20) => Y(20), 
                           Sum(19) => Y(19), Sum(18) => Y(18), Sum(17) => Y(17)
                           , Sum(16) => Y(16), Sum(15) => Y(15), Sum(14) => 
                           Y(14), Sum(13) => Y(13), Sum(12) => Y(12), Sum(11) 
                           => Y(11), Sum(10) => Y(10), Sum(9) => Y(9), Sum(8) 
                           => Y(8), Sum(7) => Y(7), Sum(6) => Y(6), Sum(5) => 
                           Y(5), Sum(4) => Y(4), Sum(3) => Y(3), Sum(2) => Y(2)
                           , Sum(1) => Y(1), Sum(0) => Y(0));
   cout_array_1_0_port <= '0';
   cout_array_2_0_port <= '0';
   cout_array_3_0_port <= '0';
   cout_array_4_0_port <= '0';
   cout_array_5_0_port <= '0';
   cout_array_0_0_port <= '0';
   muxInE_7_0_port <= '0';
   muxInE_7_1_port <= '0';
   muxInE_7_2_port <= '0';
   muxInE_7_3_port <= '0';
   muxInE_7_4_port <= '0';
   muxInE_7_5_port <= '0';
   muxInE_7_6_port <= '0';
   muxInE_7_7_port <= '0';
   muxInE_7_8_port <= '0';
   muxInE_7_9_port <= '0';
   muxInE_7_10_port <= '0';
   muxInE_7_11_port <= '0';
   muxInE_7_12_port <= '0';
   muxInE_7_13_port <= '0';
   muxInE_7_14_port <= '0';
   muxInD_7_0_port <= '0';
   muxInD_7_1_port <= '0';
   muxInD_7_2_port <= '0';
   muxInD_7_3_port <= '0';
   muxInD_7_4_port <= '0';
   muxInD_7_5_port <= '0';
   muxInD_7_6_port <= '0';
   muxInD_7_7_port <= '0';
   muxInD_7_8_port <= '0';
   muxInD_7_9_port <= '0';
   muxInD_7_10_port <= '0';
   muxInD_7_11_port <= '0';
   muxInD_7_12_port <= '0';
   muxInD_7_13_port <= '0';
   muxInD_7_14_port <= '0';
   muxInC_7_0_port <= '0';
   muxInC_7_1_port <= '0';
   muxInC_7_2_port <= '0';
   muxInC_7_3_port <= '0';
   muxInC_7_4_port <= '0';
   muxInC_7_5_port <= '0';
   muxInC_7_6_port <= '0';
   muxInC_7_7_port <= '0';
   muxInC_7_8_port <= '0';
   muxInC_7_9_port <= '0';
   muxInC_7_10_port <= '0';
   muxInC_7_11_port <= '0';
   muxInC_7_12_port <= '0';
   muxInC_7_13_port <= '0';
   muxInB_7_0_port <= '0';
   muxInB_7_1_port <= '0';
   muxInB_7_2_port <= '0';
   muxInB_7_3_port <= '0';
   muxInB_7_4_port <= '0';
   muxInB_7_5_port <= '0';
   muxInB_7_6_port <= '0';
   muxInB_7_7_port <= '0';
   muxInB_7_8_port <= '0';
   muxInB_7_9_port <= '0';
   muxInB_7_10_port <= '0';
   muxInB_7_11_port <= '0';
   muxInB_7_12_port <= '0';
   muxInB_7_13_port <= '0';
   muxInE_6_0_port <= '0';
   muxInE_6_1_port <= '0';
   muxInE_6_2_port <= '0';
   muxInE_6_3_port <= '0';
   muxInE_6_4_port <= '0';
   muxInE_6_5_port <= '0';
   muxInE_6_6_port <= '0';
   muxInE_6_7_port <= '0';
   muxInE_6_8_port <= '0';
   muxInE_6_9_port <= '0';
   muxInE_6_10_port <= '0';
   muxInE_6_11_port <= '0';
   muxInE_6_12_port <= '0';
   muxInD_6_0_port <= '0';
   muxInD_6_1_port <= '0';
   muxInD_6_2_port <= '0';
   muxInD_6_3_port <= '0';
   muxInD_6_4_port <= '0';
   muxInD_6_5_port <= '0';
   muxInD_6_6_port <= '0';
   muxInD_6_7_port <= '0';
   muxInD_6_8_port <= '0';
   muxInD_6_9_port <= '0';
   muxInD_6_10_port <= '0';
   muxInD_6_11_port <= '0';
   muxInD_6_12_port <= '0';
   muxInC_6_0_port <= '0';
   muxInC_6_1_port <= '0';
   muxInC_6_2_port <= '0';
   muxInC_6_3_port <= '0';
   muxInC_6_4_port <= '0';
   muxInC_6_5_port <= '0';
   muxInC_6_6_port <= '0';
   muxInC_6_7_port <= '0';
   muxInC_6_8_port <= '0';
   muxInC_6_9_port <= '0';
   muxInC_6_10_port <= '0';
   muxInC_6_11_port <= '0';
   muxInB_6_0_port <= '0';
   muxInB_6_1_port <= '0';
   muxInB_6_2_port <= '0';
   muxInB_6_3_port <= '0';
   muxInB_6_4_port <= '0';
   muxInB_6_5_port <= '0';
   muxInB_6_6_port <= '0';
   muxInB_6_7_port <= '0';
   muxInB_6_8_port <= '0';
   muxInB_6_9_port <= '0';
   muxInB_6_10_port <= '0';
   muxInB_6_11_port <= '0';
   muxInE_5_0_port <= '0';
   muxInE_5_1_port <= '0';
   muxInE_5_2_port <= '0';
   muxInE_5_3_port <= '0';
   muxInE_5_4_port <= '0';
   muxInE_5_5_port <= '0';
   muxInE_5_6_port <= '0';
   muxInE_5_7_port <= '0';
   muxInE_5_8_port <= '0';
   muxInE_5_9_port <= '0';
   muxInE_5_10_port <= '0';
   muxInD_5_0_port <= '0';
   muxInD_5_1_port <= '0';
   muxInD_5_2_port <= '0';
   muxInD_5_3_port <= '0';
   muxInD_5_4_port <= '0';
   muxInD_5_5_port <= '0';
   muxInD_5_6_port <= '0';
   muxInD_5_7_port <= '0';
   muxInD_5_8_port <= '0';
   muxInD_5_9_port <= '0';
   muxInD_5_10_port <= '0';
   muxInC_5_0_port <= '0';
   muxInC_5_1_port <= '0';
   muxInC_5_2_port <= '0';
   muxInC_5_3_port <= '0';
   muxInC_5_4_port <= '0';
   muxInC_5_5_port <= '0';
   muxInC_5_6_port <= '0';
   muxInC_5_7_port <= '0';
   muxInC_5_8_port <= '0';
   muxInC_5_9_port <= '0';
   muxInB_5_0_port <= '0';
   muxInB_5_1_port <= '0';
   muxInB_5_2_port <= '0';
   muxInB_5_3_port <= '0';
   muxInB_5_4_port <= '0';
   muxInB_5_5_port <= '0';
   muxInB_5_6_port <= '0';
   muxInB_5_7_port <= '0';
   muxInB_5_8_port <= '0';
   muxInB_5_9_port <= '0';
   muxInE_4_0_port <= '0';
   muxInE_4_1_port <= '0';
   muxInE_4_2_port <= '0';
   muxInE_4_3_port <= '0';
   muxInE_4_4_port <= '0';
   muxInE_4_5_port <= '0';
   muxInE_4_6_port <= '0';
   muxInE_4_7_port <= '0';
   muxInE_4_8_port <= '0';
   muxInD_4_0_port <= '0';
   muxInD_4_1_port <= '0';
   muxInD_4_2_port <= '0';
   muxInD_4_3_port <= '0';
   muxInD_4_4_port <= '0';
   muxInD_4_5_port <= '0';
   muxInD_4_6_port <= '0';
   muxInD_4_7_port <= '0';
   muxInD_4_8_port <= '0';
   muxInC_4_0_port <= '0';
   muxInC_4_1_port <= '0';
   muxInC_4_2_port <= '0';
   muxInC_4_3_port <= '0';
   muxInC_4_4_port <= '0';
   muxInC_4_5_port <= '0';
   muxInC_4_6_port <= '0';
   muxInC_4_7_port <= '0';
   muxInB_4_0_port <= '0';
   muxInB_4_1_port <= '0';
   muxInB_4_2_port <= '0';
   muxInB_4_3_port <= '0';
   muxInB_4_4_port <= '0';
   muxInB_4_5_port <= '0';
   muxInB_4_6_port <= '0';
   muxInB_4_7_port <= '0';
   muxInE_3_0_port <= '0';
   muxInE_3_1_port <= '0';
   muxInE_3_2_port <= '0';
   muxInE_3_3_port <= '0';
   muxInE_3_4_port <= '0';
   muxInE_3_5_port <= '0';
   muxInE_3_6_port <= '0';
   muxInD_3_0_port <= '0';
   muxInD_3_1_port <= '0';
   muxInD_3_2_port <= '0';
   muxInD_3_3_port <= '0';
   muxInD_3_4_port <= '0';
   muxInD_3_5_port <= '0';
   muxInD_3_6_port <= '0';
   muxInC_3_0_port <= '0';
   muxInC_3_1_port <= '0';
   muxInC_3_2_port <= '0';
   muxInC_3_3_port <= '0';
   muxInC_3_4_port <= '0';
   muxInC_3_5_port <= '0';
   muxInB_3_0_port <= '0';
   muxInB_3_1_port <= '0';
   muxInB_3_2_port <= '0';
   muxInB_3_3_port <= '0';
   muxInB_3_4_port <= '0';
   muxInB_3_5_port <= '0';
   muxInE_2_0_port <= '0';
   muxInE_2_1_port <= '0';
   muxInE_2_2_port <= '0';
   muxInE_2_3_port <= '0';
   muxInE_2_4_port <= '0';
   muxInD_2_0_port <= '0';
   muxInD_2_1_port <= '0';
   muxInD_2_2_port <= '0';
   muxInD_2_3_port <= '0';
   muxInD_2_4_port <= '0';
   muxInC_2_0_port <= '0';
   muxInC_2_1_port <= '0';
   muxInC_2_2_port <= '0';
   muxInC_2_3_port <= '0';
   muxInB_2_0_port <= '0';
   muxInB_2_1_port <= '0';
   muxInB_2_2_port <= '0';
   muxInB_2_3_port <= '0';
   muxInE_1_0_port <= '0';
   muxInE_1_1_port <= '0';
   muxInE_1_2_port <= '0';
   muxInD_1_0_port <= '0';
   muxInD_1_1_port <= '0';
   muxInD_1_2_port <= '0';
   muxInC_1_0_port <= '0';
   muxInC_1_1_port <= '0';
   muxInB_1_0_port <= '0';
   muxInB_1_1_port <= '0';
   muxInE_0_0_port <= '0';
   muxInD_0_0_port <= '0';
   U248 : BUF_X1 port map( A => A(12), Z => n25);
   U249 : BUF_X1 port map( A => A(8), Z => n18);
   U250 : BUF_X1 port map( A => A(11), Z => n22);
   U251 : BUF_X1 port map( A => A(14), Z => n27);
   U252 : BUF_X1 port map( A => A(10), Z => n21);
   U253 : BUF_X2 port map( A => A(13), Z => n26);
   U254 : BUF_X2 port map( A => A(9), Z => n19);
   U255 : BUF_X2 port map( A => A(3), Z => n11);
   U256 : BUF_X2 port map( A => A(7), Z => n17);
   U257 : BUF_X2 port map( A => A(1), Z => n10);
   U258 : BUF_X2 port map( A => A(0), Z => n2);
   U259 : BUF_X2 port map( A => A(5), Z => n14);
   U260 : BUF_X1 port map( A => A(6), Z => n15);
   U261 : BUF_X1 port map( A => A(0), Z => n3);
   U262 : BUF_X1 port map( A => A(4), Z => n13);
   U263 : BUF_X1 port map( A => A(15), Z => n28);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity adder_sub_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end adder_sub_N32;

architecture SYN_struct of adder_sub_N32 is

   component cla_adder_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component generic_xor_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, B_in_27_port,
      B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, B_in_22_port, 
      B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, B_in_17_port, 
      B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, B_in_12_port, 
      B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, B_in_7_port, 
      B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, B_in_2_port, 
      B_in_1_port, B_in_0_port : std_logic;

begin
   
   xor_g : generic_xor_N32 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => Ci, Y(31) => B_in_31_port, Y(30) => 
                           B_in_30_port, Y(29) => B_in_29_port, Y(28) => 
                           B_in_28_port, Y(27) => B_in_27_port, Y(26) => 
                           B_in_26_port, Y(25) => B_in_25_port, Y(24) => 
                           B_in_24_port, Y(23) => B_in_23_port, Y(22) => 
                           B_in_22_port, Y(21) => B_in_21_port, Y(20) => 
                           B_in_20_port, Y(19) => B_in_19_port, Y(18) => 
                           B_in_18_port, Y(17) => B_in_17_port, Y(16) => 
                           B_in_16_port, Y(15) => B_in_15_port, Y(14) => 
                           B_in_14_port, Y(13) => B_in_13_port, Y(12) => 
                           B_in_12_port, Y(11) => B_in_11_port, Y(10) => 
                           B_in_10_port, Y(9) => B_in_9_port, Y(8) => 
                           B_in_8_port, Y(7) => B_in_7_port, Y(6) => 
                           B_in_6_port, Y(5) => B_in_5_port, Y(4) => 
                           B_in_4_port, Y(3) => B_in_3_port, Y(2) => 
                           B_in_2_port, Y(1) => B_in_1_port, Y(0) => 
                           B_in_0_port);
   add : cla_adder_N32_0 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci => Ci, Cout => Cout, Sum(31) => 
                           Sum(31), Sum(30) => Sum(30), Sum(29) => Sum(29), 
                           Sum(28) => Sum(28), Sum(27) => Sum(27), Sum(26) => 
                           Sum(26), Sum(25) => Sum(25), Sum(24) => Sum(24), 
                           Sum(23) => Sum(23), Sum(22) => Sum(22), Sum(21) => 
                           Sum(21), Sum(20) => Sum(20), Sum(19) => Sum(19), 
                           Sum(18) => Sum(18), Sum(17) => Sum(17), Sum(16) => 
                           Sum(16), Sum(15) => Sum(15), Sum(14) => Sum(14), 
                           Sum(13) => Sum(13), Sum(12) => Sum(12), Sum(11) => 
                           Sum(11), Sum(10) => Sum(10), Sum(9) => Sum(9), 
                           Sum(8) => Sum(8), Sum(7) => Sum(7), Sum(6) => Sum(6)
                           , Sum(5) => Sum(5), Sum(4) => Sum(4), Sum(3) => 
                           Sum(3), Sum(2) => Sum(2), Sum(1) => Sum(1), Sum(0) 
                           => Sum(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_fwd_1 is

   port( OP, alu_out, alu_wb_in, lmd_out : in std_logic_vector (31 downto 0);  
         OPF : out std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (2 downto 0));

end mux_fwd_1;

architecture SYN_behav of mux_fwd_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n5, Z => n160);
   U2 : BUF_X1 port map( A => n5, Z => n159);
   U3 : BUF_X1 port map( A => n7, Z => n154);
   U4 : BUF_X1 port map( A => n7, Z => n153);
   U5 : BUF_X1 port map( A => n6, Z => n157);
   U6 : BUF_X1 port map( A => n6, Z => n156);
   U7 : BUF_X1 port map( A => n5, Z => n161);
   U8 : BUF_X1 port map( A => n7, Z => n155);
   U9 : BUF_X1 port map( A => n6, Z => n158);
   U10 : NOR3_X1 port map( A1 => sel(1), A2 => n164, A3 => n70, ZN => n5);
   U11 : INV_X1 port map( A => sel(0), ZN => n70);
   U12 : NOR3_X1 port map( A1 => sel(1), A2 => n164, A3 => sel(0), ZN => n6);
   U13 : BUF_X1 port map( A => sel(2), Z => n164);
   U14 : NOR2_X1 port map( A1 => n71, A2 => n164, ZN => n7);
   U15 : INV_X1 port map( A => sel(1), ZN => n71);
   U16 : BUF_X1 port map( A => sel(2), Z => n163);
   U17 : BUF_X1 port map( A => sel(2), Z => n162);
   U18 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => OPF(7));
   U19 : AOI22_X1 port map( A1 => alu_wb_in(7), A2 => n155, B1 => alu_out(7), 
                           B2 => n162, ZN => n10);
   U20 : AOI22_X1 port map( A1 => lmd_out(7), A2 => n161, B1 => OP(7), B2 => 
                           n158, ZN => n11);
   U21 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => OPF(0));
   U22 : AOI22_X1 port map( A1 => alu_wb_in(0), A2 => n153, B1 => alu_out(0), 
                           B2 => n164, ZN => n68);
   U23 : AOI22_X1 port map( A1 => lmd_out(0), A2 => n159, B1 => OP(0), B2 => 
                           n156, ZN => n69);
   U24 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => OPF(1));
   U25 : AOI22_X1 port map( A1 => alu_wb_in(1), A2 => n153, B1 => alu_out(1), 
                           B2 => n163, ZN => n46);
   U26 : AOI22_X1 port map( A1 => lmd_out(1), A2 => n159, B1 => OP(1), B2 => 
                           n156, ZN => n47);
   U27 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => OPF(2));
   U28 : AOI22_X1 port map( A1 => alu_wb_in(2), A2 => n154, B1 => alu_out(2), 
                           B2 => n162, ZN => n24);
   U29 : AOI22_X1 port map( A1 => lmd_out(2), A2 => n160, B1 => OP(2), B2 => 
                           n157, ZN => n25);
   U30 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => OPF(3));
   U31 : AOI22_X1 port map( A1 => alu_wb_in(3), A2 => n155, B1 => alu_out(3), 
                           B2 => n162, ZN => n18);
   U32 : AOI22_X1 port map( A1 => lmd_out(3), A2 => n161, B1 => OP(3), B2 => 
                           n158, ZN => n19);
   U33 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => OPF(4));
   U34 : AOI22_X1 port map( A1 => alu_wb_in(4), A2 => n155, B1 => alu_out(4), 
                           B2 => n162, ZN => n16);
   U35 : AOI22_X1 port map( A1 => lmd_out(4), A2 => n161, B1 => OP(4), B2 => 
                           n158, ZN => n17);
   U36 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => OPF(5));
   U37 : AOI22_X1 port map( A1 => alu_wb_in(5), A2 => n155, B1 => alu_out(5), 
                           B2 => n162, ZN => n14);
   U38 : AOI22_X1 port map( A1 => lmd_out(5), A2 => n161, B1 => OP(5), B2 => 
                           n158, ZN => n15);
   U39 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => OPF(6));
   U40 : AOI22_X1 port map( A1 => alu_wb_in(6), A2 => n155, B1 => alu_out(6), 
                           B2 => n162, ZN => n12);
   U41 : AOI22_X1 port map( A1 => lmd_out(6), A2 => n161, B1 => OP(6), B2 => 
                           n158, ZN => n13);
   U42 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => OPF(8));
   U43 : AOI22_X1 port map( A1 => alu_wb_in(8), A2 => n155, B1 => alu_out(8), 
                           B2 => n162, ZN => n8);
   U44 : AOI22_X1 port map( A1 => lmd_out(8), A2 => n161, B1 => OP(8), B2 => 
                           n158, ZN => n9);
   U45 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OPF(9));
   U46 : AOI22_X1 port map( A1 => alu_wb_in(9), A2 => n155, B1 => n164, B2 => 
                           alu_out(9), ZN => n3);
   U47 : AOI22_X1 port map( A1 => lmd_out(9), A2 => n161, B1 => OP(9), B2 => 
                           n158, ZN => n4);
   U48 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => OPF(10));
   U49 : AOI22_X1 port map( A1 => alu_wb_in(10), A2 => n153, B1 => alu_out(10),
                           B2 => n164, ZN => n66);
   U50 : AOI22_X1 port map( A1 => lmd_out(10), A2 => n159, B1 => OP(10), B2 => 
                           n156, ZN => n67);
   U51 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => OPF(11));
   U52 : AOI22_X1 port map( A1 => alu_wb_in(11), A2 => n153, B1 => alu_out(11),
                           B2 => n164, ZN => n64);
   U53 : AOI22_X1 port map( A1 => lmd_out(11), A2 => n159, B1 => OP(11), B2 => 
                           n156, ZN => n65);
   U54 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => OPF(12));
   U55 : AOI22_X1 port map( A1 => alu_wb_in(12), A2 => n153, B1 => alu_out(12),
                           B2 => n164, ZN => n62);
   U56 : AOI22_X1 port map( A1 => lmd_out(12), A2 => n159, B1 => OP(12), B2 => 
                           n156, ZN => n63);
   U57 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => OPF(13));
   U58 : AOI22_X1 port map( A1 => alu_wb_in(13), A2 => n153, B1 => alu_out(13),
                           B2 => n164, ZN => n60);
   U59 : AOI22_X1 port map( A1 => lmd_out(13), A2 => n159, B1 => OP(13), B2 => 
                           n156, ZN => n61);
   U60 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => OPF(14));
   U61 : AOI22_X1 port map( A1 => alu_wb_in(14), A2 => n153, B1 => alu_out(14),
                           B2 => n164, ZN => n58);
   U62 : AOI22_X1 port map( A1 => lmd_out(14), A2 => n159, B1 => OP(14), B2 => 
                           n156, ZN => n59);
   U63 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => OPF(15));
   U64 : AOI22_X1 port map( A1 => alu_wb_in(15), A2 => n153, B1 => alu_out(15),
                           B2 => n164, ZN => n56);
   U65 : AOI22_X1 port map( A1 => lmd_out(15), A2 => n159, B1 => OP(15), B2 => 
                           n156, ZN => n57);
   U66 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => OPF(31));
   U67 : AOI22_X1 port map( A1 => alu_wb_in(31), A2 => n155, B1 => alu_out(31),
                           B2 => n162, ZN => n20);
   U68 : AOI22_X1 port map( A1 => lmd_out(31), A2 => n161, B1 => OP(31), B2 => 
                           n158, ZN => n21);
   U69 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => OPF(16));
   U70 : AOI22_X1 port map( A1 => alu_wb_in(16), A2 => n153, B1 => alu_out(16),
                           B2 => n163, ZN => n54);
   U71 : AOI22_X1 port map( A1 => lmd_out(16), A2 => n159, B1 => OP(16), B2 => 
                           n156, ZN => n55);
   U72 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => OPF(17));
   U73 : AOI22_X1 port map( A1 => alu_wb_in(17), A2 => n153, B1 => alu_out(17),
                           B2 => n163, ZN => n52);
   U74 : AOI22_X1 port map( A1 => lmd_out(17), A2 => n159, B1 => OP(17), B2 => 
                           n156, ZN => n53);
   U75 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => OPF(18));
   U76 : AOI22_X1 port map( A1 => alu_wb_in(18), A2 => n153, B1 => alu_out(18),
                           B2 => n163, ZN => n50);
   U77 : AOI22_X1 port map( A1 => lmd_out(18), A2 => n159, B1 => OP(18), B2 => 
                           n156, ZN => n51);
   U78 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => OPF(19));
   U79 : AOI22_X1 port map( A1 => alu_wb_in(19), A2 => n153, B1 => alu_out(19),
                           B2 => n163, ZN => n48);
   U80 : AOI22_X1 port map( A1 => lmd_out(19), A2 => n159, B1 => OP(19), B2 => 
                           n156, ZN => n49);
   U81 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => OPF(20));
   U82 : AOI22_X1 port map( A1 => alu_wb_in(20), A2 => n154, B1 => alu_out(20),
                           B2 => n163, ZN => n44);
   U83 : AOI22_X1 port map( A1 => lmd_out(20), A2 => n160, B1 => OP(20), B2 => 
                           n157, ZN => n45);
   U84 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => OPF(21));
   U85 : AOI22_X1 port map( A1 => alu_wb_in(21), A2 => n154, B1 => alu_out(21),
                           B2 => n163, ZN => n42);
   U86 : AOI22_X1 port map( A1 => lmd_out(21), A2 => n160, B1 => OP(21), B2 => 
                           n157, ZN => n43);
   U87 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => OPF(22));
   U88 : AOI22_X1 port map( A1 => alu_wb_in(22), A2 => n154, B1 => alu_out(22),
                           B2 => n163, ZN => n40);
   U89 : AOI22_X1 port map( A1 => lmd_out(22), A2 => n160, B1 => OP(22), B2 => 
                           n157, ZN => n41);
   U90 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => OPF(23));
   U91 : AOI22_X1 port map( A1 => alu_wb_in(23), A2 => n154, B1 => alu_out(23),
                           B2 => n163, ZN => n38);
   U92 : AOI22_X1 port map( A1 => lmd_out(23), A2 => n160, B1 => OP(23), B2 => 
                           n157, ZN => n39);
   U93 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => OPF(24));
   U94 : AOI22_X1 port map( A1 => alu_wb_in(24), A2 => n154, B1 => alu_out(24),
                           B2 => n163, ZN => n36);
   U95 : AOI22_X1 port map( A1 => lmd_out(24), A2 => n160, B1 => OP(24), B2 => 
                           n157, ZN => n37);
   U96 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => OPF(25));
   U97 : AOI22_X1 port map( A1 => alu_wb_in(25), A2 => n154, B1 => alu_out(25),
                           B2 => n163, ZN => n34);
   U98 : AOI22_X1 port map( A1 => lmd_out(25), A2 => n160, B1 => OP(25), B2 => 
                           n157, ZN => n35);
   U99 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => OPF(26));
   U100 : AOI22_X1 port map( A1 => alu_wb_in(26), A2 => n154, B1 => alu_out(26)
                           , B2 => n162, ZN => n32);
   U101 : AOI22_X1 port map( A1 => lmd_out(26), A2 => n160, B1 => OP(26), B2 =>
                           n157, ZN => n33);
   U102 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => OPF(27));
   U103 : AOI22_X1 port map( A1 => alu_wb_in(27), A2 => n154, B1 => alu_out(27)
                           , B2 => n162, ZN => n30);
   U104 : AOI22_X1 port map( A1 => lmd_out(27), A2 => n160, B1 => OP(27), B2 =>
                           n157, ZN => n31);
   U105 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => OPF(28));
   U106 : AOI22_X1 port map( A1 => alu_wb_in(28), A2 => n154, B1 => alu_out(28)
                           , B2 => n162, ZN => n28);
   U107 : AOI22_X1 port map( A1 => lmd_out(28), A2 => n160, B1 => OP(28), B2 =>
                           n157, ZN => n29);
   U108 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => OPF(29));
   U109 : AOI22_X1 port map( A1 => alu_wb_in(29), A2 => n154, B1 => alu_out(29)
                           , B2 => n162, ZN => n26);
   U110 : AOI22_X1 port map( A1 => lmd_out(29), A2 => n160, B1 => OP(29), B2 =>
                           n157, ZN => n27);
   U111 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => OPF(30));
   U112 : AOI22_X1 port map( A1 => alu_wb_in(30), A2 => n154, B1 => alu_out(30)
                           , B2 => n163, ZN => n22);
   U113 : AOI22_X1 port map( A1 => lmd_out(30), A2 => n160, B1 => OP(30), B2 =>
                           n157, ZN => n23);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_fwd_0 is

   port( OP, alu_out, alu_wb_in, lmd_out : in std_logic_vector (31 downto 0);  
         OPF : out std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (2 downto 0));

end mux_fwd_0;

architecture SYN_behav of mux_fwd_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n5, Z => n89);
   U2 : BUF_X1 port map( A => n5, Z => n90);
   U3 : BUF_X1 port map( A => n7, Z => n83);
   U4 : BUF_X1 port map( A => n7, Z => n84);
   U5 : BUF_X1 port map( A => n6, Z => n86);
   U6 : BUF_X1 port map( A => n6, Z => n87);
   U7 : BUF_X1 port map( A => n5, Z => n91);
   U8 : BUF_X1 port map( A => n7, Z => n85);
   U9 : BUF_X1 port map( A => n6, Z => n88);
   U10 : NOR3_X1 port map( A1 => sel(1), A2 => n94, A3 => n70, ZN => n5);
   U11 : INV_X1 port map( A => sel(0), ZN => n70);
   U12 : NOR3_X1 port map( A1 => sel(1), A2 => n94, A3 => sel(0), ZN => n6);
   U13 : BUF_X1 port map( A => sel(2), Z => n94);
   U14 : NOR2_X1 port map( A1 => n71, A2 => n94, ZN => n7);
   U15 : INV_X1 port map( A => sel(1), ZN => n71);
   U16 : BUF_X1 port map( A => sel(2), Z => n93);
   U17 : BUF_X1 port map( A => sel(2), Z => n92);
   U18 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => OPF(31));
   U19 : AOI22_X1 port map( A1 => alu_wb_in(31), A2 => n85, B1 => alu_out(31), 
                           B2 => n92, ZN => n20);
   U20 : AOI22_X1 port map( A1 => lmd_out(31), A2 => n91, B1 => OP(31), B2 => 
                           n88, ZN => n21);
   U21 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => OPF(7));
   U22 : AOI22_X1 port map( A1 => alu_wb_in(7), A2 => n85, B1 => alu_out(7), B2
                           => n92, ZN => n10);
   U23 : AOI22_X1 port map( A1 => lmd_out(7), A2 => n91, B1 => OP(7), B2 => n88
                           , ZN => n11);
   U24 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => OPF(0));
   U25 : AOI22_X1 port map( A1 => alu_wb_in(0), A2 => n83, B1 => alu_out(0), B2
                           => n94, ZN => n68);
   U26 : AOI22_X1 port map( A1 => lmd_out(0), A2 => n89, B1 => OP(0), B2 => n86
                           , ZN => n69);
   U27 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => OPF(1));
   U28 : AOI22_X1 port map( A1 => alu_wb_in(1), A2 => n83, B1 => alu_out(1), B2
                           => n93, ZN => n46);
   U29 : AOI22_X1 port map( A1 => lmd_out(1), A2 => n89, B1 => OP(1), B2 => n86
                           , ZN => n47);
   U30 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => OPF(2));
   U31 : AOI22_X1 port map( A1 => alu_wb_in(2), A2 => n84, B1 => alu_out(2), B2
                           => n92, ZN => n24);
   U32 : AOI22_X1 port map( A1 => lmd_out(2), A2 => n90, B1 => OP(2), B2 => n87
                           , ZN => n25);
   U33 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => OPF(3));
   U34 : AOI22_X1 port map( A1 => alu_wb_in(3), A2 => n85, B1 => alu_out(3), B2
                           => n92, ZN => n18);
   U35 : AOI22_X1 port map( A1 => lmd_out(3), A2 => n91, B1 => OP(3), B2 => n88
                           , ZN => n19);
   U36 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => OPF(4));
   U37 : AOI22_X1 port map( A1 => alu_wb_in(4), A2 => n85, B1 => alu_out(4), B2
                           => n92, ZN => n16);
   U38 : AOI22_X1 port map( A1 => lmd_out(4), A2 => n91, B1 => OP(4), B2 => n88
                           , ZN => n17);
   U39 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => OPF(5));
   U40 : AOI22_X1 port map( A1 => alu_wb_in(5), A2 => n85, B1 => alu_out(5), B2
                           => n92, ZN => n14);
   U41 : AOI22_X1 port map( A1 => lmd_out(5), A2 => n91, B1 => OP(5), B2 => n88
                           , ZN => n15);
   U42 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => OPF(6));
   U43 : AOI22_X1 port map( A1 => alu_wb_in(6), A2 => n85, B1 => alu_out(6), B2
                           => n92, ZN => n12);
   U44 : AOI22_X1 port map( A1 => lmd_out(6), A2 => n91, B1 => OP(6), B2 => n88
                           , ZN => n13);
   U45 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => OPF(8));
   U46 : AOI22_X1 port map( A1 => alu_wb_in(8), A2 => n85, B1 => alu_out(8), B2
                           => n92, ZN => n8);
   U47 : AOI22_X1 port map( A1 => lmd_out(8), A2 => n91, B1 => OP(8), B2 => n88
                           , ZN => n9);
   U48 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OPF(9));
   U49 : AOI22_X1 port map( A1 => alu_wb_in(9), A2 => n85, B1 => n94, B2 => 
                           alu_out(9), ZN => n3);
   U50 : AOI22_X1 port map( A1 => lmd_out(9), A2 => n91, B1 => OP(9), B2 => n88
                           , ZN => n4);
   U51 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => OPF(10));
   U52 : AOI22_X1 port map( A1 => alu_wb_in(10), A2 => n83, B1 => alu_out(10), 
                           B2 => n94, ZN => n66);
   U53 : AOI22_X1 port map( A1 => lmd_out(10), A2 => n89, B1 => OP(10), B2 => 
                           n86, ZN => n67);
   U54 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => OPF(11));
   U55 : AOI22_X1 port map( A1 => alu_wb_in(11), A2 => n83, B1 => alu_out(11), 
                           B2 => n94, ZN => n64);
   U56 : AOI22_X1 port map( A1 => lmd_out(11), A2 => n89, B1 => OP(11), B2 => 
                           n86, ZN => n65);
   U57 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => OPF(12));
   U58 : AOI22_X1 port map( A1 => alu_wb_in(12), A2 => n83, B1 => alu_out(12), 
                           B2 => n94, ZN => n62);
   U59 : AOI22_X1 port map( A1 => lmd_out(12), A2 => n89, B1 => OP(12), B2 => 
                           n86, ZN => n63);
   U60 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => OPF(13));
   U61 : AOI22_X1 port map( A1 => alu_wb_in(13), A2 => n83, B1 => alu_out(13), 
                           B2 => n94, ZN => n60);
   U62 : AOI22_X1 port map( A1 => lmd_out(13), A2 => n89, B1 => OP(13), B2 => 
                           n86, ZN => n61);
   U63 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => OPF(14));
   U64 : AOI22_X1 port map( A1 => alu_wb_in(14), A2 => n83, B1 => alu_out(14), 
                           B2 => n94, ZN => n58);
   U65 : AOI22_X1 port map( A1 => lmd_out(14), A2 => n89, B1 => OP(14), B2 => 
                           n86, ZN => n59);
   U66 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => OPF(15));
   U67 : AOI22_X1 port map( A1 => alu_wb_in(15), A2 => n83, B1 => alu_out(15), 
                           B2 => n94, ZN => n56);
   U68 : AOI22_X1 port map( A1 => lmd_out(15), A2 => n89, B1 => OP(15), B2 => 
                           n86, ZN => n57);
   U69 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => OPF(16));
   U70 : AOI22_X1 port map( A1 => alu_wb_in(16), A2 => n83, B1 => alu_out(16), 
                           B2 => n93, ZN => n54);
   U71 : AOI22_X1 port map( A1 => lmd_out(16), A2 => n89, B1 => OP(16), B2 => 
                           n86, ZN => n55);
   U72 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => OPF(17));
   U73 : AOI22_X1 port map( A1 => alu_wb_in(17), A2 => n83, B1 => alu_out(17), 
                           B2 => n93, ZN => n52);
   U74 : AOI22_X1 port map( A1 => lmd_out(17), A2 => n89, B1 => OP(17), B2 => 
                           n86, ZN => n53);
   U75 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => OPF(18));
   U76 : AOI22_X1 port map( A1 => alu_wb_in(18), A2 => n83, B1 => alu_out(18), 
                           B2 => n93, ZN => n50);
   U77 : AOI22_X1 port map( A1 => lmd_out(18), A2 => n89, B1 => OP(18), B2 => 
                           n86, ZN => n51);
   U78 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => OPF(19));
   U79 : AOI22_X1 port map( A1 => alu_wb_in(19), A2 => n83, B1 => alu_out(19), 
                           B2 => n93, ZN => n48);
   U80 : AOI22_X1 port map( A1 => lmd_out(19), A2 => n89, B1 => OP(19), B2 => 
                           n86, ZN => n49);
   U81 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => OPF(20));
   U82 : AOI22_X1 port map( A1 => alu_wb_in(20), A2 => n84, B1 => alu_out(20), 
                           B2 => n93, ZN => n44);
   U83 : AOI22_X1 port map( A1 => lmd_out(20), A2 => n90, B1 => OP(20), B2 => 
                           n87, ZN => n45);
   U84 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => OPF(21));
   U85 : AOI22_X1 port map( A1 => alu_wb_in(21), A2 => n84, B1 => alu_out(21), 
                           B2 => n93, ZN => n42);
   U86 : AOI22_X1 port map( A1 => lmd_out(21), A2 => n90, B1 => OP(21), B2 => 
                           n87, ZN => n43);
   U87 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => OPF(22));
   U88 : AOI22_X1 port map( A1 => alu_wb_in(22), A2 => n84, B1 => alu_out(22), 
                           B2 => n93, ZN => n40);
   U89 : AOI22_X1 port map( A1 => lmd_out(22), A2 => n90, B1 => OP(22), B2 => 
                           n87, ZN => n41);
   U90 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => OPF(23));
   U91 : AOI22_X1 port map( A1 => alu_wb_in(23), A2 => n84, B1 => alu_out(23), 
                           B2 => n93, ZN => n38);
   U92 : AOI22_X1 port map( A1 => lmd_out(23), A2 => n90, B1 => OP(23), B2 => 
                           n87, ZN => n39);
   U93 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => OPF(24));
   U94 : AOI22_X1 port map( A1 => alu_wb_in(24), A2 => n84, B1 => alu_out(24), 
                           B2 => n93, ZN => n36);
   U95 : AOI22_X1 port map( A1 => lmd_out(24), A2 => n90, B1 => OP(24), B2 => 
                           n87, ZN => n37);
   U96 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => OPF(25));
   U97 : AOI22_X1 port map( A1 => alu_wb_in(25), A2 => n84, B1 => alu_out(25), 
                           B2 => n93, ZN => n34);
   U98 : AOI22_X1 port map( A1 => lmd_out(25), A2 => n90, B1 => OP(25), B2 => 
                           n87, ZN => n35);
   U99 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => OPF(26));
   U100 : AOI22_X1 port map( A1 => alu_wb_in(26), A2 => n84, B1 => alu_out(26),
                           B2 => n92, ZN => n32);
   U101 : AOI22_X1 port map( A1 => lmd_out(26), A2 => n90, B1 => OP(26), B2 => 
                           n87, ZN => n33);
   U102 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => OPF(27));
   U103 : AOI22_X1 port map( A1 => alu_wb_in(27), A2 => n84, B1 => alu_out(27),
                           B2 => n92, ZN => n30);
   U104 : AOI22_X1 port map( A1 => lmd_out(27), A2 => n90, B1 => OP(27), B2 => 
                           n87, ZN => n31);
   U105 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => OPF(28));
   U106 : AOI22_X1 port map( A1 => alu_wb_in(28), A2 => n84, B1 => alu_out(28),
                           B2 => n92, ZN => n28);
   U107 : AOI22_X1 port map( A1 => lmd_out(28), A2 => n90, B1 => OP(28), B2 => 
                           n87, ZN => n29);
   U108 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => OPF(29));
   U109 : AOI22_X1 port map( A1 => alu_wb_in(29), A2 => n84, B1 => alu_out(29),
                           B2 => n92, ZN => n26);
   U110 : AOI22_X1 port map( A1 => lmd_out(29), A2 => n90, B1 => OP(29), B2 => 
                           n87, ZN => n27);
   U111 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => OPF(30));
   U112 : AOI22_X1 port map( A1 => alu_wb_in(30), A2 => n84, B1 => alu_out(30),
                           B2 => n93, ZN => n22);
   U113 : AOI22_X1 port map( A1 => lmd_out(30), A2 => n90, B1 => OP(30), B2 => 
                           n87, ZN => n23);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity counter is

   port( clk, rst : in std_logic;  tc : out std_logic);

end counter;

architecture SYN_rtl of counter is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component counter_DW01_dec_0
      port( A : in std_logic_vector (30 downto 0);  SUM : out std_logic_vector 
            (30 downto 0));
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal i_30_port, i_29_port, i_28_port, i_27_port, i_26_port, i_25_port, 
      i_24_port, i_23_port, i_22_port, i_21_port, i_20_port, i_19_port, 
      i_18_port, i_17_port, i_16_port, i_15_port, i_14_port, i_13_port, 
      i_12_port, i_11_port, i_10_port, i_9_port, i_8_port, i_7_port, i_6_port, 
      i_5_port, i_4_port, i_3_port, i_2_port, i_1_port, i_0_port, N4, N5, N6, 
      N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, 
      N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N125, N127, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, net227481, net227482, net227483, 
      net227484, net227485, net227486, net227487, net227488, net227489, 
      net227490, net227491, net227492, net227493, net227494, net227495, 
      net227496, net227497, net227498, net227499, net227500, net227501, 
      net227502, net227503, net227504, net227505, net227506, net227507, 
      net227508, net227509, net227510, net227511, n32_port, n33_port, n34, n35,
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n119, n120, n121, n122, n123 : std_logic;

begin
   
   i_reg_0_inst : DFFR_X1 port map( D => n118, CK => clk, RN => n121, Q => 
                           i_0_port, QN => net227511);
   i_reg_30_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n122, Q => 
                           i_30_port, QN => net227510);
   i_reg_28_inst : DFFR_X1 port map( D => n116, CK => clk, RN => n122, Q => 
                           i_28_port, QN => net227509);
   i_reg_26_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n122, Q => 
                           i_26_port, QN => net227508);
   i_reg_24_inst : DFFR_X1 port map( D => n114, CK => clk, RN => n122, Q => 
                           i_24_port, QN => net227507);
   i_reg_22_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n122, Q => 
                           i_22_port, QN => net227506);
   i_reg_20_inst : DFFR_X1 port map( D => n112, CK => clk, RN => n122, Q => 
                           i_20_port, QN => net227505);
   i_reg_18_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n121, Q => 
                           i_18_port, QN => net227504);
   i_reg_16_inst : DFFR_X1 port map( D => n110, CK => clk, RN => n121, Q => 
                           i_16_port, QN => net227503);
   i_reg_14_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n121, Q => 
                           i_14_port, QN => net227502);
   i_reg_12_inst : DFFR_X1 port map( D => n108, CK => clk, RN => n121, Q => 
                           i_12_port, QN => net227501);
   i_reg_10_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n121, Q => 
                           i_10_port, QN => net227500);
   i_reg_8_inst : DFFR_X1 port map( D => n106, CK => clk, RN => n122, Q => 
                           i_8_port, QN => net227499);
   i_reg_6_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n123, Q => 
                           i_6_port, QN => net227498);
   i_reg_4_inst : DFFR_X1 port map( D => n104, CK => clk, RN => n123, Q => 
                           i_4_port, QN => net227497);
   i_reg_2_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n122, Q => 
                           i_2_port, QN => net227496);
   i_reg_1_inst : DFFS_X1 port map( D => n102, CK => clk, SN => n123, Q => 
                           i_1_port, QN => net227495);
   i_reg_3_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n123, Q => 
                           i_3_port, QN => net227494);
   i_reg_5_inst : DFFR_X1 port map( D => n100, CK => clk, RN => n123, Q => 
                           i_5_port, QN => net227493);
   i_reg_7_inst : DFFR_X1 port map( D => n99, CK => clk, RN => n123, Q => 
                           i_7_port, QN => net227492);
   i_reg_9_inst : DFFR_X1 port map( D => n98, CK => clk, RN => n123, Q => 
                           i_9_port, QN => net227491);
   i_reg_11_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n122, Q => 
                           i_11_port, QN => net227490);
   i_reg_13_inst : DFFR_X1 port map( D => n96, CK => clk, RN => n122, Q => 
                           i_13_port, QN => net227489);
   i_reg_15_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n122, Q => 
                           i_15_port, QN => net227488);
   i_reg_17_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n121, Q => 
                           i_17_port, QN => net227487);
   i_reg_19_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n122, Q => 
                           i_19_port, QN => net227486);
   i_reg_21_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n121, Q => 
                           i_21_port, QN => net227485);
   i_reg_23_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n121, Q => 
                           i_23_port, QN => net227484);
   i_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n121, Q => 
                           i_25_port, QN => net227483);
   i_reg_27_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n121, Q => 
                           i_27_port, QN => net227482);
   i_reg_29_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n121, Q => 
                           i_29_port, QN => net227481);
   tc_reg : DFFS_X1 port map( D => N125, CK => clk, SN => n123, Q => tc, QN => 
                           n87);
   sub_19 : counter_DW01_dec_0 port map( A(30) => i_30_port, A(29) => i_29_port
                           , A(28) => i_28_port, A(27) => i_27_port, A(26) => 
                           i_26_port, A(25) => i_25_port, A(24) => i_24_port, 
                           A(23) => i_23_port, A(22) => i_22_port, A(21) => 
                           i_21_port, A(20) => i_20_port, A(19) => i_19_port, 
                           A(18) => i_18_port, A(17) => i_17_port, A(16) => 
                           i_16_port, A(15) => i_15_port, A(14) => i_14_port, 
                           A(13) => i_13_port, A(12) => i_12_port, A(11) => 
                           i_11_port, A(10) => i_10_port, A(9) => i_9_port, 
                           A(8) => i_8_port, A(7) => i_7_port, A(6) => i_6_port
                           , A(5) => i_5_port, A(4) => i_4_port, A(3) => 
                           i_3_port, A(2) => i_2_port, A(1) => i_1_port, A(0) 
                           => i_0_port, SUM(30) => N33, SUM(29) => N32, SUM(28)
                           => N31, SUM(27) => N30, SUM(26) => N29, SUM(25) => 
                           N28, SUM(24) => N27, SUM(23) => N26, SUM(22) => N25,
                           SUM(21) => N24, SUM(20) => N23, SUM(19) => N22, 
                           SUM(18) => N21, SUM(17) => N20, SUM(16) => N19, 
                           SUM(15) => N18, SUM(14) => N17, SUM(13) => N16, 
                           SUM(12) => N15, SUM(11) => N14, SUM(10) => N13, 
                           SUM(9) => N12, SUM(8) => N11, SUM(7) => N10, SUM(6) 
                           => N9, SUM(5) => N8, SUM(4) => N7, SUM(3) => N6, 
                           SUM(2) => N5, SUM(1) => N127, SUM(0) => N4);
   U3 : OR3_X1 port map( A1 => n77, A2 => n78, A3 => n76, ZN => n84);
   U4 : NOR2_X1 port map( A1 => n120, A2 => n39, ZN => n93);
   U5 : NOR2_X1 port map( A1 => n120, A2 => n37, ZN => n95);
   U6 : NOR2_X1 port map( A1 => n119, A2 => n47, ZN => n116);
   U7 : INV_X1 port map( A => N31, ZN => n47);
   U8 : NOR2_X1 port map( A1 => n119, A2 => n41, ZN => n91);
   U9 : INV_X1 port map( A => N26, ZN => n41);
   U10 : NOR2_X1 port map( A1 => n119, A2 => n52, ZN => n111);
   U11 : NOR2_X1 port map( A1 => n119, A2 => n51, ZN => n112);
   U12 : NOR2_X1 port map( A1 => n119, A2 => n50, ZN => n113);
   U13 : INV_X1 port map( A => N25, ZN => n50);
   U14 : NOR2_X1 port map( A1 => n119, A2 => n48, ZN => n115);
   U15 : INV_X1 port map( A => N29, ZN => n48);
   U16 : NOR2_X1 port map( A1 => n86, A2 => n57, ZN => n106);
   U17 : NOR2_X1 port map( A1 => n86, A2 => n56, ZN => n107);
   U18 : INV_X1 port map( A => N13, ZN => n56);
   U19 : NOR4_X1 port map( A1 => N15, A2 => N14, A3 => N13, A4 => N127, ZN => 
                           n79);
   U20 : NOR4_X1 port map( A1 => N9, A2 => N8, A3 => N7, A4 => N6, ZN => n83);
   U21 : NOR4_X1 port map( A1 => N31, A2 => N30, A3 => N29, A4 => N28, ZN => 
                           n81);
   U22 : NOR4_X1 port map( A1 => N27, A2 => N26, A3 => N25, A4 => N24, ZN => 
                           n80);
   U23 : OR2_X1 port map( A1 => N5, A2 => N4, ZN => n85);
   U24 : INV_X1 port map( A => N21, ZN => n52);
   U25 : NOR2_X1 port map( A1 => n120, A2 => n40, ZN => n92);
   U26 : INV_X1 port map( A => N24, ZN => n40);
   U27 : NOR2_X1 port map( A1 => n120, A2 => n38, ZN => n94);
   U28 : NOR2_X1 port map( A1 => n120, A2 => n36, ZN => n96);
   U29 : NOR2_X1 port map( A1 => n120, A2 => n35, ZN => n97);
   U30 : INV_X1 port map( A => N14, ZN => n35);
   U31 : NOR2_X1 port map( A1 => n120, A2 => n34, ZN => n98);
   U32 : NOR2_X1 port map( A1 => n120, A2 => n33_port, ZN => n99);
   U33 : NOR2_X1 port map( A1 => n119, A2 => n44, ZN => n88);
   U34 : INV_X1 port map( A => N32, ZN => n44);
   U35 : NOR2_X1 port map( A1 => n119, A2 => n43, ZN => n89);
   U36 : INV_X1 port map( A => N30, ZN => n43);
   U37 : NOR2_X1 port map( A1 => n119, A2 => n46, ZN => n117);
   U38 : NOR2_X1 port map( A1 => n119, A2 => n42, ZN => n90);
   U39 : INV_X1 port map( A => N28, ZN => n42);
   U40 : NOR2_X1 port map( A1 => n119, A2 => n49, ZN => n114);
   U41 : INV_X1 port map( A => N27, ZN => n49);
   U42 : NOR2_X1 port map( A1 => n86, A2 => n55, ZN => n108);
   U43 : INV_X1 port map( A => N15, ZN => n55);
   U44 : NOR2_X1 port map( A1 => n86, A2 => n54, ZN => n109);
   U45 : NOR2_X1 port map( A1 => n86, A2 => n53, ZN => n110);
   U46 : INV_X1 port map( A => N18, ZN => n37);
   U47 : INV_X1 port map( A => N22, ZN => n39);
   U48 : INV_X1 port map( A => N11, ZN => n57);
   U49 : INV_X1 port map( A => N23, ZN => n51);
   U50 : BUF_X1 port map( A => n32_port, Z => n119);
   U51 : BUF_X1 port map( A => n32_port, Z => n86);
   U52 : BUF_X1 port map( A => n32_port, Z => n120);
   U53 : NOR2_X1 port map( A1 => n86, A2 => n61, ZN => n102);
   U54 : INV_X1 port map( A => N127, ZN => n61);
   U55 : NOR2_X1 port map( A1 => n119, A2 => n45, ZN => n118);
   U56 : INV_X1 port map( A => N4, ZN => n45);
   U57 : NOR2_X1 port map( A1 => n86, A2 => n63, ZN => n100);
   U58 : INV_X1 port map( A => N8, ZN => n63);
   U59 : NOR2_X1 port map( A1 => n86, A2 => n62, ZN => n101);
   U60 : INV_X1 port map( A => N6, ZN => n62);
   U61 : NOR2_X1 port map( A1 => n86, A2 => n60, ZN => n103);
   U62 : INV_X1 port map( A => N5, ZN => n60);
   U63 : NOR2_X1 port map( A1 => n86, A2 => n59, ZN => n104);
   U64 : INV_X1 port map( A => N7, ZN => n59);
   U65 : NOR2_X1 port map( A1 => n86, A2 => n58, ZN => n105);
   U66 : INV_X1 port map( A => N9, ZN => n58);
   U67 : BUF_X1 port map( A => rst, Z => n122);
   U68 : BUF_X1 port map( A => rst, Z => n121);
   U69 : BUF_X1 port map( A => rst, Z => n123);
   U70 : INV_X1 port map( A => N19, ZN => n53);
   U71 : INV_X1 port map( A => N20, ZN => n38);
   U72 : INV_X1 port map( A => N17, ZN => n54);
   U73 : INV_X1 port map( A => N10, ZN => n33_port);
   U74 : INV_X1 port map( A => N12, ZN => n34);
   U75 : INV_X1 port map( A => N16, ZN => n36);
   U76 : NOR4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           n69);
   U77 : NAND4_X1 port map( A1 => net227484, A2 => net227483, A3 => net227482, 
                           A4 => net227481, ZN => n70);
   U78 : NAND4_X1 port map( A1 => net227488, A2 => net227487, A3 => net227486, 
                           A4 => net227485, ZN => n71);
   U79 : NAND4_X1 port map( A1 => net227492, A2 => net227491, A3 => net227490, 
                           A4 => net227489, ZN => n72);
   U80 : NAND4_X1 port map( A1 => net227496, A2 => net227495, A3 => net227494, 
                           A4 => net227493, ZN => n73);
   U81 : NAND4_X1 port map( A1 => net227508, A2 => net227507, A3 => net227506, 
                           A4 => net227505, ZN => n74);
   U82 : AND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n69, ZN => 
                           n32_port);
   U83 : NOR4_X1 port map( A1 => i_12_port, A2 => i_14_port, A3 => i_16_port, 
                           A4 => i_18_port, ZN => n65);
   U84 : NOR4_X1 port map( A1 => i_4_port, A2 => i_6_port, A3 => i_8_port, A4 
                           => i_10_port, ZN => n66);
   U85 : NOR3_X1 port map( A1 => N33, A2 => N32, A3 => n85, ZN => n82);
   U86 : NOR2_X1 port map( A1 => n75, A2 => n84, ZN => n64);
   U87 : NAND4_X1 port map( A1 => n57, A2 => n34, A3 => n33_port, A4 => n79, ZN
                           => n76);
   U88 : NAND4_X1 port map( A1 => n38, A2 => n52, A3 => n39, A4 => n51, ZN => 
                           n77);
   U89 : NAND4_X1 port map( A1 => n36, A2 => n54, A3 => n37, A4 => n53, ZN => 
                           n78);
   U90 : NOR2_X1 port map( A1 => n64, A2 => n86, ZN => N125);
   U91 : NOR4_X1 port map( A1 => n74, A2 => i_0_port, A3 => i_28_port, A4 => 
                           i_30_port, ZN => n67);
   U92 : INV_X1 port map( A => N33, ZN => n46);
   U93 : NAND4_X1 port map( A1 => n80, A2 => n81, A3 => n82, A4 => n83, ZN => 
                           n75);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N2_0 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (1 downto 0);  
         d_out : out std_logic_vector (1 downto 0));

end reg_N2_0;

architecture SYN_behav of reg_N2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, n1, n3_port : std_logic;

begin
   
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n1);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n3_port);
   U3 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U4 : AND2_X1 port map( A1 => rst, A2 => d_in(1), ZN => N3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity mux_pc is

   port( A, B, C, D, E, F : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux_pc;

architecture SYN_behav of mux_pc is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n23, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   Y_tri_12_inst : TBUF_X1 port map( A => n126, EN => n169, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n125, EN => n169, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n124, EN => n169, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n123, EN => n169, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n122, EN => n169, Z => Y(16));
   Y_tri_18_inst : TBUF_X1 port map( A => n120, EN => n169, Z => Y(18));
   Y_tri_21_inst : TBUF_X1 port map( A => n117, EN => n169, Z => Y(21));
   Y_tri_23_inst : TBUF_X1 port map( A => n115, EN => n169, Z => Y(23));
   Y_tri_3_inst : TBUF_X1 port map( A => n136, EN => n167, Z => Y(3));
   Y_tri_5_inst : TBUF_X1 port map( A => n134, EN => n167, Z => Y(5));
   Y_tri_7_inst : TBUF_X1 port map( A => n132, EN => n167, Z => Y(7));
   Y_tri_9_inst : TBUF_X1 port map( A => n129, EN => n167, Z => Y(9));
   Y_tri_25_inst : TBUF_X1 port map( A => n113, EN => n167, Z => Y(25));
   Y_tri_27_inst : TBUF_X1 port map( A => n111, EN => n167, Z => Y(27));
   Y_tri_2_inst : TBUF_X1 port map( A => n137, EN => n167, Z => Y(2));
   Y_tri_4_inst : TBUF_X1 port map( A => n135, EN => n167, Z => Y(4));
   Y_tri_6_inst : TBUF_X1 port map( A => n133, EN => n167, Z => Y(6));
   Y_tri_8_inst : TBUF_X1 port map( A => n131, EN => n168, Z => Y(8));
   Y_tri_17_inst : TBUF_X1 port map( A => n121, EN => n168, Z => Y(17));
   Y_tri_19_inst : TBUF_X1 port map( A => n119, EN => n168, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n118, EN => n168, Z => Y(20));
   Y_tri_22_inst : TBUF_X1 port map( A => n116, EN => n168, Z => Y(22));
   Y_tri_24_inst : TBUF_X1 port map( A => n114, EN => n168, Z => Y(24));
   Y_tri_26_inst : TBUF_X1 port map( A => n112, EN => n168, Z => Y(26));
   Y_tri_28_inst : TBUF_X1 port map( A => n110, EN => n168, Z => Y(28));
   Y_tri_0_inst : TBUF_X1 port map( A => n139, EN => n168, Z => Y(0));
   Y_tri_1_inst : TBUF_X1 port map( A => n138, EN => n168, Z => Y(1));
   Y_tri_10_inst : TBUF_X1 port map( A => n128, EN => n168, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n127, EN => n168, Z => Y(11));
   Y_tri_31_inst : TBUF_X1 port map( A => n107, EN => n167, Z => Y(31));
   Y_tri_29_inst : TBUF_X1 port map( A => n109, EN => n167, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n108, EN => n167, Z => Y(30));
   U1 : BUF_X1 port map( A => n23, Z => n168);
   U2 : BUF_X1 port map( A => n23, Z => n167);
   U3 : BUF_X1 port map( A => n9, Z => n162);
   U4 : BUF_X1 port map( A => n9, Z => n161);
   U5 : BUF_X1 port map( A => n10, Z => n159);
   U6 : BUF_X1 port map( A => n10, Z => n158);
   U7 : BUF_X1 port map( A => n9, Z => n163);
   U8 : BUF_X1 port map( A => n10, Z => n160);
   U9 : BUF_X1 port map( A => n23, Z => n169);
   U10 : BUF_X1 port map( A => n12, Z => n153);
   U11 : BUF_X1 port map( A => n12, Z => n152);
   U12 : NOR2_X1 port map( A1 => n77, A2 => n4, ZN => n10);
   U13 : NOR2_X1 port map( A1 => n77, A2 => n5, ZN => n9);
   U14 : BUF_X1 port map( A => n13, Z => n150);
   U15 : BUF_X1 port map( A => n13, Z => n149);
   U16 : BUF_X1 port map( A => n11, Z => n156);
   U17 : BUF_X1 port map( A => n8, Z => n165);
   U18 : BUF_X1 port map( A => n11, Z => n155);
   U19 : BUF_X1 port map( A => n8, Z => n164);
   U20 : BUF_X1 port map( A => n12, Z => n154);
   U21 : BUF_X1 port map( A => n13, Z => n151);
   U22 : BUF_X1 port map( A => n11, Z => n157);
   U23 : BUF_X1 port map( A => n8, Z => n166);
   U24 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n23);
   U25 : NOR3_X1 port map( A1 => sel(1), A2 => sel(2), A3 => n77, ZN => n13);
   U26 : NOR3_X1 port map( A1 => sel(1), A2 => sel(2), A3 => sel(0), ZN => n12)
                           ;
   U27 : NOR2_X1 port map( A1 => n5, A2 => sel(0), ZN => n11);
   U28 : NOR2_X1 port map( A1 => n4, A2 => sel(0), ZN => n8);
   U29 : INV_X1 port map( A => sel(1), ZN => n5);
   U30 : INV_X1 port map( A => sel(0), ZN => n77);
   U31 : INV_X1 port map( A => sel(2), ZN => n4);
   U32 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => n108);
   U33 : AOI222_X1 port map( A1 => E(30), A2 => n164, B1 => D(30), B2 => n161, 
                           C1 => F(30), C2 => n158, ZN => n74);
   U34 : AOI222_X1 port map( A1 => C(30), A2 => n155, B1 => A(30), B2 => n152, 
                           C1 => B(30), C2 => n149, ZN => n73);
   U35 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n109);
   U36 : AOI222_X1 port map( A1 => E(29), A2 => n164, B1 => D(29), B2 => n161, 
                           C1 => F(29), C2 => n158, ZN => n72);
   U37 : AOI222_X1 port map( A1 => C(29), A2 => n155, B1 => A(29), B2 => n152, 
                           C1 => B(29), C2 => n149, ZN => n71);
   U38 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => n115);
   U39 : AOI222_X1 port map( A1 => E(23), A2 => n164, B1 => D(23), B2 => n161, 
                           C1 => F(23), C2 => n158, ZN => n60);
   U40 : AOI222_X1 port map( A1 => C(23), A2 => n155, B1 => A(23), B2 => n152, 
                           C1 => B(23), C2 => n149, ZN => n59);
   U41 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => n110);
   U42 : AOI222_X1 port map( A1 => E(28), A2 => n164, B1 => D(28), B2 => n161, 
                           C1 => F(28), C2 => n158, ZN => n70);
   U43 : AOI222_X1 port map( A1 => C(28), A2 => n155, B1 => A(28), B2 => n152, 
                           C1 => B(28), C2 => n149, ZN => n69);
   U44 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => n112);
   U45 : AOI222_X1 port map( A1 => E(26), A2 => n164, B1 => D(26), B2 => n161, 
                           C1 => F(26), C2 => n158, ZN => n66);
   U46 : AOI222_X1 port map( A1 => C(26), A2 => n155, B1 => A(26), B2 => n152, 
                           C1 => B(26), C2 => n149, ZN => n65);
   U47 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n114);
   U48 : AOI222_X1 port map( A1 => E(24), A2 => n164, B1 => D(24), B2 => n161, 
                           C1 => F(24), C2 => n158, ZN => n62);
   U49 : AOI222_X1 port map( A1 => C(24), A2 => n155, B1 => A(24), B2 => n152, 
                           C1 => B(24), C2 => n149, ZN => n61);
   U50 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => n111);
   U51 : AOI222_X1 port map( A1 => E(27), A2 => n164, B1 => D(27), B2 => n161, 
                           C1 => F(27), C2 => n158, ZN => n68);
   U52 : AOI222_X1 port map( A1 => C(27), A2 => n155, B1 => A(27), B2 => n152, 
                           C1 => B(27), C2 => n149, ZN => n67);
   U53 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n113);
   U54 : AOI222_X1 port map( A1 => E(25), A2 => n164, B1 => D(25), B2 => n161, 
                           C1 => F(25), C2 => n158, ZN => n64);
   U55 : AOI222_X1 port map( A1 => C(25), A2 => n155, B1 => A(25), B2 => n152, 
                           C1 => B(25), C2 => n149, ZN => n63);
   U56 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n138);
   U57 : AOI222_X1 port map( A1 => E(1), A2 => n166, B1 => D(1), B2 => n163, C1
                           => F(1), C2 => n160, ZN => n15);
   U58 : AOI222_X1 port map( A1 => C(1), A2 => n157, B1 => A(1), B2 => n154, C1
                           => B(1), C2 => n151, ZN => n14);
   U59 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => n139);
   U60 : AOI222_X1 port map( A1 => E(0), A2 => n166, B1 => D(0), B2 => n163, C1
                           => F(0), C2 => n160, ZN => n7);
   U61 : AOI222_X1 port map( A1 => C(0), A2 => n157, B1 => A(0), B2 => n154, C1
                           => B(0), C2 => n151, ZN => n6);
   U62 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n133);
   U63 : AOI222_X1 port map( A1 => E(6), A2 => n166, B1 => D(6), B2 => n163, C1
                           => F(6), C2 => n160, ZN => n26);
   U64 : AOI222_X1 port map( A1 => C(6), A2 => n157, B1 => A(6), B2 => n154, C1
                           => B(6), C2 => n151, ZN => n25);
   U65 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n135);
   U66 : AOI222_X1 port map( A1 => E(4), A2 => n166, B1 => D(4), B2 => n163, C1
                           => F(4), C2 => n160, ZN => n21);
   U67 : AOI222_X1 port map( A1 => C(4), A2 => n157, B1 => A(4), B2 => n154, C1
                           => B(4), C2 => n151, ZN => n20);
   U68 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n137);
   U69 : AOI222_X1 port map( A1 => E(2), A2 => n166, B1 => D(2), B2 => n163, C1
                           => F(2), C2 => n160, ZN => n17);
   U70 : AOI222_X1 port map( A1 => C(2), A2 => n157, B1 => A(2), B2 => n154, C1
                           => B(2), C2 => n151, ZN => n16);
   U71 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => n132);
   U72 : AOI222_X1 port map( A1 => E(7), A2 => n166, B1 => D(7), B2 => n163, C1
                           => F(7), C2 => n160, ZN => n28);
   U73 : AOI222_X1 port map( A1 => C(7), A2 => n157, B1 => A(7), B2 => n154, C1
                           => B(7), C2 => n151, ZN => n27);
   U74 : NAND2_X1 port map( A1 => n22, A2 => n24, ZN => n134);
   U75 : AOI222_X1 port map( A1 => E(5), A2 => n166, B1 => D(5), B2 => n163, C1
                           => F(5), C2 => n160, ZN => n24);
   U76 : AOI222_X1 port map( A1 => C(5), A2 => n157, B1 => A(5), B2 => n154, C1
                           => B(5), C2 => n151, ZN => n22);
   U77 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n136);
   U78 : AOI222_X1 port map( A1 => E(3), A2 => n166, B1 => D(3), B2 => n163, C1
                           => F(3), C2 => n160, ZN => n19);
   U79 : AOI222_X1 port map( A1 => C(3), A2 => n157, B1 => A(3), B2 => n154, C1
                           => B(3), C2 => n151, ZN => n18);
   U80 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => n107);
   U81 : AOI222_X1 port map( A1 => E(31), A2 => n164, B1 => D(31), B2 => n161, 
                           C1 => F(31), C2 => n158, ZN => n76);
   U82 : AOI222_X1 port map( A1 => C(31), A2 => n155, B1 => A(31), B2 => n152, 
                           C1 => B(31), C2 => n149, ZN => n75);
   U83 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n117);
   U84 : AOI222_X1 port map( A1 => E(21), A2 => n164, B1 => D(21), B2 => n161, 
                           C1 => F(21), C2 => n158, ZN => n56);
   U85 : AOI222_X1 port map( A1 => C(21), A2 => n155, B1 => A(21), B2 => n152, 
                           C1 => B(21), C2 => n149, ZN => n55);
   U86 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n120);
   U87 : AOI222_X1 port map( A1 => E(18), A2 => n165, B1 => D(18), B2 => n162, 
                           C1 => F(18), C2 => n159, ZN => n50);
   U88 : AOI222_X1 port map( A1 => C(18), A2 => n156, B1 => A(18), B2 => n153, 
                           C1 => B(18), C2 => n150, ZN => n49);
   U89 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n122);
   U90 : AOI222_X1 port map( A1 => E(16), A2 => n165, B1 => D(16), B2 => n162, 
                           C1 => F(16), C2 => n159, ZN => n46);
   U91 : AOI222_X1 port map( A1 => C(16), A2 => n156, B1 => A(16), B2 => n153, 
                           C1 => B(16), C2 => n150, ZN => n45);
   U92 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n123);
   U93 : AOI222_X1 port map( A1 => E(15), A2 => n165, B1 => D(15), B2 => n162, 
                           C1 => F(15), C2 => n159, ZN => n44);
   U94 : AOI222_X1 port map( A1 => C(15), A2 => n156, B1 => A(15), B2 => n153, 
                           C1 => B(15), C2 => n150, ZN => n43);
   U95 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n124);
   U96 : AOI222_X1 port map( A1 => E(14), A2 => n165, B1 => D(14), B2 => n162, 
                           C1 => F(14), C2 => n159, ZN => n42);
   U97 : AOI222_X1 port map( A1 => C(14), A2 => n156, B1 => A(14), B2 => n153, 
                           C1 => B(14), C2 => n150, ZN => n41);
   U98 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n125);
   U99 : AOI222_X1 port map( A1 => E(13), A2 => n165, B1 => D(13), B2 => n162, 
                           C1 => F(13), C2 => n159, ZN => n40);
   U100 : AOI222_X1 port map( A1 => C(13), A2 => n156, B1 => A(13), B2 => n153,
                           C1 => B(13), C2 => n150, ZN => n39);
   U101 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => n126);
   U102 : AOI222_X1 port map( A1 => E(12), A2 => n165, B1 => D(12), B2 => n162,
                           C1 => F(12), C2 => n159, ZN => n38);
   U103 : AOI222_X1 port map( A1 => C(12), A2 => n156, B1 => A(12), B2 => n153,
                           C1 => B(12), C2 => n150, ZN => n37);
   U104 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => n127);
   U105 : AOI222_X1 port map( A1 => E(11), A2 => n165, B1 => D(11), B2 => n162,
                           C1 => F(11), C2 => n159, ZN => n36);
   U106 : AOI222_X1 port map( A1 => C(11), A2 => n156, B1 => A(11), B2 => n153,
                           C1 => B(11), C2 => n150, ZN => n35);
   U107 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => n128);
   U108 : AOI222_X1 port map( A1 => E(10), A2 => n165, B1 => D(10), B2 => n162,
                           C1 => F(10), C2 => n159, ZN => n34);
   U109 : AOI222_X1 port map( A1 => C(10), A2 => n156, B1 => A(10), B2 => n153,
                           C1 => B(10), C2 => n150, ZN => n33);
   U110 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n116);
   U111 : AOI222_X1 port map( A1 => E(22), A2 => n164, B1 => D(22), B2 => n161,
                           C1 => F(22), C2 => n158, ZN => n58);
   U112 : AOI222_X1 port map( A1 => C(22), A2 => n155, B1 => A(22), B2 => n152,
                           C1 => B(22), C2 => n149, ZN => n57);
   U113 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n118);
   U114 : AOI222_X1 port map( A1 => E(20), A2 => n164, B1 => D(20), B2 => n161,
                           C1 => F(20), C2 => n158, ZN => n54);
   U115 : AOI222_X1 port map( A1 => C(20), A2 => n155, B1 => A(20), B2 => n152,
                           C1 => B(20), C2 => n149, ZN => n53);
   U116 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => n119);
   U117 : AOI222_X1 port map( A1 => E(19), A2 => n165, B1 => D(19), B2 => n162,
                           C1 => F(19), C2 => n159, ZN => n52);
   U118 : AOI222_X1 port map( A1 => C(19), A2 => n156, B1 => A(19), B2 => n153,
                           C1 => B(19), C2 => n150, ZN => n51);
   U119 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => n121);
   U120 : AOI222_X1 port map( A1 => E(17), A2 => n165, B1 => D(17), B2 => n162,
                           C1 => F(17), C2 => n159, ZN => n48);
   U121 : AOI222_X1 port map( A1 => C(17), A2 => n156, B1 => A(17), B2 => n153,
                           C1 => B(17), C2 => n150, ZN => n47);
   U122 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => n131);
   U123 : AOI222_X1 port map( A1 => E(8), A2 => n165, B1 => D(8), B2 => n162, 
                           C1 => F(8), C2 => n159, ZN => n30);
   U124 : AOI222_X1 port map( A1 => C(8), A2 => n156, B1 => A(8), B2 => n153, 
                           C1 => B(8), C2 => n150, ZN => n29);
   U125 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => n129);
   U126 : AOI222_X1 port map( A1 => E(9), A2 => n165, B1 => D(9), B2 => n162, 
                           C1 => F(9), C2 => n159, ZN => n32);
   U127 : AOI222_X1 port map( A1 => C(9), A2 => n156, B1 => A(9), B2 => n153, 
                           C1 => B(9), C2 => n150, ZN => n31);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity ff_0 is

   port( clk, rst, d_in : in std_logic;  d_out : out std_logic);

end ff_0;

architecture SYN_behav of ff_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, n1 : std_logic;

begin
   
   d_out_reg : DFF_X1 port map( D => N2, CK => clk, Q => d_out, QN => n1);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in, ZN => N2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_4 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_4;

architecture SYN_behav of reg_N32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U4 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U5 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U6 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U7 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U8 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U9 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U10 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U11 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U12 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U13 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U14 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U15 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U16 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U17 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U18 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U19 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U20 : BUF_X1 port map( A => rst, Z => n68);
   U21 : BUF_X1 port map( A => rst, Z => n69);
   U22 : BUF_X1 port map( A => rst, Z => n70);
   U23 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U24 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U25 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U26 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U27 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U28 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U29 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U30 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U31 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U32 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U33 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U34 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U35 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U36 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U37 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity PC_incr is

   port( PC : in std_logic_vector (31 downto 0);  NPC : out std_logic_vector 
         (31 downto 0));

end PC_incr;

architecture SYN_behav of PC_incr is

   component PC_incr_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal net227480, n4, n5, n6 : std_logic;

begin
   
   n4 <= '0';
   n5 <= '1';
   n6 <= '0';
   add_14 : PC_incr_DW01_add_1 port map( A(31) => PC(31), A(30) => PC(30), 
                           A(29) => PC(29), A(28) => PC(28), A(27) => PC(27), 
                           A(26) => PC(26), A(25) => PC(25), A(24) => PC(24), 
                           A(23) => PC(23), A(22) => PC(22), A(21) => PC(21), 
                           A(20) => PC(20), A(19) => PC(19), A(18) => PC(18), 
                           A(17) => PC(17), A(16) => PC(16), A(15) => PC(15), 
                           A(14) => PC(14), A(13) => PC(13), A(12) => PC(12), 
                           A(11) => PC(11), A(10) => PC(10), A(9) => PC(9), 
                           A(8) => PC(8), A(7) => PC(7), A(6) => PC(6), A(5) =>
                           PC(5), A(4) => PC(4), A(3) => PC(3), A(2) => PC(2), 
                           A(1) => PC(1), A(0) => PC(0), B(31) => n6, B(30) => 
                           n6, B(29) => n6, B(28) => n6, B(27) => n6, B(26) => 
                           n6, B(25) => n6, B(24) => n6, B(23) => n6, B(22) => 
                           n6, B(21) => n6, B(20) => n6, B(19) => n6, B(18) => 
                           n6, B(17) => n6, B(16) => n6, B(15) => n6, B(14) => 
                           n6, B(13) => n6, B(12) => n6, B(11) => n6, B(10) => 
                           n6, B(9) => n6, B(8) => n6, B(7) => n6, B(6) => n6, 
                           B(5) => n6, B(4) => n6, B(3) => n6, B(2) => n5, B(1)
                           => n4, B(0) => n4, CI => n6, SUM(31) => NPC(31), 
                           SUM(30) => NPC(30), SUM(29) => NPC(29), SUM(28) => 
                           NPC(28), SUM(27) => NPC(27), SUM(26) => NPC(26), 
                           SUM(25) => NPC(25), SUM(24) => NPC(24), SUM(23) => 
                           NPC(23), SUM(22) => NPC(22), SUM(21) => NPC(21), 
                           SUM(20) => NPC(20), SUM(19) => NPC(19), SUM(18) => 
                           NPC(18), SUM(17) => NPC(17), SUM(16) => NPC(16), 
                           SUM(15) => NPC(15), SUM(14) => NPC(14), SUM(13) => 
                           NPC(13), SUM(12) => NPC(12), SUM(11) => NPC(11), 
                           SUM(10) => NPC(10), SUM(9) => NPC(9), SUM(8) => 
                           NPC(8), SUM(7) => NPC(7), SUM(6) => NPC(6), SUM(5) 
                           => NPC(5), SUM(4) => NPC(4), SUM(3) => NPC(3), 
                           SUM(2) => NPC(2), SUM(1) => NPC(1), SUM(0) => NPC(0)
                           , CO => net227480);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_en_N32 is

   port( clk, rst, en : in std_logic;  d_in : in std_logic_vector (31 downto 0)
         ;  d_out : out std_logic_vector (31 downto 0));

end reg_en_N32;

architecture SYN_behav of reg_en_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, net227477, net227478, net227479, n34, n35, n36, n66, 
      n67, n68, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => n100, CK => clk, Q => d_out(31), 
                           QN => net227479);
   d_out_reg_30_inst : DFF_X1 port map( D => n99, CK => clk, Q => d_out(30), QN
                           => net227478);
   d_out_reg_29_inst : DFF_X1 port map( D => n98, CK => clk, Q => d_out(29), QN
                           => net227477);
   d_out_reg_28_inst : DFF_X1 port map( D => n97, CK => clk, Q => d_out(28), QN
                           => n65);
   d_out_reg_27_inst : DFF_X1 port map( D => n96, CK => clk, Q => d_out(27), QN
                           => n64);
   d_out_reg_26_inst : DFF_X1 port map( D => n95, CK => clk, Q => d_out(26), QN
                           => n63);
   d_out_reg_25_inst : DFF_X1 port map( D => n94, CK => clk, Q => d_out(25), QN
                           => n62);
   d_out_reg_24_inst : DFF_X1 port map( D => n93, CK => clk, Q => d_out(24), QN
                           => n61);
   d_out_reg_23_inst : DFF_X1 port map( D => n92, CK => clk, Q => d_out(23), QN
                           => n60);
   d_out_reg_22_inst : DFF_X1 port map( D => n91, CK => clk, Q => d_out(22), QN
                           => n59);
   d_out_reg_21_inst : DFF_X1 port map( D => n90, CK => clk, Q => d_out(21), QN
                           => n58);
   d_out_reg_20_inst : DFF_X1 port map( D => n89, CK => clk, Q => d_out(20), QN
                           => n57);
   d_out_reg_19_inst : DFF_X1 port map( D => n88, CK => clk, Q => d_out(19), QN
                           => n56);
   d_out_reg_18_inst : DFF_X1 port map( D => n87, CK => clk, Q => d_out(18), QN
                           => n55);
   d_out_reg_17_inst : DFF_X1 port map( D => n86, CK => clk, Q => d_out(17), QN
                           => n54);
   d_out_reg_16_inst : DFF_X1 port map( D => n85, CK => clk, Q => d_out(16), QN
                           => n53);
   d_out_reg_15_inst : DFF_X1 port map( D => n84, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => n83, CK => clk, Q => d_out(14), QN
                           => n51);
   d_out_reg_13_inst : DFF_X1 port map( D => n82, CK => clk, Q => d_out(13), QN
                           => n50);
   d_out_reg_12_inst : DFF_X1 port map( D => n81, CK => clk, Q => d_out(12), QN
                           => n49);
   d_out_reg_11_inst : DFF_X1 port map( D => n80, CK => clk, Q => d_out(11), QN
                           => n48);
   d_out_reg_10_inst : DFF_X1 port map( D => n79, CK => clk, Q => d_out(10), QN
                           => n47);
   d_out_reg_9_inst : DFF_X1 port map( D => n78, CK => clk, Q => d_out(9), QN 
                           => n46);
   d_out_reg_8_inst : DFF_X1 port map( D => n77, CK => clk, Q => d_out(8), QN 
                           => n45);
   d_out_reg_7_inst : DFF_X1 port map( D => n76, CK => clk, Q => d_out(7), QN 
                           => n44);
   d_out_reg_6_inst : DFF_X1 port map( D => n75, CK => clk, Q => d_out(6), QN 
                           => n43);
   d_out_reg_5_inst : DFF_X1 port map( D => n74, CK => clk, Q => d_out(5), QN 
                           => n42);
   d_out_reg_4_inst : DFF_X1 port map( D => n73, CK => clk, Q => d_out(4), QN 
                           => n41);
   d_out_reg_3_inst : DFF_X1 port map( D => n72, CK => clk, Q => d_out(3), QN 
                           => n40);
   d_out_reg_2_inst : DFF_X1 port map( D => n71, CK => clk, Q => d_out(2), QN 
                           => n39);
   d_out_reg_1_inst : DFF_X1 port map( D => n70, CK => clk, Q => d_out(1), QN 
                           => n38);
   d_out_reg_0_inst : DFF_X1 port map( D => n69, CK => clk, Q => d_out(0), QN 
                           => n37);
   U3 : BUF_X1 port map( A => n35, Z => n131);
   U4 : BUF_X1 port map( A => n35, Z => n130);
   U5 : BUF_X1 port map( A => n35, Z => n132);
   U6 : BUF_X1 port map( A => n34, Z => n135);
   U7 : BUF_X1 port map( A => n34, Z => n133);
   U8 : BUF_X1 port map( A => n34, Z => n134);
   U9 : NAND2_X1 port map( A1 => rst, A2 => n133, ZN => n35);
   U10 : OAI22_X1 port map( A1 => net227477, A2 => n135, B1 => n132, B2 => n66,
                           ZN => n98);
   U11 : INV_X1 port map( A => d_in(29), ZN => n66);
   U12 : OAI22_X1 port map( A1 => net227478, A2 => n135, B1 => n132, B2 => n36,
                           ZN => n99);
   U13 : INV_X1 port map( A => d_in(30), ZN => n36);
   U14 : OAI22_X1 port map( A1 => n60, A2 => n135, B1 => n132, B2 => n104, ZN 
                           => n92);
   U15 : INV_X1 port map( A => d_in(23), ZN => n104);
   U16 : OAI22_X1 port map( A1 => n61, A2 => n135, B1 => n132, B2 => n103, ZN 
                           => n93);
   U17 : INV_X1 port map( A => d_in(24), ZN => n103);
   U18 : OAI22_X1 port map( A1 => n62, A2 => n135, B1 => n132, B2 => n102, ZN 
                           => n94);
   U19 : INV_X1 port map( A => d_in(25), ZN => n102);
   U20 : OAI22_X1 port map( A1 => n63, A2 => n135, B1 => n132, B2 => n101, ZN 
                           => n95);
   U21 : INV_X1 port map( A => d_in(26), ZN => n101);
   U22 : OAI22_X1 port map( A1 => n64, A2 => n135, B1 => n132, B2 => n68, ZN =>
                           n96);
   U23 : INV_X1 port map( A => d_in(27), ZN => n68);
   U24 : OAI22_X1 port map( A1 => n65, A2 => n135, B1 => n132, B2 => n67, ZN =>
                           n97);
   U25 : INV_X1 port map( A => d_in(28), ZN => n67);
   U26 : OAI22_X1 port map( A1 => net227479, A2 => n133, B1 => n130, B2 => n128
                           , ZN => n100);
   U27 : INV_X1 port map( A => d_in(31), ZN => n128);
   U28 : OAI22_X1 port map( A1 => n37, A2 => n133, B1 => n130, B2 => n127, ZN 
                           => n69);
   U29 : INV_X1 port map( A => d_in(0), ZN => n127);
   U30 : OAI22_X1 port map( A1 => n38, A2 => n133, B1 => n130, B2 => n126, ZN 
                           => n70);
   U31 : INV_X1 port map( A => d_in(1), ZN => n126);
   U32 : OAI22_X1 port map( A1 => n39, A2 => n133, B1 => n130, B2 => n125, ZN 
                           => n71);
   U33 : INV_X1 port map( A => d_in(2), ZN => n125);
   U34 : OAI22_X1 port map( A1 => n40, A2 => n133, B1 => n130, B2 => n124, ZN 
                           => n72);
   U35 : INV_X1 port map( A => d_in(3), ZN => n124);
   U36 : OAI22_X1 port map( A1 => n41, A2 => n133, B1 => n130, B2 => n123, ZN 
                           => n73);
   U37 : INV_X1 port map( A => d_in(4), ZN => n123);
   U38 : OAI22_X1 port map( A1 => n42, A2 => n133, B1 => n130, B2 => n122, ZN 
                           => n74);
   U39 : INV_X1 port map( A => d_in(5), ZN => n122);
   U40 : OAI22_X1 port map( A1 => n43, A2 => n133, B1 => n130, B2 => n121, ZN 
                           => n75);
   U41 : INV_X1 port map( A => d_in(6), ZN => n121);
   U42 : OAI22_X1 port map( A1 => n44, A2 => n133, B1 => n130, B2 => n120, ZN 
                           => n76);
   U43 : INV_X1 port map( A => d_in(7), ZN => n120);
   U44 : OAI22_X1 port map( A1 => n45, A2 => n133, B1 => n130, B2 => n119, ZN 
                           => n77);
   U45 : INV_X1 port map( A => d_in(8), ZN => n119);
   U46 : OAI22_X1 port map( A1 => n46, A2 => n133, B1 => n130, B2 => n118, ZN 
                           => n78);
   U47 : INV_X1 port map( A => d_in(9), ZN => n118);
   U48 : OAI22_X1 port map( A1 => n47, A2 => n134, B1 => n130, B2 => n117, ZN 
                           => n79);
   U49 : INV_X1 port map( A => d_in(10), ZN => n117);
   U50 : OAI22_X1 port map( A1 => n48, A2 => n134, B1 => n131, B2 => n116, ZN 
                           => n80);
   U51 : INV_X1 port map( A => d_in(11), ZN => n116);
   U52 : OAI22_X1 port map( A1 => n49, A2 => n134, B1 => n131, B2 => n115, ZN 
                           => n81);
   U53 : INV_X1 port map( A => d_in(12), ZN => n115);
   U54 : OAI22_X1 port map( A1 => n50, A2 => n134, B1 => n131, B2 => n114, ZN 
                           => n82);
   U55 : INV_X1 port map( A => d_in(13), ZN => n114);
   U56 : OAI22_X1 port map( A1 => n51, A2 => n134, B1 => n131, B2 => n113, ZN 
                           => n83);
   U57 : INV_X1 port map( A => d_in(14), ZN => n113);
   U58 : OAI22_X1 port map( A1 => n52, A2 => n134, B1 => n131, B2 => n112, ZN 
                           => n84);
   U59 : INV_X1 port map( A => d_in(15), ZN => n112);
   U60 : OAI22_X1 port map( A1 => n53, A2 => n134, B1 => n131, B2 => n111, ZN 
                           => n85);
   U61 : INV_X1 port map( A => d_in(16), ZN => n111);
   U62 : OAI22_X1 port map( A1 => n54, A2 => n134, B1 => n131, B2 => n110, ZN 
                           => n86);
   U63 : INV_X1 port map( A => d_in(17), ZN => n110);
   U64 : OAI22_X1 port map( A1 => n55, A2 => n134, B1 => n131, B2 => n109, ZN 
                           => n87);
   U65 : INV_X1 port map( A => d_in(18), ZN => n109);
   U66 : OAI22_X1 port map( A1 => n56, A2 => n134, B1 => n131, B2 => n108, ZN 
                           => n88);
   U67 : INV_X1 port map( A => d_in(19), ZN => n108);
   U68 : OAI22_X1 port map( A1 => n57, A2 => n134, B1 => n131, B2 => n107, ZN 
                           => n89);
   U69 : INV_X1 port map( A => d_in(20), ZN => n107);
   U70 : OAI22_X1 port map( A1 => n58, A2 => n134, B1 => n131, B2 => n106, ZN 
                           => n90);
   U71 : INV_X1 port map( A => d_in(21), ZN => n106);
   U72 : OAI22_X1 port map( A1 => n59, A2 => n135, B1 => n131, B2 => n105, ZN 
                           => n91);
   U73 : INV_X1 port map( A => d_in(22), ZN => n105);
   U74 : NAND2_X1 port map( A1 => n129, A2 => rst, ZN => n34);
   U75 : INV_X1 port map( A => en, ZN => n129);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_1;

architecture SYN_struct of MUX21_GENERIC_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   M_0 : MUX21_90 port map( A => A(0), B => B(0), S => n4, Y => Y(0));
   M_1 : MUX21_89 port map( A => A(1), B => B(1), S => n4, Y => Y(1));
   M_2 : MUX21_88 port map( A => A(2), B => B(2), S => n4, Y => Y(2));
   M_3 : MUX21_87 port map( A => A(3), B => B(3), S => n4, Y => Y(3));
   M_4 : MUX21_86 port map( A => A(4), B => B(4), S => n4, Y => Y(4));
   M_5 : MUX21_85 port map( A => A(5), B => B(5), S => n4, Y => Y(5));
   M_6 : MUX21_84 port map( A => A(6), B => B(6), S => n4, Y => Y(6));
   M_7 : MUX21_83 port map( A => A(7), B => B(7), S => n4, Y => Y(7));
   M_8 : MUX21_82 port map( A => A(8), B => B(8), S => n4, Y => Y(8));
   M_9 : MUX21_81 port map( A => A(9), B => B(9), S => n4, Y => Y(9));
   M_10 : MUX21_80 port map( A => A(10), B => B(10), S => n4, Y => Y(10));
   M_11 : MUX21_79 port map( A => A(11), B => B(11), S => n4, Y => Y(11));
   M_12 : MUX21_78 port map( A => A(12), B => B(12), S => n5, Y => Y(12));
   M_13 : MUX21_77 port map( A => A(13), B => B(13), S => n5, Y => Y(13));
   M_14 : MUX21_76 port map( A => A(14), B => B(14), S => n5, Y => Y(14));
   M_15 : MUX21_75 port map( A => A(15), B => B(15), S => n5, Y => Y(15));
   M_16 : MUX21_74 port map( A => A(16), B => B(16), S => n5, Y => Y(16));
   M_17 : MUX21_73 port map( A => A(17), B => B(17), S => n5, Y => Y(17));
   M_18 : MUX21_72 port map( A => A(18), B => B(18), S => n5, Y => Y(18));
   M_19 : MUX21_71 port map( A => A(19), B => B(19), S => n5, Y => Y(19));
   M_20 : MUX21_70 port map( A => A(20), B => B(20), S => n5, Y => Y(20));
   M_21 : MUX21_69 port map( A => A(21), B => B(21), S => n5, Y => Y(21));
   M_22 : MUX21_68 port map( A => A(22), B => B(22), S => n5, Y => Y(22));
   M_23 : MUX21_67 port map( A => A(23), B => B(23), S => n5, Y => Y(23));
   M_24 : MUX21_66 port map( A => A(24), B => B(24), S => n6, Y => Y(24));
   M_25 : MUX21_65 port map( A => A(25), B => B(25), S => n6, Y => Y(25));
   M_26 : MUX21_64 port map( A => A(26), B => B(26), S => n6, Y => Y(26));
   M_27 : MUX21_63 port map( A => A(27), B => B(27), S => n6, Y => Y(27));
   M_28 : MUX21_62 port map( A => A(28), B => B(28), S => n6, Y => Y(28));
   M_29 : MUX21_61 port map( A => A(29), B => B(29), S => n6, Y => Y(29));
   M_30 : MUX21_31 port map( A => A(30), B => B(30), S => n6, Y => Y(30));
   M_31 : MUX21_30 port map( A => A(31), B => B(31), S => n6, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n4);
   U2 : BUF_X1 port map( A => SEL, Z => n5);
   U3 : BUF_X1 port map( A => SEL, Z => n6);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_5 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_5;

architecture SYN_behav of reg_N32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U7 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U8 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U9 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U10 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U11 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U12 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U13 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U14 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U15 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U16 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U17 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U20 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U21 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U22 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U23 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U24 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U25 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U26 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U27 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U28 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U29 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U30 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U31 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U32 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U33 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U34 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U35 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_6 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_6;

architecture SYN_behav of reg_N32_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U10 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U11 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U14 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U15 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U16 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U17 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U18 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U19 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U20 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U21 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U22 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U23 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U24 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U25 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U26 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U27 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U28 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U29 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U30 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U31 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U32 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U33 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U34 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U35 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U36 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U37 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_10 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_10;

architecture SYN_behav of reg_N32_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U4 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U5 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U6 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U7 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U8 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U9 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U10 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U11 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U12 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U13 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U14 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U15 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U16 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U17 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U18 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U19 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U20 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U21 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U22 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U23 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U24 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U25 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U26 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U27 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U28 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U29 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U30 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U31 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U32 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U33 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U34 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);
   U35 : BUF_X1 port map( A => rst, Z => n68);
   U36 : BUF_X1 port map( A => rst, Z => n69);
   U37 : BUF_X1 port map( A => rst, Z => n70);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity MUX21_GENERIC_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_0;

architecture SYN_struct of MUX21_GENERIC_N32_0 is

   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_0 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_217 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_216 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_215 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   M_4 : MUX21_214 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   M_5 : MUX21_213 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   M_6 : MUX21_212 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   M_7 : MUX21_211 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   M_8 : MUX21_210 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   M_9 : MUX21_209 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   M_10 : MUX21_208 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   M_11 : MUX21_207 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   M_12 : MUX21_206 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   M_13 : MUX21_205 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   M_14 : MUX21_204 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   M_15 : MUX21_203 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   M_16 : MUX21_202 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   M_17 : MUX21_201 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   M_18 : MUX21_200 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   M_19 : MUX21_199 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   M_20 : MUX21_198 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   M_21 : MUX21_197 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   M_22 : MUX21_196 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   M_23 : MUX21_195 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   M_24 : MUX21_194 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   M_25 : MUX21_193 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   M_26 : MUX21_192 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   M_27 : MUX21_191 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   M_28 : MUX21_190 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   M_29 : MUX21_189 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   M_30 : MUX21_188 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   M_31 : MUX21_187 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity sign_ext_Nstart26_Nend32 is

   port( Ain : in std_logic_vector (25 downto 0);  Aout : out std_logic_vector 
         (31 downto 0));

end sign_ext_Nstart26_Nend32;

architecture SYN_behav of sign_ext_Nstart26_Nend32 is

begin
   Aout <= ( Ain(25), Ain(25), Ain(25), Ain(25), Ain(25), Ain(25), Ain(25), 
      Ain(24), Ain(23), Ain(22), Ain(21), Ain(20), Ain(19), Ain(18), Ain(17), 
      Ain(16), Ain(15), Ain(14), Ain(13), Ain(12), Ain(11), Ain(10), Ain(9), 
      Ain(8), Ain(7), Ain(6), Ain(5), Ain(4), Ain(3), Ain(2), Ain(1), Ain(0) );

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity sign_ext_Nstart16_Nend32 is

   port( Ain : in std_logic_vector (15 downto 0);  Aout : out std_logic_vector 
         (31 downto 0));

end sign_ext_Nstart16_Nend32;

architecture SYN_behav of sign_ext_Nstart16_Nend32 is

begin
   Aout <= ( Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), 
      Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), Ain(15), 
      Ain(15), Ain(15), Ain(14), Ain(13), Ain(12), Ain(11), Ain(10), Ain(9), 
      Ain(8), Ain(7), Ain(6), Ain(5), Ain(4), Ain(3), Ain(2), Ain(1), Ain(0) );

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_13 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_13;

architecture SYN_behav of reg_N32_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity w_reg_file_M8_N8_F4_Nbit32 is

   port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  datain : in 
         std_logic_vector (31 downto 0);  out1, out2 : out std_logic_vector (31
         downto 0);  call, ret : in std_logic;  spill, fill : out std_logic;  
         to_mem : out std_logic_vector (31 downto 0);  from_mem : in 
         std_logic_vector (31 downto 0));

end w_reg_file_M8_N8_F4_Nbit32;

architecture SYN_behav of w_reg_file_M8_N8_F4_Nbit32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0
      port( A : in std_logic_vector (5 downto 0);  SUM : out std_logic_vector 
            (5 downto 0));
   end component;
   
   component w_reg_file_M8_N8_F4_Nbit32_DW01_add_1
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   component w_reg_file_M8_N8_F4_Nbit32_DW01_add_0
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal registers_0_31_port, registers_0_30_port, registers_0_29_port, 
      registers_0_28_port, registers_0_27_port, registers_0_26_port, 
      registers_0_25_port, registers_0_24_port, registers_0_23_port, 
      registers_0_22_port, registers_0_21_port, registers_0_20_port, 
      registers_0_19_port, registers_0_18_port, registers_0_17_port, 
      registers_0_16_port, registers_0_15_port, registers_0_14_port, 
      registers_0_13_port, registers_0_12_port, registers_0_11_port, 
      registers_0_10_port, registers_0_9_port, registers_0_8_port, 
      registers_0_7_port, registers_0_6_port, registers_0_5_port, 
      registers_0_4_port, registers_0_3_port, registers_0_2_port, 
      registers_0_1_port, registers_0_0_port, registers_1_31_port, 
      registers_1_30_port, registers_1_29_port, registers_1_28_port, 
      registers_1_27_port, registers_1_26_port, registers_1_25_port, 
      registers_1_24_port, registers_1_23_port, registers_1_22_port, 
      registers_1_21_port, registers_1_20_port, registers_1_19_port, 
      registers_1_18_port, registers_1_17_port, registers_1_16_port, 
      registers_1_15_port, registers_1_14_port, registers_1_13_port, 
      registers_1_12_port, registers_1_11_port, registers_1_10_port, 
      registers_1_9_port, registers_1_8_port, registers_1_7_port, 
      registers_1_6_port, registers_1_5_port, registers_1_4_port, 
      registers_1_3_port, registers_1_2_port, registers_1_1_port, 
      registers_1_0_port, registers_2_31_port, registers_2_30_port, 
      registers_2_29_port, registers_2_28_port, registers_2_27_port, 
      registers_2_26_port, registers_2_25_port, registers_2_24_port, 
      registers_2_23_port, registers_2_22_port, registers_2_21_port, 
      registers_2_20_port, registers_2_19_port, registers_2_18_port, 
      registers_2_17_port, registers_2_16_port, registers_2_15_port, 
      registers_2_14_port, registers_2_13_port, registers_2_12_port, 
      registers_2_11_port, registers_2_10_port, registers_2_9_port, 
      registers_2_8_port, registers_2_7_port, registers_2_6_port, 
      registers_2_5_port, registers_2_4_port, registers_2_3_port, 
      registers_2_2_port, registers_2_1_port, registers_2_0_port, 
      registers_4_31_port, registers_4_30_port, registers_4_29_port, 
      registers_4_28_port, registers_4_27_port, registers_4_26_port, 
      registers_4_25_port, registers_4_24_port, registers_4_23_port, 
      registers_4_22_port, registers_4_21_port, registers_4_20_port, 
      registers_4_19_port, registers_4_18_port, registers_4_17_port, 
      registers_4_16_port, registers_4_15_port, registers_4_14_port, 
      registers_4_13_port, registers_4_12_port, registers_4_11_port, 
      registers_4_10_port, registers_4_9_port, registers_4_8_port, 
      registers_4_7_port, registers_4_6_port, registers_4_5_port, 
      registers_4_4_port, registers_4_3_port, registers_4_2_port, 
      registers_4_1_port, registers_4_0_port, registers_5_31_port, 
      registers_5_30_port, registers_5_29_port, registers_5_28_port, 
      registers_5_27_port, registers_5_26_port, registers_5_25_port, 
      registers_5_24_port, registers_5_23_port, registers_5_22_port, 
      registers_5_21_port, registers_5_20_port, registers_5_19_port, 
      registers_5_18_port, registers_5_17_port, registers_5_16_port, 
      registers_5_15_port, registers_5_14_port, registers_5_13_port, 
      registers_5_12_port, registers_5_11_port, registers_5_10_port, 
      registers_5_9_port, registers_5_8_port, registers_5_7_port, 
      registers_5_6_port, registers_5_5_port, registers_5_4_port, 
      registers_5_3_port, registers_5_2_port, registers_5_1_port, 
      registers_5_0_port, registers_7_31_port, registers_7_30_port, 
      registers_7_29_port, registers_7_28_port, registers_7_27_port, 
      registers_7_26_port, registers_7_25_port, registers_7_24_port, 
      registers_7_23_port, registers_7_22_port, registers_7_21_port, 
      registers_7_20_port, registers_7_19_port, registers_7_18_port, 
      registers_7_17_port, registers_7_16_port, registers_7_15_port, 
      registers_7_14_port, registers_7_13_port, registers_7_12_port, 
      registers_7_11_port, registers_7_10_port, registers_7_9_port, 
      registers_7_8_port, registers_7_7_port, registers_7_6_port, 
      registers_7_5_port, registers_7_4_port, registers_7_3_port, 
      registers_7_2_port, registers_7_1_port, registers_7_0_port, 
      registers_9_31_port, registers_9_30_port, registers_9_29_port, 
      registers_9_28_port, registers_9_27_port, registers_9_26_port, 
      registers_9_25_port, registers_9_24_port, registers_9_23_port, 
      registers_9_22_port, registers_9_21_port, registers_9_20_port, 
      registers_9_19_port, registers_9_18_port, registers_9_17_port, 
      registers_9_16_port, registers_9_15_port, registers_9_14_port, 
      registers_9_13_port, registers_9_12_port, registers_9_11_port, 
      registers_9_10_port, registers_9_9_port, registers_9_8_port, 
      registers_9_7_port, registers_9_6_port, registers_9_5_port, 
      registers_9_4_port, registers_9_3_port, registers_9_2_port, 
      registers_9_1_port, registers_9_0_port, registers_10_31_port, 
      registers_10_30_port, registers_10_29_port, registers_10_28_port, 
      registers_10_27_port, registers_10_26_port, registers_10_25_port, 
      registers_10_24_port, registers_10_23_port, registers_10_22_port, 
      registers_10_21_port, registers_10_20_port, registers_10_19_port, 
      registers_10_18_port, registers_10_17_port, registers_10_16_port, 
      registers_10_15_port, registers_10_14_port, registers_10_13_port, 
      registers_10_12_port, registers_10_11_port, registers_10_10_port, 
      registers_10_9_port, registers_10_8_port, registers_10_7_port, 
      registers_10_6_port, registers_10_5_port, registers_10_4_port, 
      registers_10_3_port, registers_10_2_port, registers_10_1_port, 
      registers_10_0_port, registers_11_31_port, registers_11_30_port, 
      registers_11_29_port, registers_11_28_port, registers_11_27_port, 
      registers_11_26_port, registers_11_25_port, registers_11_24_port, 
      registers_11_23_port, registers_11_22_port, registers_11_21_port, 
      registers_11_20_port, registers_11_19_port, registers_11_18_port, 
      registers_11_17_port, registers_11_16_port, registers_11_15_port, 
      registers_11_14_port, registers_11_13_port, registers_11_12_port, 
      registers_11_11_port, registers_11_10_port, registers_11_9_port, 
      registers_11_8_port, registers_11_7_port, registers_11_6_port, 
      registers_11_5_port, registers_11_4_port, registers_11_3_port, 
      registers_11_2_port, registers_11_1_port, registers_11_0_port, 
      registers_12_31_port, registers_12_30_port, registers_12_29_port, 
      registers_12_28_port, registers_12_27_port, registers_12_26_port, 
      registers_12_25_port, registers_12_24_port, registers_12_23_port, 
      registers_12_22_port, registers_12_21_port, registers_12_20_port, 
      registers_12_19_port, registers_12_18_port, registers_12_17_port, 
      registers_12_16_port, registers_12_15_port, registers_12_14_port, 
      registers_12_13_port, registers_12_12_port, registers_12_11_port, 
      registers_12_10_port, registers_12_9_port, registers_12_8_port, 
      registers_12_7_port, registers_12_6_port, registers_12_5_port, 
      registers_12_4_port, registers_12_3_port, registers_12_2_port, 
      registers_12_1_port, registers_12_0_port, registers_15_31_port, 
      registers_15_30_port, registers_15_29_port, registers_15_28_port, 
      registers_15_27_port, registers_15_26_port, registers_15_25_port, 
      registers_15_24_port, registers_15_23_port, registers_15_22_port, 
      registers_15_21_port, registers_15_20_port, registers_15_19_port, 
      registers_15_18_port, registers_15_17_port, registers_15_16_port, 
      registers_15_15_port, registers_15_14_port, registers_15_13_port, 
      registers_15_12_port, registers_15_11_port, registers_15_10_port, 
      registers_15_9_port, registers_15_8_port, registers_15_7_port, 
      registers_15_6_port, registers_15_5_port, registers_15_4_port, 
      registers_15_3_port, registers_15_2_port, registers_15_1_port, 
      registers_15_0_port, registers_16_31_port, registers_16_30_port, 
      registers_16_29_port, registers_16_28_port, registers_16_27_port, 
      registers_16_26_port, registers_16_25_port, registers_16_24_port, 
      registers_16_23_port, registers_16_22_port, registers_16_21_port, 
      registers_16_20_port, registers_16_19_port, registers_16_18_port, 
      registers_16_17_port, registers_16_16_port, registers_16_15_port, 
      registers_16_14_port, registers_16_13_port, registers_16_12_port, 
      registers_16_11_port, registers_16_10_port, registers_16_9_port, 
      registers_16_8_port, registers_16_7_port, registers_16_6_port, 
      registers_16_5_port, registers_16_4_port, registers_16_3_port, 
      registers_16_2_port, registers_16_1_port, registers_16_0_port, 
      registers_17_31_port, registers_17_30_port, registers_17_29_port, 
      registers_17_28_port, registers_17_27_port, registers_17_26_port, 
      registers_17_25_port, registers_17_24_port, registers_17_23_port, 
      registers_17_22_port, registers_17_21_port, registers_17_20_port, 
      registers_17_19_port, registers_17_18_port, registers_17_17_port, 
      registers_17_16_port, registers_17_15_port, registers_17_14_port, 
      registers_17_13_port, registers_17_12_port, registers_17_11_port, 
      registers_17_10_port, registers_17_9_port, registers_17_8_port, 
      registers_17_7_port, registers_17_6_port, registers_17_5_port, 
      registers_17_4_port, registers_17_3_port, registers_17_2_port, 
      registers_17_1_port, registers_17_0_port, registers_18_31_port, 
      registers_18_30_port, registers_18_29_port, registers_18_28_port, 
      registers_18_27_port, registers_18_26_port, registers_18_25_port, 
      registers_18_24_port, registers_18_23_port, registers_18_22_port, 
      registers_18_21_port, registers_18_20_port, registers_18_19_port, 
      registers_18_18_port, registers_18_17_port, registers_18_16_port, 
      registers_18_15_port, registers_18_14_port, registers_18_13_port, 
      registers_18_12_port, registers_18_11_port, registers_18_10_port, 
      registers_18_9_port, registers_18_8_port, registers_18_7_port, 
      registers_18_6_port, registers_18_5_port, registers_18_4_port, 
      registers_18_3_port, registers_18_2_port, registers_18_1_port, 
      registers_18_0_port, registers_19_31_port, registers_19_30_port, 
      registers_19_29_port, registers_19_28_port, registers_19_27_port, 
      registers_19_26_port, registers_19_25_port, registers_19_24_port, 
      registers_19_23_port, registers_19_22_port, registers_19_21_port, 
      registers_19_20_port, registers_19_19_port, registers_19_18_port, 
      registers_19_17_port, registers_19_16_port, registers_19_15_port, 
      registers_19_14_port, registers_19_13_port, registers_19_12_port, 
      registers_19_11_port, registers_19_10_port, registers_19_9_port, 
      registers_19_8_port, registers_19_7_port, registers_19_6_port, 
      registers_19_5_port, registers_19_4_port, registers_19_3_port, 
      registers_19_2_port, registers_19_1_port, registers_19_0_port, 
      registers_22_31_port, registers_22_30_port, registers_22_29_port, 
      registers_22_28_port, registers_22_27_port, registers_22_26_port, 
      registers_22_25_port, registers_22_24_port, registers_22_23_port, 
      registers_22_22_port, registers_22_21_port, registers_22_20_port, 
      registers_22_19_port, registers_22_18_port, registers_22_17_port, 
      registers_22_16_port, registers_22_15_port, registers_22_14_port, 
      registers_22_13_port, registers_22_12_port, registers_22_11_port, 
      registers_22_10_port, registers_22_9_port, registers_22_8_port, 
      registers_22_7_port, registers_22_6_port, registers_22_5_port, 
      registers_22_4_port, registers_22_3_port, registers_22_2_port, 
      registers_22_1_port, registers_22_0_port, registers_23_31_port, 
      registers_23_30_port, registers_23_29_port, registers_23_28_port, 
      registers_23_27_port, registers_23_26_port, registers_23_25_port, 
      registers_23_24_port, registers_23_23_port, registers_23_22_port, 
      registers_23_21_port, registers_23_20_port, registers_23_19_port, 
      registers_23_18_port, registers_23_17_port, registers_23_16_port, 
      registers_23_15_port, registers_23_14_port, registers_23_13_port, 
      registers_23_12_port, registers_23_11_port, registers_23_10_port, 
      registers_23_9_port, registers_23_8_port, registers_23_7_port, 
      registers_23_6_port, registers_23_5_port, registers_23_4_port, 
      registers_23_3_port, registers_23_2_port, registers_23_1_port, 
      registers_23_0_port, registers_25_31_port, registers_25_30_port, 
      registers_25_29_port, registers_25_28_port, registers_25_27_port, 
      registers_25_26_port, registers_25_25_port, registers_25_24_port, 
      registers_25_23_port, registers_25_22_port, registers_25_21_port, 
      registers_25_20_port, registers_25_19_port, registers_25_18_port, 
      registers_25_17_port, registers_25_16_port, registers_25_15_port, 
      registers_25_14_port, registers_25_13_port, registers_25_12_port, 
      registers_25_11_port, registers_25_10_port, registers_25_9_port, 
      registers_25_8_port, registers_25_7_port, registers_25_6_port, 
      registers_25_5_port, registers_25_4_port, registers_25_3_port, 
      registers_25_2_port, registers_25_1_port, registers_25_0_port, 
      registers_29_31_port, registers_29_30_port, registers_29_29_port, 
      registers_29_28_port, registers_29_27_port, registers_29_26_port, 
      registers_29_25_port, registers_29_24_port, registers_29_23_port, 
      registers_29_22_port, registers_29_21_port, registers_29_20_port, 
      registers_29_19_port, registers_29_18_port, registers_29_17_port, 
      registers_29_16_port, registers_29_15_port, registers_29_14_port, 
      registers_29_13_port, registers_29_12_port, registers_29_11_port, 
      registers_29_10_port, registers_29_9_port, registers_29_8_port, 
      registers_29_7_port, registers_29_6_port, registers_29_5_port, 
      registers_29_4_port, registers_29_3_port, registers_29_2_port, 
      registers_29_1_port, registers_29_0_port, registers_30_31_port, 
      registers_30_30_port, registers_30_29_port, registers_30_28_port, 
      registers_30_27_port, registers_30_26_port, registers_30_25_port, 
      registers_30_24_port, registers_30_23_port, registers_30_22_port, 
      registers_30_21_port, registers_30_20_port, registers_30_19_port, 
      registers_30_18_port, registers_30_17_port, registers_30_16_port, 
      registers_30_15_port, registers_30_14_port, registers_30_13_port, 
      registers_30_12_port, registers_30_11_port, registers_30_10_port, 
      registers_30_9_port, registers_30_8_port, registers_30_7_port, 
      registers_30_6_port, registers_30_5_port, registers_30_4_port, 
      registers_30_3_port, registers_30_2_port, registers_30_1_port, 
      registers_30_0_port, registers_34_31_port, registers_34_30_port, 
      registers_34_29_port, registers_34_28_port, registers_34_27_port, 
      registers_34_26_port, registers_34_25_port, registers_34_24_port, 
      registers_34_23_port, registers_34_22_port, registers_34_21_port, 
      registers_34_20_port, registers_34_19_port, registers_34_18_port, 
      registers_34_17_port, registers_34_16_port, registers_34_15_port, 
      registers_34_14_port, registers_34_13_port, registers_34_12_port, 
      registers_34_11_port, registers_34_10_port, registers_34_9_port, 
      registers_34_8_port, registers_34_7_port, registers_34_6_port, 
      registers_34_5_port, registers_34_4_port, registers_34_3_port, 
      registers_34_2_port, registers_34_1_port, registers_34_0_port, 
      registers_36_31_port, registers_36_30_port, registers_36_29_port, 
      registers_36_28_port, registers_36_27_port, registers_36_26_port, 
      registers_36_25_port, registers_36_24_port, registers_36_23_port, 
      registers_36_22_port, registers_36_21_port, registers_36_20_port, 
      registers_36_19_port, registers_36_18_port, registers_36_17_port, 
      registers_36_16_port, registers_36_15_port, registers_36_14_port, 
      registers_36_13_port, registers_36_12_port, registers_36_11_port, 
      registers_36_10_port, registers_36_9_port, registers_36_8_port, 
      registers_36_7_port, registers_36_6_port, registers_36_5_port, 
      registers_36_4_port, registers_36_3_port, registers_36_2_port, 
      registers_36_1_port, registers_36_0_port, registers_37_31_port, 
      registers_37_30_port, registers_37_29_port, registers_37_28_port, 
      registers_37_27_port, registers_37_26_port, registers_37_25_port, 
      registers_37_24_port, registers_37_23_port, registers_37_22_port, 
      registers_37_21_port, registers_37_20_port, registers_37_19_port, 
      registers_37_18_port, registers_37_17_port, registers_37_16_port, 
      registers_37_15_port, registers_37_14_port, registers_37_13_port, 
      registers_37_12_port, registers_37_11_port, registers_37_10_port, 
      registers_37_9_port, registers_37_8_port, registers_37_7_port, 
      registers_37_6_port, registers_37_5_port, registers_37_4_port, 
      registers_37_3_port, registers_37_2_port, registers_37_1_port, 
      registers_37_0_port, registers_38_31_port, registers_38_30_port, 
      registers_38_29_port, registers_38_28_port, registers_38_27_port, 
      registers_38_26_port, registers_38_25_port, registers_38_24_port, 
      registers_38_23_port, registers_38_22_port, registers_38_21_port, 
      registers_38_20_port, registers_38_19_port, registers_38_18_port, 
      registers_38_17_port, registers_38_16_port, registers_38_15_port, 
      registers_38_14_port, registers_38_13_port, registers_38_12_port, 
      registers_38_11_port, registers_38_10_port, registers_38_9_port, 
      registers_38_8_port, registers_38_7_port, registers_38_6_port, 
      registers_38_5_port, registers_38_4_port, registers_38_3_port, 
      registers_38_2_port, registers_38_1_port, registers_38_0_port, 
      registers_40_31_port, registers_40_30_port, registers_40_29_port, 
      registers_40_28_port, registers_40_27_port, registers_40_26_port, 
      registers_40_25_port, registers_40_24_port, registers_40_23_port, 
      registers_40_22_port, registers_40_21_port, registers_40_20_port, 
      registers_40_19_port, registers_40_18_port, registers_40_17_port, 
      registers_40_16_port, registers_40_15_port, registers_40_14_port, 
      registers_40_13_port, registers_40_12_port, registers_40_11_port, 
      registers_40_10_port, registers_40_9_port, registers_40_8_port, 
      registers_40_7_port, registers_40_6_port, registers_40_5_port, 
      registers_40_4_port, registers_40_3_port, registers_40_2_port, 
      registers_40_1_port, registers_40_0_port, registers_41_31_port, 
      registers_41_30_port, registers_41_29_port, registers_41_28_port, 
      registers_41_27_port, registers_41_26_port, registers_41_25_port, 
      registers_41_24_port, registers_41_23_port, registers_41_22_port, 
      registers_41_21_port, registers_41_20_port, registers_41_19_port, 
      registers_41_18_port, registers_41_17_port, registers_41_16_port, 
      registers_41_15_port, registers_41_14_port, registers_41_13_port, 
      registers_41_12_port, registers_41_11_port, registers_41_10_port, 
      registers_41_9_port, registers_41_8_port, registers_41_7_port, 
      registers_41_6_port, registers_41_5_port, registers_41_4_port, 
      registers_41_3_port, registers_41_2_port, registers_41_1_port, 
      registers_41_0_port, registers_42_31_port, registers_42_30_port, 
      registers_42_29_port, registers_42_28_port, registers_42_27_port, 
      registers_42_26_port, registers_42_25_port, registers_42_24_port, 
      registers_42_23_port, registers_42_22_port, registers_42_21_port, 
      registers_42_20_port, registers_42_19_port, registers_42_18_port, 
      registers_42_17_port, registers_42_16_port, registers_42_15_port, 
      registers_42_14_port, registers_42_13_port, registers_42_12_port, 
      registers_42_11_port, registers_42_10_port, registers_42_9_port, 
      registers_42_8_port, registers_42_7_port, registers_42_6_port, 
      registers_42_5_port, registers_42_4_port, registers_42_3_port, 
      registers_42_2_port, registers_42_1_port, registers_42_0_port, 
      registers_43_31_port, registers_43_30_port, registers_43_29_port, 
      registers_43_28_port, registers_43_27_port, registers_43_26_port, 
      registers_43_25_port, registers_43_24_port, registers_43_23_port, 
      registers_43_22_port, registers_43_21_port, registers_43_20_port, 
      registers_43_19_port, registers_43_18_port, registers_43_17_port, 
      registers_43_16_port, registers_43_15_port, registers_43_14_port, 
      registers_43_13_port, registers_43_12_port, registers_43_11_port, 
      registers_43_10_port, registers_43_9_port, registers_43_8_port, 
      registers_43_7_port, registers_43_6_port, registers_43_5_port, 
      registers_43_4_port, registers_43_3_port, registers_43_2_port, 
      registers_43_1_port, registers_43_0_port, registers_44_31_port, 
      registers_44_30_port, registers_44_29_port, registers_44_28_port, 
      registers_44_27_port, registers_44_26_port, registers_44_25_port, 
      registers_44_24_port, registers_44_23_port, registers_44_22_port, 
      registers_44_21_port, registers_44_20_port, registers_44_19_port, 
      registers_44_18_port, registers_44_17_port, registers_44_16_port, 
      registers_44_15_port, registers_44_14_port, registers_44_13_port, 
      registers_44_12_port, registers_44_11_port, registers_44_10_port, 
      registers_44_9_port, registers_44_8_port, registers_44_7_port, 
      registers_44_6_port, registers_44_5_port, registers_44_4_port, 
      registers_44_3_port, registers_44_2_port, registers_44_1_port, 
      registers_44_0_port, registers_45_31_port, registers_45_30_port, 
      registers_45_29_port, registers_45_28_port, registers_45_27_port, 
      registers_45_26_port, registers_45_25_port, registers_45_24_port, 
      registers_45_23_port, registers_45_22_port, registers_45_21_port, 
      registers_45_20_port, registers_45_19_port, registers_45_18_port, 
      registers_45_17_port, registers_45_16_port, registers_45_15_port, 
      registers_45_14_port, registers_45_13_port, registers_45_12_port, 
      registers_45_11_port, registers_45_10_port, registers_45_9_port, 
      registers_45_8_port, registers_45_7_port, registers_45_6_port, 
      registers_45_5_port, registers_45_4_port, registers_45_3_port, 
      registers_45_2_port, registers_45_1_port, registers_45_0_port, 
      registers_47_31_port, registers_47_30_port, registers_47_29_port, 
      registers_47_28_port, registers_47_27_port, registers_47_26_port, 
      registers_47_25_port, registers_47_24_port, registers_47_23_port, 
      registers_47_22_port, registers_47_21_port, registers_47_20_port, 
      registers_47_19_port, registers_47_18_port, registers_47_17_port, 
      registers_47_16_port, registers_47_15_port, registers_47_14_port, 
      registers_47_13_port, registers_47_12_port, registers_47_11_port, 
      registers_47_10_port, registers_47_9_port, registers_47_8_port, 
      registers_47_7_port, registers_47_6_port, registers_47_5_port, 
      registers_47_4_port, registers_47_3_port, registers_47_2_port, 
      registers_47_1_port, registers_47_0_port, registers_48_31_port, 
      registers_48_30_port, registers_48_29_port, registers_48_28_port, 
      registers_48_27_port, registers_48_26_port, registers_48_25_port, 
      registers_48_24_port, registers_48_23_port, registers_48_22_port, 
      registers_48_21_port, registers_48_20_port, registers_48_19_port, 
      registers_48_18_port, registers_48_17_port, registers_48_16_port, 
      registers_48_15_port, registers_48_14_port, registers_48_13_port, 
      registers_48_12_port, registers_48_11_port, registers_48_10_port, 
      registers_48_9_port, registers_48_8_port, registers_48_7_port, 
      registers_48_6_port, registers_48_5_port, registers_48_4_port, 
      registers_48_3_port, registers_48_2_port, registers_48_1_port, 
      registers_48_0_port, registers_49_31_port, registers_49_30_port, 
      registers_49_29_port, registers_49_28_port, registers_49_27_port, 
      registers_49_26_port, registers_49_25_port, registers_49_24_port, 
      registers_49_23_port, registers_49_22_port, registers_49_21_port, 
      registers_49_20_port, registers_49_19_port, registers_49_18_port, 
      registers_49_17_port, registers_49_16_port, registers_49_15_port, 
      registers_49_14_port, registers_49_13_port, registers_49_12_port, 
      registers_49_11_port, registers_49_10_port, registers_49_9_port, 
      registers_49_8_port, registers_49_7_port, registers_49_6_port, 
      registers_49_5_port, registers_49_4_port, registers_49_3_port, 
      registers_49_2_port, registers_49_1_port, registers_49_0_port, 
      registers_50_31_port, registers_50_30_port, registers_50_29_port, 
      registers_50_28_port, registers_50_27_port, registers_50_26_port, 
      registers_50_25_port, registers_50_24_port, registers_50_23_port, 
      registers_50_22_port, registers_50_21_port, registers_50_20_port, 
      registers_50_19_port, registers_50_18_port, registers_50_17_port, 
      registers_50_16_port, registers_50_15_port, registers_50_14_port, 
      registers_50_13_port, registers_50_12_port, registers_50_11_port, 
      registers_50_10_port, registers_50_9_port, registers_50_8_port, 
      registers_50_7_port, registers_50_6_port, registers_50_5_port, 
      registers_50_4_port, registers_50_3_port, registers_50_2_port, 
      registers_50_1_port, registers_50_0_port, registers_51_31_port, 
      registers_51_30_port, registers_51_29_port, registers_51_28_port, 
      registers_51_27_port, registers_51_26_port, registers_51_25_port, 
      registers_51_24_port, registers_51_23_port, registers_51_22_port, 
      registers_51_21_port, registers_51_20_port, registers_51_19_port, 
      registers_51_18_port, registers_51_17_port, registers_51_16_port, 
      registers_51_15_port, registers_51_14_port, registers_51_13_port, 
      registers_51_12_port, registers_51_11_port, registers_51_10_port, 
      registers_51_9_port, registers_51_8_port, registers_51_7_port, 
      registers_51_6_port, registers_51_5_port, registers_51_4_port, 
      registers_51_3_port, registers_51_2_port, registers_51_1_port, 
      registers_51_0_port, registers_54_31_port, registers_54_30_port, 
      registers_54_29_port, registers_54_28_port, registers_54_27_port, 
      registers_54_26_port, registers_54_25_port, registers_54_24_port, 
      registers_54_23_port, registers_54_22_port, registers_54_21_port, 
      registers_54_20_port, registers_54_19_port, registers_54_18_port, 
      registers_54_17_port, registers_54_16_port, registers_54_15_port, 
      registers_54_14_port, registers_54_13_port, registers_54_12_port, 
      registers_54_11_port, registers_54_10_port, registers_54_9_port, 
      registers_54_8_port, registers_54_7_port, registers_54_6_port, 
      registers_54_5_port, registers_54_4_port, registers_54_3_port, 
      registers_54_2_port, registers_54_1_port, registers_54_0_port, 
      registers_55_31_port, registers_55_30_port, registers_55_29_port, 
      registers_55_28_port, registers_55_27_port, registers_55_26_port, 
      registers_55_25_port, registers_55_24_port, registers_55_23_port, 
      registers_55_22_port, registers_55_21_port, registers_55_20_port, 
      registers_55_19_port, registers_55_18_port, registers_55_17_port, 
      registers_55_16_port, registers_55_15_port, registers_55_14_port, 
      registers_55_13_port, registers_55_12_port, registers_55_11_port, 
      registers_55_10_port, registers_55_9_port, registers_55_8_port, 
      registers_55_7_port, registers_55_6_port, registers_55_5_port, 
      registers_55_4_port, registers_55_3_port, registers_55_2_port, 
      registers_55_1_port, registers_55_0_port, registers_56_31_port, 
      registers_56_30_port, registers_56_29_port, registers_56_28_port, 
      registers_56_27_port, registers_56_26_port, registers_56_25_port, 
      registers_56_24_port, registers_56_23_port, registers_56_22_port, 
      registers_56_21_port, registers_56_20_port, registers_56_19_port, 
      registers_56_18_port, registers_56_17_port, registers_56_16_port, 
      registers_56_15_port, registers_56_14_port, registers_56_13_port, 
      registers_56_12_port, registers_56_11_port, registers_56_10_port, 
      registers_56_9_port, registers_56_8_port, registers_56_7_port, 
      registers_56_6_port, registers_56_5_port, registers_56_4_port, 
      registers_56_3_port, registers_56_2_port, registers_56_1_port, 
      registers_56_0_port, registers_59_31_port, registers_59_30_port, 
      registers_59_29_port, registers_59_28_port, registers_59_27_port, 
      registers_59_26_port, registers_59_25_port, registers_59_24_port, 
      registers_59_23_port, registers_59_22_port, registers_59_21_port, 
      registers_59_20_port, registers_59_19_port, registers_59_18_port, 
      registers_59_17_port, registers_59_16_port, registers_59_15_port, 
      registers_59_14_port, registers_59_13_port, registers_59_12_port, 
      registers_59_11_port, registers_59_10_port, registers_59_9_port, 
      registers_59_8_port, registers_59_7_port, registers_59_6_port, 
      registers_59_5_port, registers_59_4_port, registers_59_3_port, 
      registers_59_2_port, registers_59_1_port, registers_59_0_port, 
      registers_60_31_port, registers_60_30_port, registers_60_29_port, 
      registers_60_28_port, registers_60_27_port, registers_60_26_port, 
      registers_60_25_port, registers_60_24_port, registers_60_23_port, 
      registers_60_22_port, registers_60_21_port, registers_60_20_port, 
      registers_60_19_port, registers_60_18_port, registers_60_17_port, 
      registers_60_16_port, registers_60_15_port, registers_60_14_port, 
      registers_60_13_port, registers_60_12_port, registers_60_11_port, 
      registers_60_10_port, registers_60_9_port, registers_60_8_port, 
      registers_60_7_port, registers_60_6_port, registers_60_5_port, 
      registers_60_4_port, registers_60_3_port, registers_60_2_port, 
      registers_60_1_port, registers_60_0_port, registers_62_31_port, 
      registers_62_30_port, registers_62_29_port, registers_62_28_port, 
      registers_62_27_port, registers_62_26_port, registers_62_25_port, 
      registers_62_24_port, registers_62_23_port, registers_62_22_port, 
      registers_62_21_port, registers_62_20_port, registers_62_19_port, 
      registers_62_18_port, registers_62_17_port, registers_62_16_port, 
      registers_62_15_port, registers_62_14_port, registers_62_13_port, 
      registers_62_12_port, registers_62_11_port, registers_62_10_port, 
      registers_62_9_port, registers_62_8_port, registers_62_7_port, 
      registers_62_6_port, registers_62_5_port, registers_62_4_port, 
      registers_62_3_port, registers_62_2_port, registers_62_1_port, 
      registers_62_0_port, registers_63_31_port, registers_63_30_port, 
      registers_63_29_port, registers_63_28_port, registers_63_27_port, 
      registers_63_26_port, registers_63_25_port, registers_63_24_port, 
      registers_63_23_port, registers_63_22_port, registers_63_21_port, 
      registers_63_20_port, registers_63_19_port, registers_63_18_port, 
      registers_63_17_port, registers_63_16_port, registers_63_15_port, 
      registers_63_14_port, registers_63_13_port, registers_63_12_port, 
      registers_63_11_port, registers_63_10_port, registers_63_9_port, 
      registers_63_8_port, registers_63_7_port, registers_63_6_port, 
      registers_63_5_port, registers_63_4_port, registers_63_3_port, 
      registers_63_2_port, registers_63_1_port, registers_63_0_port, 
      registers_68_31_port, registers_68_30_port, registers_68_29_port, 
      registers_68_28_port, registers_68_27_port, registers_68_26_port, 
      registers_68_25_port, registers_68_24_port, registers_68_23_port, 
      registers_68_22_port, registers_68_21_port, registers_68_20_port, 
      registers_68_19_port, registers_68_18_port, registers_68_17_port, 
      registers_68_16_port, registers_68_15_port, registers_68_14_port, 
      registers_68_13_port, registers_68_12_port, registers_68_11_port, 
      registers_68_10_port, registers_68_9_port, registers_68_8_port, 
      registers_68_7_port, registers_68_6_port, registers_68_5_port, 
      registers_68_4_port, registers_68_3_port, registers_68_2_port, 
      registers_68_1_port, registers_68_0_port, swp_5_port, swp_4_port, 
      swp_3_port, swp_2_port, swp_1_port, swp_0_port, lastcwp_4_port, 
      lastcwp_3_port, lastcwp_2_port, lastcwp_1_port, N273, N274, N275, N276, 
      N9641, i_5_port, i_4_port, i_3_port, i_2_port, i_1_port, i_0_port, N9908,
      N9909, N9910, N9921, N9922, N9923, N9924, N9925, N9926, N45784, N45785, 
      N45786, N45787, N45788, N45789, N46298, N46299, N46300, N46301, N46302, 
      N46303, N51637, n7587, n7588, n7589, n7590, n7591, n7592, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
      n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, 
      n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, 
      n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
      n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
      n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
      n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
      n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
      n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
      n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641_port, n9642, n9643
      , n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
      n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
      n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, 
      n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, 
      n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, 
      n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
      n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
      n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, 
      n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, 
      n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
      n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, 
      n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, 
      n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, 
      n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
      n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, 
      n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, 
      n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, 
      n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, 
      n9904, n9905, n9906, n9907, n9908_port, n9909_port, n9910_port, n9911, 
      n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921_port
      , n9922_port, n9923_port, n9924_port, n9925_port, n9926_port, n9927, 
      n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, 
      n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, 
      n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, 
      n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
      n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, 
      n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, 
      n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, 
      n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
      n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, 
      n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, 
      n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, 
      n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, 
      n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, 
      n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, 
      n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
      n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, 
      n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, 
      n10124, n10125, n10127, n10128, n10129, n10130, n10131, n10132, n10133, 
      n10134, n10135, n10136, n10137, n10138, n10140, n10141, n10142, n10143, 
      n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, 
      n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, 
      n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, 
      n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, 
      n10180, n10181, n10182, n10183, n10184, n10185, n10187, n10188, n10189, 
      n10190, add_73_carry_1_port, add_73_carry_2_port, add_73_carry_3_port, 
      add_73_carry_4_port, add_73_carry_5_port, r590_carry_5_port, n3043, n5522
      , n6613, n6620, n6621, n6624, n6630, n6632, n6634, n6641, n6642, n6646, 
      n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, 
      n6657, n6658, n6659, n6660, n6671, n6674, n6676, n6683, n6684, n6687, 
      n6693, n6695, net226799, net226800, net226801, net226802, net226803, 
      net226804, net226805, net226806, net226807, net226808, net226809, 
      net226810, net226811, net226812, net226813, net226814, net226815, 
      net226816, net226817, net226818, net226819, net226820, net226821, 
      net226822, net226823, net226824, net226825, net226826, net226827, 
      net226828, net226829, net226830, net226831, net226832, net226833, 
      net226834, net226835, net226836, net226837, net226838, net226839, 
      net226840, net226841, net226842, net226843, net226844, net226845, 
      net226846, net226847, net226848, net226849, net226850, net226851, 
      net226852, net226853, net226854, net226855, net226856, net226857, 
      net226858, net226859, net226860, net226861, net226862, net226863, 
      net226864, net226865, net226866, net226867, net226868, net226869, 
      net226870, net226871, net226872, net226873, net226874, net226875, 
      net226876, net226877, net226878, net226879, net226880, net226881, 
      net226882, net226883, net226884, net226885, net226886, net226887, 
      net226888, net226889, net226890, net226891, net226892, net226893, 
      net226894, net226895, net226896, net226897, net226898, net226899, 
      net226900, net226901, net226902, net226903, net226904, net226905, 
      net226906, net226907, net226908, net226909, net226910, net226911, 
      net226912, net226913, net226914, net226915, net226916, net226917, 
      net226918, net226919, net226920, net226921, net226922, net226923, 
      net226924, net226925, net226926, net226927, net226928, net226929, 
      net226930, net226931, net226932, net226933, net226934, net226935, 
      net226936, net226937, net226938, net226939, net226940, net226941, 
      net226942, net226943, net226944, net226945, net226946, net226947, 
      net226948, net226949, net226950, net226951, net226952, net226953, 
      net226954, net226955, net226956, net226957, net226958, net226959, 
      net226960, net226961, net226962, net226963, net226964, net226965, 
      net226966, net226967, net226968, net226969, net226970, net226971, 
      net226972, net226973, net226974, net226975, net226976, net226977, 
      net226978, net226979, net226980, net226981, net226982, net226983, 
      net226984, net226985, net226986, net226987, net226988, net226989, 
      net226990, net226991, net226992, net226993, net226994, net226995, 
      net226996, net226997, net226998, net226999, net227000, net227001, 
      net227002, net227003, net227004, net227005, net227006, net227007, 
      net227008, net227009, net227010, net227011, net227012, net227013, 
      net227014, net227015, net227016, net227017, net227018, net227019, 
      net227020, net227021, net227022, net227023, net227024, net227025, 
      net227026, net227027, net227028, net227029, net227030, net227031, 
      net227032, net227033, net227034, net227035, net227036, net227037, 
      net227038, net227039, net227040, net227041, net227042, net227043, 
      net227044, net227045, net227046, net227047, net227048, net227049, 
      net227050, net227051, net227052, net227053, net227054, net227055, 
      net227056, net227057, net227058, net227059, net227060, net227061, 
      net227062, net227063, net227064, net227065, net227066, net227067, 
      net227068, net227069, net227070, net227071, net227072, net227073, 
      net227074, net227075, net227076, net227077, net227078, net227079, 
      net227080, net227081, net227082, net227083, net227084, net227085, 
      net227086, net227087, net227088, net227089, net227090, net227091, 
      net227092, net227093, net227094, net227095, net227096, net227097, 
      net227098, net227099, net227100, net227101, net227102, net227103, 
      net227104, net227105, net227106, net227107, net227108, net227109, 
      net227110, net227111, net227112, net227113, net227114, net227115, 
      net227116, net227117, net227118, net227119, net227120, net227121, 
      net227122, net227123, net227124, net227125, net227126, net227127, 
      net227128, net227129, net227130, net227131, net227132, net227133, 
      net227134, net227135, net227136, net227137, net227138, net227139, 
      net227140, net227141, net227142, net227143, net227144, net227145, 
      net227146, net227147, net227148, net227149, net227150, net227151, 
      net227152, net227153, net227154, net227155, net227156, net227157, 
      net227158, net227159, net227160, net227161, net227162, net227163, 
      net227164, net227165, net227166, net227167, net227168, net227169, 
      net227170, net227171, net227172, net227173, net227174, net227175, 
      net227176, net227177, net227178, net227179, net227180, net227181, 
      net227182, net227183, net227184, net227185, net227186, net227187, 
      net227188, net227189, net227190, net227191, net227192, net227193, 
      net227194, net227195, net227196, net227197, net227198, net227199, 
      net227200, net227201, net227202, net227203, net227204, net227205, 
      net227206, net227207, net227208, net227209, net227210, net227211, 
      net227212, net227213, net227214, net227215, net227216, net227217, 
      net227218, net227219, net227220, net227221, net227222, net227223, 
      net227224, net227225, net227226, net227227, net227228, net227229, 
      net227230, net227231, net227232, net227233, net227234, net227235, 
      net227236, net227237, net227238, net227239, net227240, net227241, 
      net227242, net227243, net227244, net227245, net227246, net227247, 
      net227248, net227249, net227250, net227251, net227252, net227253, 
      net227254, net227255, net227256, net227257, net227258, net227259, 
      net227260, net227261, net227262, net227263, net227264, net227265, 
      net227266, net227267, net227268, net227269, net227270, net227271, 
      net227272, net227273, net227274, net227275, net227276, net227277, 
      net227278, net227279, net227280, net227281, net227282, net227283, 
      net227284, net227285, net227286, net227287, net227288, net227289, 
      net227290, net227291, net227292, net227293, net227294, net227295, 
      net227296, net227297, net227298, net227299, net227300, net227301, 
      net227302, net227303, net227304, net227305, net227306, net227307, 
      net227308, net227309, net227310, net227311, net227312, net227313, 
      net227314, net227315, net227316, net227317, net227318, net227319, 
      net227320, net227321, net227322, net227323, net227324, net227325, 
      net227326, net227327, net227328, net227329, net227330, net227331, 
      net227332, net227333, net227334, net227335, net227336, net227337, 
      net227338, net227339, net227340, net227341, net227342, net227343, 
      net227344, net227345, net227346, net227347, net227348, net227349, 
      net227350, net227351, net227352, net227353, net227354, net227355, 
      net227356, net227357, net227358, net227359, net227360, net227361, 
      net227362, net227363, net227364, net227365, net227366, net227367, 
      net227368, net227369, net227370, net227371, net227372, net227373, 
      net227374, net227375, net227376, net227377, net227378, net227379, 
      net227380, net227381, net227382, net227383, net227384, net227385, 
      net227386, net227387, net227388, net227389, net227390, net227391, 
      net227392, net227393, net227394, net227395, net227396, net227397, 
      net227398, net227399, net227400, net227401, net227402, net227403, 
      net227404, net227405, net227406, net227407, net227408, net227409, 
      net227410, net227411, net227412, net227413, net227414, net227415, 
      net227416, net227417, net227418, net227419, net227420, net227421, 
      net227422, net227423, net227424, net227425, net227426, net227427, 
      net227428, net227429, net227430, net227431, net227432, net227433, 
      net227434, net227435, net227436, net227437, net227438, net227439, 
      net227440, net227441, net227442, net227443, net227444, net227445, 
      net227446, net227447, net227448, net227449, net227450, net227451, 
      net227452, net227453, net227454, net227455, net227456, net227457, 
      net227458, net227459, net227460, net227461, net227462, net227463, 
      net227464, net227465, net227466, net227467, net227468, net227469, 
      net227470, net227471, net227472, net227473, net227474, net227475, 
      net227476, net226798, net226797, n4, n76, n77, n4058, n4059, n4062, n4067
      , n4070, n4073, n4076, n4079, n4082, n4085, n4088, n4090, n4091, n4095, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4106, n4107, n4108, n4109, 
      n4110, n4112, n4114, n4117, n4118, n4119, n4121, n4123, n4124, n4125, 
      n4126, n4128, n4130, n4131, n4132, n4133, n4135, n4137, n4138, n4139, 
      n4140, n4141, n4142, n4145, n4148, n4150, n4152, n4153, n4156, n4157, 
      n4159, n4161, n4162, n4163, n4164, n4168, n4170, n4171, n4172, n4173, 
      n4175, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4186, 
      n4188, n4189, n4190, n4191, n4192, n4195, n4198, n4199, n4200, n4202, 
      n4206, n4207, n4208, n4209, n4211, n4213, n4214, n4217, n4218, n4219, 
      n4220, n4221, n4222, n4223, n4225, n4226, n4227, n4228, n4230, n4232, 
      n4233, n4234, n4235, n4237, n4239, n4240, n4241, n4242, n4248, n4251, 
      n4256, n4259, n4262, n4267, n4270, n4273, n4275, n4278, n4279, n4282, 
      n4285, n4288, n4291, n4298, n4301, n4306, n4309, n4312, n4317, n4320, 
      n4323, n4326, n4329, n4332, n4335, n4338, n4341, n4348, n4351, n4356, 
      n4359, n4362, n4367, n4370, n4373, n4376, n4379, n4382, n4385, n4388, 
      n4391, n4398, n4401, n4406, n4409, n4412, n4417, n4420, n4423, n4426, 
      n4429, n4432, n4435, n4438, n4441, n4448, n4451, n4456, n4459, n4462, 
      n4467, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4495, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
      n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4533, n4611, 
      n4612, n4613, n4614, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4645, 
      n4648, n4649, n4650, n4651, n4652, n4653, n4664, n4738, n4739, n4740, 
      n4741, n4742, n4745, n4748, n4749, n4750, n4751, n4752, n4753, n4756, 
      n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4767, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4791, n4871, n4872, n4873, n4874, n4875, 
      n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, 
      n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4895, n4898, n4899, 
      n4900, n4901, n4902, n4903, n4906, n4907, n4908, n4909, n4910, n4911, 
      n4912, n4913, n4924, n4993, n4994, n4995, n4996, n4997, n4998, n4999, 
      n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, 
      n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5020, n5021, 
      n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, 
      n5040, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5146, n5147, n5157, n5257, 
      n5259, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5285, n5286, n5288, n5290, n5291, n5292, n5293, n5294, n5295, 
      n5298, n5299, n5301, n5302, n5303, n5304, n5305, n5307, n5309, n5311, 
      n5312, n5313, n5314, n5315, n5316, n5319, n5343, n5442, n5443, n5446, 
      n5447, n5448, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
      n5472, n5473, n5475, n5476, n5478, n5480, n5481, n5482, n5483, n5484, 
      n5485, n5488, n5489, n5491, n5492, n5493, n5494, n5495, n5497, n5499, 
      n5501, n5502, n5503, n5504, n5530, n5629, n5630, n5631, n5632, n5635, 
      n5636, n5637, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, 
      n5661, n5662, n5664, n5665, n5667, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5677, n5678, n5680, n5681, n5682, n5683, n5684, n5686, n5688, 
      n5690, n5691, n5717, n5816, n5817, n5818, n5819, n5820, n5821, n5824, 
      n5825, n5826, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, 
      n5850, n5851, n5853, n5854, n5856, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5866, n5867, n5869, n5870, n5871, n5872, n5873, n5875, n5877, 
      n5889, n6001, n6003, n6005, n6006, n6007, n6008, n6009, n6010, n6013, 
      n6014, n6015, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, 
      n6039, n6040, n6042, n6043, n6045, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6055, n6056, n6058, n6059, n6060, n6061, n6062, n6076, n6187, 
      n6188, n6190, n6192, n6194, n6195, n6196, n6197, n6198, n6199, n6202, 
      n6203, n6204, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6231, n6232, n6234, n6236, n6237, n6238, n6239, n6240, 
      n6241, n6244, n6245, n6247, n6248, n6249, n6261, n6374, n6375, n6376, 
      n6377, n6379, n6381, n6383, n6384, n6385, n6386, n6387, n6388, n6391, 
      n6392, n6393, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, 
      n6417, n6418, n6420, n6421, n6423, n6425, n6426, n6427, n6428, n6429, 
      n6430, n6433, n6434, n6436, n6448, n6560, n6562, n6563, n6564, n6565, 
      n6566, n6568, n6570, n6572, n6573, n6574, n6575, n6576, n6577, n6580, 
      n6581, n6582, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
      n6606, n6607, n6609, n6610, n6612, n6614, n6615, n6616, n6617, n6618, 
      n6619, n6622, n6635, n6724, n6725, n6726, n6727, n6728, n6729, n6730, 
      n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, 
      n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, 
      n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, 
      n6769, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6878, n6942, 
      n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, 
      n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, 
      n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
      n6973, n6974, n6975, n6976, n6977, n6978, n6987, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7096, n7160, n7161, n7162, n7163, n7164, 
      n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, 
      n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, 
      n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, 
      n7195, n7196, n7205, n7274, n7275, n7276, n7277, n7278, n7279, n7280, 
      n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, 
      n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, 
      n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, 
      n7319, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7428, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, 
      n7523, n7524, n7525, n7526, n7527, n7528, n7537, n7607, n7608, n7609, 
      n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, 
      n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, 
      n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, 
      n7640, n7641, n7642, n7643, n7652, n10243, n10244, n10245, n10246, n10247
      , n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
      n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, 
      n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, 
      n10275, n10276, n10277, n10278, n10279, n10280, n10282, n10283, n10285, 
      n10286, n10287, n10288, n10290, n10292, n10300, n10303, n10306, n10315, 
      n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, 
      n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, 
      n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, 
      n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10400, n10405, n10410, n10413, n10416, n10425, n10444, n10448, 
      n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, 
      n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, 
      n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, 
      n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, 
      n10501, n10510, n10511, n10513, n10514, n10515, n10516, n10517, n10518, 
      n10519, n10520, n10522, n10523, n10524, n10525, n10526, n10527, n10528, 
      n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, 
      n10538, n10540, n10542, n10543, n10544, n10545, n10547, n10549, n10550, 
      n10551, n10552, n10554, n10556, n10557, n10558, n10560, n10562, n10563, 
      n10564, n10565, n10566, n10567, n10568, n10569, n10571, n10573, n10575, 
      n10576, n10577, n10578, n10580, n10582, n10583, n10584, n10585, n10587, 
      n10589, n10590, n10591, n10592, n10594, n10596, n10597, n10598, n10599, 
      n10600, n10601, n10602, n10603, n10605, n10607, n10608, n10609, n10610, 
      n10612, n10614, n10615, n10616, n10617, n10619, n10621, n10622, n10623, 
      n10624, n10626, n10628, n10629, n10630, n10631, n10632, n10633, n10634, 
      n10635, n10637, n10639, n10641, n10642, n10643, n10644, n10646, n10648, 
      n10649, n10650, n10651, n10653, n10655, n10656, n10657, n10658, n10660, 
      n10662, n10663, n10665, n10666, n10667, n10668, n10669, n10670, n10671, 
      n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10682, 
      n10683, n10685, n10687, n10688, n10689, n10690, n10691, n10694, n10695, 
      n10698, n10700, n10701, n10702, n10703, n10704, n10707, n10709, n10711, 
      n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10724, 
      n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, 
      n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, 
      n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, 
      n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, 
      n10761, n10762, n10763, n10764, n10765, n10767, n10768, n10769, n10770, 
      n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, 
      n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, 
      n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, 
      n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, 
      n10807, n10808, n10810, n10811, n10812, n10813, n10814, n10815, n10816, 
      n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, 
      n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, 
      n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, 
      n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10853, 
      n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, 
      n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, 
      n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, 
      n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, 
      n10890, n10891, n10892, n10893, n10894, n10896, n10897, n10898, n10899, 
      n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, 
      n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, 
      n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, 
      n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, 
      n10936, n10937, n10939, n10940, n10941, n10942, n10943, n10944, n10945, 
      n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, 
      n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, 
      n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, 
      n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11025, n11026, n11027, n11028, 
      n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, 
      n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, 
      n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, 
      n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, 
      n11065, n11066, n11068, n11069, n11070, n11071, n11072, n11073, n11074, 
      n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, 
      n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, 
      n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, 
      n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11111, 
      n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, 
      n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, 
      n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, 
      n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, 
      n11148, n11149, n11150, n11151, n11152, n11154, n11155, n11156, n11157, 
      n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, 
      n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, 
      n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, 
      n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, 
      n11194, n11195, n11197, n11198, n11199, n11200, n11201, n11202, n11203, 
      n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, 
      n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, 
      n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, 
      n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11240, 
      n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
      n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, 
      n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, 
      n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, 
      n11277, n11278, n11279, n11280, n11281, n11283, n11284, n11285, n11286, 
      n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, 
      n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, 
      n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, 
      n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, 
      n11323, n11324, n11326, n11327, n11328, n11329, n11330, n11331, n11332, 
      n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, 
      n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, 
      n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, 
      n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11369, 
      n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, 
      n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, 
      n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, 
      n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, 
      n11406, n11407, n11408, n11409, n11410, n11412, n11413, n11414, n11415, 
      n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, 
      n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, 
      n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, 
      n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, 
      n11452, n11453, n11455, n11456, n11457, n11458, n11459, n11460, n11462, 
      n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, 
      n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, 
      n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, 
      n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11499, 
      n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, 
      n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, 
      n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, 
      n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, 
      n11536, n11537, n11538, n11539, n11540, n11542, n11543, n11544, n11545, 
      n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, 
      n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
      n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, 
      n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, 
      n11582, n11583, n11585, n11586, n11587, n11588, n11589, n11590, n11591, 
      n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, 
      n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, 
      n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, 
      n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11628, 
      n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, 
      n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, 
      n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, 
      n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, 
      n11665, n11666, n11667, n11668, n11669, n11671, n11672, n11673, n11674, 
      n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, 
      n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, 
      n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, 
      n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, 
      n11711, n11712, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, 
      n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11757, 
      n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, 
      n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, 
      n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, 
      n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, 
      n11794, n11795, n11796, n11797, n11798, n11800, n11801, n11802, n11803, 
      n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, 
      n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, 
      n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, 
      n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, 
      n11840, n11841, n11843, n11848, n11853, n11859, n11868, n11908, n11909, 
      n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, 
      n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, 
      n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, 
      n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11953, 
      n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, 
      n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, 
      n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, 
      n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, 
      n11990, n11991, n11992, n11993, n11994, n11996, n12029, n12061, n12062, 
      n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, 
      n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, 
      n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, 
      n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12106, 
      n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, 
      n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, 
      n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, 
      n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, 
      n12143, n12144, n12145, n12146, n12147, n12149, n12184, n12216, n12217, 
      n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, 
      n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, 
      n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, 
      n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12259, 
      n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, 
      n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, 
      n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, 
      n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, 
      n12296, n12297, n12298, n12299, n12300, n12302, n12338, n12370, n12371, 
      n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, 
      n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, 
      n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, 
      n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12412, 
      n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, 
      n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, 
      n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, 
      n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, 
      n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, 
      n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, 
      n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, 
      n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, 
      n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, 
      n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, 
      n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, 
      n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, 
      n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, 
      n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, 
      n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, 
      n12548, n12549, n12550, n12552, n12553, n12554, n12555, n12556, n12557, 
      n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, 
      n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, 
      n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, 
      n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, 
      n12594, n12595, n12596, n12597, n12598, n12599, n12601, n12603, n12604, 
      n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, 
      n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, 
      n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, 
      n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, 
      n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, 
      n12650, n12651, n12653, n12654, n12655, n12656, n12657, n12658, n12659, 
      n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, 
      n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, 
      n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, 
      n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, 
      n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, 
      n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, 
      n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, 
      n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, 
      n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, 
      n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, 
      n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, 
      n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, 
      n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, 
      n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, 
      n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, 
      n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, 
      n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, 
      n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, 
      n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, 
      n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, 
      n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, 
      n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, 
      n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, 
      n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, 
      n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, 
      n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, 
      n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, 
      n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, 
      n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, 
      n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, 
      n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, 
      n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, 
      n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, 
      n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, 
      n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, 
      n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, 
      n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, 
      n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, 
      n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, 
      n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, 
      n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, 
      n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, 
      n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, 
      n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, 
      n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, 
      n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, 
      n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, 
      n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, 
      n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, 
      n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, 
      n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, 
      n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, 
      n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, 
      n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, 
      n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, 
      n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, 
      n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, 
      n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, 
      n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, 
      n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, 
      n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, 
      n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, 
      n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, 
      n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, 
      n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, 
      n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, 
      n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, 
      n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, 
      n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, 
      n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, 
      n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, 
      n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, 
      n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, 
      n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, 
      n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, 
      n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, 
      n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, 
      n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, 
      n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, 
      n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, 
      n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, 
      n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, 
      n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, 
      n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, 
      n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, 
      n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, 
      n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, 
      n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, 
      n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, 
      n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, 
      n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, 
      n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, 
      n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, 
      n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, 
      n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, 
      n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, 
      n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, 
      n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, 
      n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, 
      n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, 
      n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, 
      n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, 
      n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, 
      n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, 
      n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, 
      n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, 
      n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, 
      n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, 
      n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, 
      n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, 
      n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, 
      n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, 
      n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, 
      n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, 
      n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, 
      n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, 
      n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, 
      n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, 
      n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, 
      n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, 
      n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
      n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, 
      n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, 
      n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, 
      n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, 
      n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, 
      n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, 
      n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, 
      n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, 
      n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, 
      n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, 
      n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, 
      n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, 
      n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, 
      n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, 
      n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, 
      n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, 
      n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, 
      n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, 
      n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, 
      n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, 
      n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, 
      n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, 
      n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, 
      n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, 
      n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, 
      n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, 
      n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, 
      n13993, n13994, n13995, n13997, n13998, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14009, n14010, n14011, n14012, n14013, 
      n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, 
      n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14033, n14034, 
      n14058, n14059, n14061, n14062, n14063, n14064, n14066, n14067, n14068, 
      n14070, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, 
      n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, 
      n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, 
      n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, 
      n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, 
      n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, 
      n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, 
      n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, 
      n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, 
      n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, 
      n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, 
      n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, 
      n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, 
      n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, 
      n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, 
      n14206, n14207, n14208, n14209, n14210, n14211, n14213, n14214, n14215, 
      n14217, n14218, n14220, n14221, n14222, n14223, n14224, n14226, n14228, 
      n14229, n14231, n14232, n14233, n14234, n14236, n14237, n14238, n14239, 
      n14240, n14241, n14244, n14245, n14247, n14248, n14249, n14250, n14251, 
      n14252, n14253, n14254, n14256, n14257, n14258, n14259, n14260, n14262, 
      n14263, n14265, n14266, n14267, n11498, n11541, n11584, n11627, n11670, 
      n11713, n11756, n11799, n11842, n11844, n11845, n11846, n11847, n11849, 
      n11850, n11851, n11852, n11854, n11855, n11856, n11857, n11858, n11860, 
      n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11869, n11870, 
      n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, 
      n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, 
      n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, 
      n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, 
      n11907, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, 
      n11995, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, 
      n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, 
      n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, 
      n12023, n12024, n12025, n12026, n12027, n12028, n12030, n12031, n12032, 
      n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, 
      n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, 
      n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, 
      n12060, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, 
      n12148, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, 
      n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, 
      n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, 
      n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12185, 
      n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, 
      n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, 
      n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, 
      n12213, n12214, n12215, n12253, n12254, n12255, n12256, n12257, n12258, 
      n12301, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, 
      n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, 
      n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, 
      n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, 
      n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, 
      n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, 
      n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, 
      n12366, n12367, n12368, n12369, n12407, n12408, n12409, n12410, n12411, 
      n12551, n12600, n12602, n12652, n12669, n13996, n13999, n14008, n14014, 
      n14015, n14032, n14035, n14036, n14037, n14038, n14039, n14040, n14041, 
      n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, 
      n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14060, n14065, 
      n14069, n14071, n14212, n14216, n14219, n14225, n14227, n14230, n14235, 
      n14242, n14243, n14246, n14255, n14261, n14264, n14268, n14269, n14270, 
      n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, 
      n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, 
      n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, 
      n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, 
      n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, 
      n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, 
      n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, 
      n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, 
      n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, 
      n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, 
      n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, 
      n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, 
      n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, 
      n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, 
      n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, 
      n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, 
      n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, 
      n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, 
      n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, 
      n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, 
      n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, 
      n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, 
      n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, 
      n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, 
      n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, 
      n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, 
      n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, 
      n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, 
      n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, 
      n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, 
      n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, 
      n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, 
      n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, 
      n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, 
      n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, 
      n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, 
      n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, 
      n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, 
      n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, 
      n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, 
      n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, 
      n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, 
      n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, 
      n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, 
      n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, 
      n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, 
      n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, 
      n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, 
      n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, 
      n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, 
      n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, 
      n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, 
      n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, 
      n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, 
      n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, 
      n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, 
      n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, 
      n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, 
      n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, 
      n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, 
      n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, 
      n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, 
      n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, 
      n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, 
      n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, 
      n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, 
      n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, 
      n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, 
      n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, 
      n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, 
      n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, 
      n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, 
      n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, 
      n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, 
      n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, 
      n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, 
      n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, 
      n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, 
      n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, 
      n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, 
      n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, 
      n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, 
      n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, 
      n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, 
      n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, 
      n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, 
      n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, 
      n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, 
      n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, 
      n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, 
      n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, 
      n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, 
      n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
      n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, 
      n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, 
      n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, 
      n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, 
      n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, 
      n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, 
      n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, 
      n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, 
      n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, 
      n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, 
      n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, 
      n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, 
      n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, 
      n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, 
      n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, 
      n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, 
      n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, 
      n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, 
      n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, 
      n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, 
      n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, 
      n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, 
      n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, 
      n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, 
      n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, 
      n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, 
      n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, 
      n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, 
      n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, 
      n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, 
      n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, 
      n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, 
      n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, 
      n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, 
      n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, 
      n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, 
      n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, 
      n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, 
      n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, 
      n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, 
      n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, 
      n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, 
      n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, 
      n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, 
      n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, 
      n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, 
      n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, 
      n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, 
      n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, 
      n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, 
      n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, 
      n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, 
      n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, 
      n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, 
      n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, 
      n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, 
      n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, 
      n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, 
      n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, 
      n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, 
      n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, 
      n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, 
      n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, 
      n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, 
      n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, 
      n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, 
      n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, 
      n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, 
      n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, 
      n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, 
      n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, 
      n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, 
      n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, 
      n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, 
      n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, 
      n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, 
      n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, 
      n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, 
      n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, 
      n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, 
      n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, 
      n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, 
      n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, 
      n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, 
      n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, 
      n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, 
      n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, 
      n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, 
      n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, 
      n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, 
      n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, 
      n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, 
      n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, 
      n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, 
      n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, 
      n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, 
      n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, 
      n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, 
      n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, 
      n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, 
      n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, 
      n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, 
      n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, 
      n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, 
      n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, 
      n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, 
      n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, 
      n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, 
      n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, 
      n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, 
      n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, 
      n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, 
      n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, 
      n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, 
      n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, 
      n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, 
      n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, 
      n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, 
      n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, 
      n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, 
      n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, 
      n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, 
      n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, 
      n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, 
      n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, 
      n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, 
      n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, 
      n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, 
      n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, 
      n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, 
      n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, 
      n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, 
      n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, 
      n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, 
      n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, 
      n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, 
      n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, 
      n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, 
      n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, 
      n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, 
      n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, 
      n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, 
      n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, 
      n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, 
      n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, 
      n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, 
      n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, 
      n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, 
      n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, 
      n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, 
      n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, 
      n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, 
      n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, 
      n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, 
      n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, 
      n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, 
      n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, 
      n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, 
      n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, 
      n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, 
      n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, 
      n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, 
      n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, 
      n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, 
      n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, 
      n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, 
      n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, 
      n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, 
      n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, 
      n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, 
      n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, 
      n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, 
      n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, 
      n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, 
      n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, 
      n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, 
      n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, 
      n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, 
      n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, 
      n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, 
      n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, 
      n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, 
      n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, 
      n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, 
      n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, 
      n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, 
      n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, 
      n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, 
      n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, 
      n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, 
      n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, 
      n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, 
      n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, 
      n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, 
      n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, 
      n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, 
      n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, 
      n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, 
      n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, 
      n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, 
      n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, 
      n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, 
      n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, 
      n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, 
      n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, 
      n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, 
      n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, 
      n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, 
      n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, 
      n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, 
      n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, 
      n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, 
      n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, 
      n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, 
      n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, 
      n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, 
      n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, 
      n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, 
      n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, 
      n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, 
      n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, 
      n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, 
      n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, 
      n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, 
      n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, 
      n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, 
      n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, 
      n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, 
      n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, 
      n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, 
      n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, 
      n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, 
      n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, 
      n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, 
      n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, 
      n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, 
      n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, 
      n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, 
      n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, 
      n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, 
      n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, 
      n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, 
      n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, 
      n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, 
      n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, 
      n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, 
      n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, 
      n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, 
      n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, 
      n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, 
      n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, 
      n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, 
      n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, 
      n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, 
      n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, 
      n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, 
      n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, 
      n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, 
      n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, 
      n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, 
      n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, 
      n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, 
      n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, 
      n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, 
      n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, 
      n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, 
      n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, 
      n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, 
      n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, 
      n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, 
      n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, 
      n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, 
      n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, 
      n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, 
      n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, 
      n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, 
      n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, 
      n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, 
      n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, 
      n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, 
      n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, 
      n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, 
      n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, 
      n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, 
      n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, 
      n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, 
      n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, 
      n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, 
      n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, 
      n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, 
      n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, 
      n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, 
      n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, 
      n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, 
      n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, 
      n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, 
      n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, 
      n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, 
      n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, 
      n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, 
      n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, 
      n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, 
      n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, 
      n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, 
      n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, 
      n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, 
      n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, 
      n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, 
      n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, 
      n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, 
      n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, 
      n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, 
      n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, 
      n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, 
      n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, 
      n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, 
      n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, 
      n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, 
      n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, 
      n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, 
      n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, 
      n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, 
      n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, 
      n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, 
      n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, 
      n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, 
      n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, 
      n18051, n18052, n18053, n18054, n18055, net271227, net271228, net271229, 
      net271230, net271231, net271232, net271233, net271234, net271235, 
      net271236, net271237, net271238, net271239, net271240, net271241, 
      net271242, net271243, net271244, net271245, net271246, net271247, 
      net271248, net271249, net271250, net271251, net271252, net271253, 
      net271254, net271255, net271256, net271257, net271258, net271259, 
      net271260, net271261, net271262, net271263, net271264, net271265, 
      net271266, net271267, net271268, net271269, net271270, net271271, 
      net271272, net271273, net271274, net271275, net271276, net271277, 
      net271278, net271279, net271280, net271281, net271282, net271283, 
      net271284, net271285, net271286, net271287, net271288, net271289, 
      net271290, net271291, net271292, net271293, net271294, net271295, 
      net271296, net271297, net271298, net271299, net271300, net271301, 
      net271302, net271303, net271304, net271305, net271306, net271307, 
      net271308, net271309, net271310, net271311, net271312, net271313, 
      net271314, net271315, net271316, net271317, net271318, net271319, 
      net271320, net271321, net271322, net271323, net271324, net271325, 
      net271326, net271327, net271328, net271329, net271330, net271331, 
      net271332, net271333, net271334, net271335, net271336, net271337, 
      net271338, net271339, net271340, net271341, net271342, net271343, 
      net271344, net271345, net271346, net271347, net271348, net271349, 
      net271350, net271351, net271352, net271353, net271354, net271355, 
      net271356, net271357, net271358, net271359, net271360, net271361, 
      net271362, net271363, net271364, net271365, net271366, net271367, 
      net271368, net271369, net271370, net271371, net271372, net271373, 
      net271374, net271375, net271376, net271377, net271378, net271379, 
      net271380, net271381, net271382, net271383, net271384, net271385, 
      net271386, net271387, net271388, net271389, net271390, net271391, 
      net271392, net271393, net271394, net271395, net271396, net271397, 
      net271398, net271399, net271400, net271401, net271402, net271403, 
      net271404, net271405, net271406, net271407, net271408, net271409, 
      net271410, net271411, net271412, net271413, net271414, net271415, 
      net271416, net271417, net271418, net271419, net271420, net271421, 
      net271422, net271423, net271424, net271425, net271426, net271427, 
      net271428, net271429, net271430, net271431, net271432, net271433, 
      net271434, net271435, net271436, net271437, net271438, net271439, 
      net271440, net271441, net271442, net271443, net271444, net271445, 
      net271446, net271447, net271448, net271449, net271450, net271451, 
      net271452, net271453, net271454, net271455, net271456, net271457, 
      net271458, net271459, net271460, net271461, net271462, net271463, 
      net271464, net271465, net271466, net271467, net271468, net271469, 
      net271470, net271471, net271472, net271473, net271474, net271475, 
      net271476, net271477, net271478, net271479, net271480, net271481, 
      net271482, net271483, net271484, net271485, net271486, net271487, 
      net271488, net271489, net271490, net271491, net271492, net271493, 
      net271494, net271495, net271496, net271497, net271498, net271499, 
      net271500, net271501, net271502, net271503, net271504, net271505, 
      net271506, net271507, net271508, net271509, net271510, net271511, 
      net271512, net271513, net271514, net271515, net271516, net271517, 
      net271518, net271519, net271520, net271521, net271522, net271523, 
      net271524, net271525, net271526, net271527, net271528, net271529, 
      net271530, net271531, net271532, net271533, net271534, net271535, 
      net271536, net271537, net271538, net271539, net271540, net271541, 
      net271542, net271543, net271544, net271545, net271546, net271547, 
      net271548, net271549, net271550, net271551, net271552, net271553, 
      net271554, net271555, net271556, net271557, net271558, net271559, 
      net271560, net271561, net271562, net271563, net271564, net271565, 
      net271566, net271567, net271568, net271569, net271570, net271571, 
      net271572, net271573, net271574, net271575, net271576, net271577, 
      net271578, net271579, net271580, net271581, net271582, net271583, 
      net271584, net271585, net271586, net271587, net271588, net271589, 
      net271590, net271591, net271592, net271593, net271594, net271595, 
      net271596, net271597, net271598, net271599, net271600, net271601, 
      net271602, net271603, net271604, net271605 : std_logic;

begin
   
   imspilling_reg : DFF_X1 port map( D => n10185, CK => clk, Q => spill, QN => 
                           n14821);
   swp_reg_0_inst : DFF_X1 port map( D => n10184, CK => clk, Q => swp_0_port, 
                           QN => net271605);
   imfilling_reg : DFF_X1 port map( D => n10183, CK => clk, Q => fill, QN => 
                           n5522);
   cwp_reg_5_inst : DFF_X1 port map( D => n10181, CK => clk, Q => N51637, QN =>
                           n3043);
   swp_reg_1_inst : DFF_X1 port map( D => n10178, CK => clk, Q => swp_1_port, 
                           QN => net271604);
   swp_reg_2_inst : DFF_X1 port map( D => n10176, CK => clk, Q => swp_2_port, 
                           QN => net271603);
   swp_reg_3_inst : DFF_X1 port map( D => n10174, CK => clk, Q => swp_3_port, 
                           QN => net271602);
   swp_reg_5_inst : DFF_X1 port map( D => n10173, CK => clk, Q => swp_5_port, 
                           QN => net271601);
   swp_reg_4_inst : DFF_X1 port map( D => n10172, CK => clk, Q => swp_4_port, 
                           QN => net271600);
   to_mem_tri_enable_reg_31_inst : DFF_X1 port map( D => n10171, CK => clk, Q 
                           => n6613, QN => n7662);
   to_mem_tri_enable_reg_30_inst : DFF_X1 port map( D => n10170, CK => clk, Q 
                           => n6620, QN => n7663);
   to_mem_tri_enable_reg_29_inst : DFF_X1 port map( D => n10169, CK => clk, Q 
                           => n6621, QN => n7664);
   to_mem_tri_enable_reg_28_inst : DFF_X1 port map( D => n10168, CK => clk, Q 
                           => n6624, QN => n7665);
   to_mem_tri_enable_reg_27_inst : DFF_X1 port map( D => n10167, CK => clk, Q 
                           => n6630, QN => n7666);
   to_mem_tri_enable_reg_26_inst : DFF_X1 port map( D => n10166, CK => clk, Q 
                           => n6632, QN => n7667);
   to_mem_tri_enable_reg_25_inst : DFF_X1 port map( D => n10165, CK => clk, Q 
                           => n6634, QN => n7668);
   to_mem_tri_enable_reg_24_inst : DFF_X1 port map( D => n10164, CK => clk, Q 
                           => n6641, QN => n7669);
   to_mem_tri_enable_reg_23_inst : DFF_X1 port map( D => n10163, CK => clk, Q 
                           => n6642, QN => n7670);
   to_mem_tri_enable_reg_22_inst : DFF_X1 port map( D => n10162, CK => clk, Q 
                           => n6646, QN => n7671);
   to_mem_tri_enable_reg_21_inst : DFF_X1 port map( D => n10161, CK => clk, Q 
                           => n6647, QN => n7672);
   to_mem_tri_enable_reg_20_inst : DFF_X1 port map( D => n10160, CK => clk, Q 
                           => n6648, QN => n7673);
   to_mem_tri_enable_reg_19_inst : DFF_X1 port map( D => n10159, CK => clk, Q 
                           => n6649, QN => n7674);
   to_mem_tri_enable_reg_18_inst : DFF_X1 port map( D => n10158, CK => clk, Q 
                           => n6650, QN => n7675);
   to_mem_tri_enable_reg_17_inst : DFF_X1 port map( D => n10157, CK => clk, Q 
                           => n6651, QN => n7676);
   to_mem_tri_enable_reg_16_inst : DFF_X1 port map( D => n10156, CK => clk, Q 
                           => n6652, QN => n7677);
   to_mem_tri_enable_reg_15_inst : DFF_X1 port map( D => n10155, CK => clk, Q 
                           => n6653, QN => n7678);
   to_mem_tri_enable_reg_14_inst : DFF_X1 port map( D => n10154, CK => clk, Q 
                           => n6654, QN => n7679);
   to_mem_tri_enable_reg_13_inst : DFF_X1 port map( D => n10153, CK => clk, Q 
                           => n6655, QN => n7680);
   to_mem_tri_enable_reg_12_inst : DFF_X1 port map( D => n10152, CK => clk, Q 
                           => n6656, QN => n7681);
   to_mem_tri_enable_reg_11_inst : DFF_X1 port map( D => n10151, CK => clk, Q 
                           => n6657, QN => n7682);
   to_mem_tri_enable_reg_10_inst : DFF_X1 port map( D => n10150, CK => clk, Q 
                           => n6658, QN => n7683);
   to_mem_tri_enable_reg_9_inst : DFF_X1 port map( D => n10149, CK => clk, Q =>
                           n6659, QN => n7684);
   to_mem_tri_enable_reg_8_inst : DFF_X1 port map( D => n10148, CK => clk, Q =>
                           n6660, QN => n7685);
   to_mem_tri_enable_reg_7_inst : DFF_X1 port map( D => n10147, CK => clk, Q =>
                           n6671, QN => n7686);
   to_mem_tri_enable_reg_6_inst : DFF_X1 port map( D => n10146, CK => clk, Q =>
                           n6674, QN => n7687);
   to_mem_tri_enable_reg_5_inst : DFF_X1 port map( D => n10145, CK => clk, Q =>
                           n6676, QN => n7688);
   to_mem_tri_enable_reg_4_inst : DFF_X1 port map( D => n10144, CK => clk, Q =>
                           n6683, QN => n7689);
   to_mem_tri_enable_reg_3_inst : DFF_X1 port map( D => n10143, CK => clk, Q =>
                           n6684, QN => n7690);
   to_mem_tri_enable_reg_2_inst : DFF_X1 port map( D => n10142, CK => clk, Q =>
                           n6687, QN => n7691);
   to_mem_tri_enable_reg_1_inst : DFF_X1 port map( D => n10141, CK => clk, Q =>
                           n6693, QN => n7692);
   to_mem_tri_enable_reg_0_inst : DFF_X1 port map( D => n10140, CK => clk, Q =>
                           n6695, QN => n7693);
   i_reg_0_inst : DFF_X1 port map( D => n10138, CK => clk, Q => i_0_port, QN =>
                           net227476);
   i_reg_5_inst : DFF_X1 port map( D => n10137, CK => clk, Q => i_5_port, QN =>
                           net227475);
   i_reg_1_inst : DFF_X1 port map( D => n10136, CK => clk, Q => i_1_port, QN =>
                           net227474);
   i_reg_2_inst : DFF_X1 port map( D => n10135, CK => clk, Q => i_2_port, QN =>
                           net227473);
   i_reg_3_inst : DFF_X1 port map( D => n10134, CK => clk, Q => i_3_port, QN =>
                           net227472);
   i_reg_4_inst : DFF_X1 port map( D => n10133, CK => clk, Q => i_4_port, QN =>
                           net227471);
   lastcwp_reg_5_inst : DFF_X1 port map( D => n10132, CK => clk, Q => net271599
                           , QN => n7592);
   lastcwp_reg_4_inst : DFF_X1 port map( D => n10131, CK => clk, Q => 
                           lastcwp_4_port, QN => n7591);
   lastcwp_reg_3_inst : DFF_X1 port map( D => n10130, CK => clk, Q => 
                           lastcwp_3_port, QN => n7590);
   lastcwp_reg_2_inst : DFF_X1 port map( D => n10129, CK => clk, Q => 
                           lastcwp_2_port, QN => n7589);
   lastcwp_reg_1_inst : DFF_X1 port map( D => n10128, CK => clk, Q => 
                           lastcwp_1_port, QN => n7588);
   lastcwp_reg_0_inst : DFF_X1 port map( D => n10127, CK => clk, Q => net271598
                           , QN => n7587);
   registers_reg_0_31_inst : DFF_X1 port map( D => n10125, CK => clk, Q => 
                           registers_0_31_port, QN => n15801);
   registers_reg_1_31_inst : DFF_X1 port map( D => n10124, CK => clk, Q => 
                           registers_1_31_port, QN => n15585);
   registers_reg_2_31_inst : DFF_X1 port map( D => n10123, CK => clk, Q => 
                           registers_2_31_port, QN => n14815);
   registers_reg_3_31_inst : DFF_X1 port map( D => n10122, CK => clk, Q => 
                           net227470, QN => n15781);
   registers_reg_4_31_inst : DFF_X1 port map( D => n10121, CK => clk, Q => 
                           registers_4_31_port, QN => n15458);
   registers_reg_5_31_inst : DFF_X1 port map( D => n10120, CK => clk, Q => 
                           registers_5_31_port, QN => n15318);
   registers_reg_6_31_inst : DFF_X1 port map( D => n10119, CK => clk, Q => 
                           net271597, QN => n12348);
   registers_reg_7_31_inst : DFF_X1 port map( D => n10118, CK => clk, Q => 
                           registers_7_31_port, QN => n15349);
   registers_reg_8_31_inst : DFF_X1 port map( D => n10117, CK => clk, Q => 
                           net227469, QN => n15239);
   registers_reg_9_31_inst : DFF_X1 port map( D => n10116, CK => clk, Q => 
                           registers_9_31_port, QN => n14358);
   registers_reg_10_31_inst : DFF_X1 port map( D => n10115, CK => clk, Q => 
                           registers_10_31_port, QN => n14756);
   registers_reg_11_31_inst : DFF_X1 port map( D => n10114, CK => clk, Q => 
                           registers_11_31_port, QN => n14425);
   registers_reg_12_31_inst : DFF_X1 port map( D => n10113, CK => clk, Q => 
                           registers_12_31_port, QN => n15691);
   registers_reg_13_31_inst : DFF_X1 port map( D => n10112, CK => clk, Q => 
                           net227468, QN => n15071);
   registers_reg_14_31_inst : DFF_X1 port map( D => n10111, CK => clk, Q => 
                           net271596, QN => n11903);
   registers_reg_15_31_inst : DFF_X1 port map( D => n10110, CK => clk, Q => 
                           registers_15_31_port, QN => n15314);
   registers_reg_16_31_inst : DFF_X1 port map( D => n10109, CK => clk, Q => 
                           registers_16_31_port, QN => n15721);
   registers_reg_17_31_inst : DFF_X1 port map( D => n10108, CK => clk, Q => 
                           registers_17_31_port, QN => n14627);
   registers_reg_18_31_inst : DFF_X1 port map( D => n10107, CK => clk, Q => 
                           registers_18_31_port, QN => n14371);
   registers_reg_19_31_inst : DFF_X1 port map( D => n10106, CK => clk, Q => 
                           registers_19_31_port, QN => n15814);
   registers_reg_20_31_inst : DFF_X1 port map( D => n10105, CK => clk, Q => 
                           net271595, QN => n14853);
   registers_reg_21_31_inst : DFF_X1 port map( D => n10104, CK => clk, Q => 
                           net271594, QN => n12307);
   registers_reg_22_31_inst : DFF_X1 port map( D => n10103, CK => clk, Q => 
                           registers_22_31_port, QN => n15377);
   registers_reg_23_31_inst : DFF_X1 port map( D => n10102, CK => clk, Q => 
                           registers_23_31_port, QN => n15889);
   registers_reg_24_31_inst : DFF_X1 port map( D => n10101, CK => clk, Q => 
                           net227467, QN => n15209);
   registers_reg_25_31_inst : DFF_X1 port map( D => n10100, CK => clk, Q => 
                           registers_25_31_port, QN => n14328);
   registers_reg_26_31_inst : DFF_X1 port map( D => n10099, CK => clk, Q => 
                           net271593, QN => n12355);
   registers_reg_27_31_inst : DFF_X1 port map( D => n10098, CK => clk, Q => 
                           net271592, QN => n12047);
   registers_reg_28_31_inst : DFF_X1 port map( D => n10097, CK => clk, Q => 
                           net227466, QN => n15032);
   registers_reg_29_31_inst : DFF_X1 port map( D => n10096, CK => clk, Q => 
                           registers_29_31_port, QN => n15813);
   registers_reg_30_31_inst : DFF_X1 port map( D => n10095, CK => clk, Q => 
                           registers_30_31_port, QN => n14699);
   registers_reg_31_31_inst : DFF_X1 port map( D => n10094, CK => clk, Q => 
                           net227465, QN => n15757);
   registers_reg_32_31_inst : DFF_X1 port map( D => n10093, CK => clk, Q => 
                           net271591, QN => n12314);
   registers_reg_33_31_inst : DFF_X1 port map( D => n10092, CK => clk, Q => 
                           net271590, QN => n11845);
   registers_reg_34_31_inst : DFF_X1 port map( D => n10091, CK => clk, Q => 
                           registers_34_31_port, QN => n15517);
   registers_reg_35_31_inst : DFF_X1 port map( D => n10090, CK => clk, Q => 
                           net227464, QN => n15590);
   registers_reg_36_31_inst : DFF_X1 port map( D => n10089, CK => clk, Q => 
                           registers_36_31_port, QN => n15156);
   registers_reg_37_31_inst : DFF_X1 port map( D => n10088, CK => clk, Q => 
                           registers_37_31_port, QN => n14370);
   registers_reg_38_31_inst : DFF_X1 port map( D => n10087, CK => clk, Q => 
                           registers_38_31_port, QN => n15041);
   registers_reg_39_31_inst : DFF_X1 port map( D => n10086, CK => clk, Q => 
                           net271589, QN => n12194);
   registers_reg_40_31_inst : DFF_X1 port map( D => n10085, CK => clk, Q => 
                           registers_40_31_port, QN => n15150);
   registers_reg_41_31_inst : DFF_X1 port map( D => n10084, CK => clk, Q => 
                           registers_41_31_port, QN => n14533);
   registers_reg_42_31_inst : DFF_X1 port map( D => n10083, CK => clk, Q => 
                           registers_42_31_port, QN => n15926);
   registers_reg_43_31_inst : DFF_X1 port map( D => n10082, CK => clk, Q => 
                           registers_43_31_port, QN => n14887);
   registers_reg_44_31_inst : DFF_X1 port map( D => n10081, CK => clk, Q => 
                           registers_44_31_port, QN => n15487);
   registers_reg_45_31_inst : DFF_X1 port map( D => n10080, CK => clk, Q => 
                           registers_45_31_port, QN => n14816);
   registers_reg_46_31_inst : DFF_X1 port map( D => n10079, CK => clk, Q => 
                           net227463, QN => n11950);
   registers_reg_47_31_inst : DFF_X1 port map( D => n10078, CK => clk, Q => 
                           registers_47_31_port, QN => n14546);
   registers_reg_48_31_inst : DFF_X1 port map( D => n10077, CK => clk, Q => 
                           registers_48_31_port, QN => n15551);
   registers_reg_49_31_inst : DFF_X1 port map( D => n10076, CK => clk, Q => 
                           registers_49_31_port, QN => n14477);
   registers_reg_50_31_inst : DFF_X1 port map( D => n10075, CK => clk, Q => 
                           registers_50_31_port, QN => n15975);
   registers_reg_51_31_inst : DFF_X1 port map( D => n10074, CK => clk, Q => 
                           registers_51_31_port, QN => n15427);
   registers_reg_52_31_inst : DFF_X1 port map( D => n10073, CK => clk, Q => 
                           net227462, QN => n14937);
   registers_reg_53_31_inst : DFF_X1 port map( D => n10072, CK => clk, Q => 
                           net227461, QN => n15920);
   registers_reg_54_31_inst : DFF_X1 port map( D => n10071, CK => clk, Q => 
                           registers_54_31_port, QN => n14535);
   registers_reg_55_31_inst : DFF_X1 port map( D => n10070, CK => clk, Q => 
                           registers_55_31_port, QN => n12049);
   registers_reg_56_31_inst : DFF_X1 port map( D => n10069, CK => clk, Q => 
                           registers_56_31_port, QN => n15790);
   registers_reg_57_31_inst : DFF_X1 port map( D => n10068, CK => clk, Q => 
                           net227460, QN => n15034);
   registers_reg_58_31_inst : DFF_X1 port map( D => n10067, CK => clk, Q => 
                           net227459, QN => n14859);
   registers_reg_59_31_inst : DFF_X1 port map( D => n10066, CK => clk, Q => 
                           registers_59_31_port, QN => n14670);
   registers_reg_60_31_inst : DFF_X1 port map( D => n10065, CK => clk, Q => 
                           registers_60_31_port, QN => n14634);
   registers_reg_61_31_inst : DFF_X1 port map( D => n10064, CK => clk, Q => 
                           net227458, QN => n15317);
   registers_reg_62_31_inst : DFF_X1 port map( D => n10063, CK => clk, Q => 
                           registers_62_31_port, QN => n14992);
   registers_reg_63_31_inst : DFF_X1 port map( D => n10062, CK => clk, Q => 
                           registers_63_31_port, QN => n14281);
   to_mem_reg_31_inst : DFF_X1 port map( D => n10061, CK => clk, Q => net271588
                           , QN => n7694);
   registers_reg_64_31_inst : DFF_X1 port map( D => n10060, CK => clk, Q => 
                           net227457, QN => n16034);
   registers_reg_65_31_inst : DFF_X1 port map( D => n10059, CK => clk, Q => 
                           net227456, QN => n16028);
   registers_reg_66_31_inst : DFF_X1 port map( D => n10058, CK => clk, Q => 
                           net227455, QN => n16029);
   registers_reg_67_31_inst : DFF_X1 port map( D => n10057, CK => clk, Q => 
                           net271587, QN => n14856);
   registers_reg_68_31_inst : DFF_X1 port map( D => n10056, CK => clk, Q => 
                           registers_68_31_port, QN => n16035);
   registers_reg_69_31_inst : DFF_X1 port map( D => n10055, CK => clk, Q => 
                           net227454, QN => n16033);
   registers_reg_70_31_inst : DFF_X1 port map( D => n10054, CK => clk, Q => 
                           net227453, QN => n16123);
   registers_reg_0_30_inst : DFF_X1 port map( D => n10053, CK => clk, Q => 
                           registers_0_30_port, QN => n15785);
   registers_reg_1_30_inst : DFF_X1 port map( D => n10052, CK => clk, Q => 
                           registers_1_30_port, QN => n15279);
   registers_reg_2_30_inst : DFF_X1 port map( D => n10051, CK => clk, Q => 
                           registers_2_30_port, QN => n14630);
   registers_reg_3_30_inst : DFF_X1 port map( D => n10050, CK => clk, Q => 
                           net227452, QN => n15283);
   registers_reg_4_30_inst : DFF_X1 port map( D => n10049, CK => clk, Q => 
                           registers_4_30_port, QN => n15274);
   registers_reg_5_30_inst : DFF_X1 port map( D => n10048, CK => clk, Q => 
                           registers_5_30_port, QN => n14632);
   registers_reg_6_30_inst : DFF_X1 port map( D => n10047, CK => clk, Q => 
                           net271586, QN => n12196);
   registers_reg_7_30_inst : DFF_X1 port map( D => n10046, CK => clk, Q => 
                           registers_7_30_port, QN => n15271);
   registers_reg_8_30_inst : DFF_X1 port map( D => n10045, CK => clk, Q => 
                           net227451, QN => n14874);
   registers_reg_9_30_inst : DFF_X1 port map( D => n10044, CK => clk, Q => 
                           registers_9_30_port, QN => n14055);
   registers_reg_10_30_inst : DFF_X1 port map( D => n10043, CK => clk, Q => 
                           registers_10_30_port, QN => n14629);
   registers_reg_11_30_inst : DFF_X1 port map( D => n10042, CK => clk, Q => 
                           registers_11_30_port, QN => n14060);
   registers_reg_12_30_inst : DFF_X1 port map( D => n10041, CK => clk, Q => 
                           registers_12_30_port, QN => n15280);
   registers_reg_13_30_inst : DFF_X1 port map( D => n10040, CK => clk, Q => 
                           net227450, QN => n14870);
   registers_reg_14_30_inst : DFF_X1 port map( D => n10039, CK => clk, Q => 
                           net271585, QN => n11541);
   registers_reg_15_30_inst : DFF_X1 port map( D => n10038, CK => clk, Q => 
                           registers_15_30_port, QN => n15270);
   registers_reg_16_30_inst : DFF_X1 port map( D => n10037, CK => clk, Q => 
                           registers_16_30_port, QN => n15281);
   registers_reg_17_30_inst : DFF_X1 port map( D => n10036, CK => clk, Q => 
                           registers_17_30_port, QN => n14299);
   registers_reg_18_30_inst : DFF_X1 port map( D => n10035, CK => clk, Q => 
                           registers_18_30_port, QN => n14057);
   registers_reg_19_30_inst : DFF_X1 port map( D => n10034, CK => clk, Q => 
                           registers_19_30_port, QN => n15784);
   registers_reg_20_30_inst : DFF_X1 port map( D => n10033, CK => clk, Q => 
                           net271584, QN => n14822);
   registers_reg_21_30_inst : DFF_X1 port map( D => n10032, CK => clk, Q => 
                           net271583, QN => n12161);
   registers_reg_22_30_inst : DFF_X1 port map( D => n10031, CK => clk, Q => 
                           registers_22_30_port, QN => n15273);
   registers_reg_23_30_inst : DFF_X1 port map( D => n10030, CK => clk, Q => 
                           registers_23_30_port, QN => n15786);
   registers_reg_24_30_inst : DFF_X1 port map( D => n10029, CK => clk, Q => 
                           net227449, QN => n14873);
   registers_reg_25_30_inst : DFF_X1 port map( D => n10028, CK => clk, Q => 
                           registers_25_30_port, QN => n14054);
   registers_reg_26_30_inst : DFF_X1 port map( D => n10027, CK => clk, Q => 
                           net271582, QN => n12197);
   registers_reg_27_30_inst : DFF_X1 port map( D => n10026, CK => clk, Q => 
                           net271581, QN => n11904);
   registers_reg_28_30_inst : DFF_X1 port map( D => n10025, CK => clk, Q => 
                           net227448, QN => n14857);
   registers_reg_29_30_inst : DFF_X1 port map( D => n10024, CK => clk, Q => 
                           registers_29_30_port, QN => n15783);
   registers_reg_30_30_inst : DFF_X1 port map( D => n10023, CK => clk, Q => 
                           registers_30_30_port, QN => n14628);
   registers_reg_31_30_inst : DFF_X1 port map( D => n10022, CK => clk, Q => 
                           net227447, QN => n15282);
   registers_reg_32_30_inst : DFF_X1 port map( D => n10021, CK => clk, Q => 
                           net271580, QN => n12163);
   registers_reg_33_30_inst : DFF_X1 port map( D => n10020, CK => clk, Q => 
                           net271579, QN => n11498);
   registers_reg_34_30_inst : DFF_X1 port map( D => n10019, CK => clk, Q => 
                           registers_34_30_port, QN => n15276);
   registers_reg_35_30_inst : DFF_X1 port map( D => n10018, CK => clk, Q => 
                           net227446, QN => n15278);
   registers_reg_36_30_inst : DFF_X1 port map( D => n10017, CK => clk, Q => 
                           registers_36_30_port, QN => n14872);
   registers_reg_37_30_inst : DFF_X1 port map( D => n10016, CK => clk, Q => 
                           registers_37_30_port, QN => n14056);
   registers_reg_38_30_inst : DFF_X1 port map( D => n10015, CK => clk, Q => 
                           registers_38_30_port, QN => n14869);
   registers_reg_39_30_inst : DFF_X1 port map( D => n10014, CK => clk, Q => 
                           net271578, QN => n12160);
   registers_reg_40_30_inst : DFF_X1 port map( D => n10013, CK => clk, Q => 
                           registers_40_30_port, QN => n14871);
   registers_reg_41_30_inst : DFF_X1 port map( D => n10012, CK => clk, Q => 
                           registers_41_30_port, QN => n14069);
   registers_reg_42_30_inst : DFF_X1 port map( D => n10011, CK => clk, Q => 
                           registers_42_30_port, QN => n15787);
   registers_reg_43_30_inst : DFF_X1 port map( D => n10010, CK => clk, Q => 
                           registers_43_30_port, QN => n14854);
   registers_reg_44_30_inst : DFF_X1 port map( D => n10009, CK => clk, Q => 
                           registers_44_30_port, QN => n15275);
   registers_reg_45_30_inst : DFF_X1 port map( D => n10008, CK => clk, Q => 
                           registers_45_30_port, QN => n14631);
   registers_reg_46_30_inst : DFF_X1 port map( D => n10007, CK => clk, Q => 
                           net227445, QN => n11670);
   registers_reg_47_30_inst : DFF_X1 port map( D => n10006, CK => clk, Q => 
                           registers_47_30_port, QN => n14279);
   registers_reg_48_30_inst : DFF_X1 port map( D => n10005, CK => clk, Q => 
                           registers_48_30_port, QN => n15277);
   registers_reg_49_30_inst : DFF_X1 port map( D => n10004, CK => clk, Q => 
                           registers_49_30_port, QN => n14065);
   registers_reg_50_30_inst : DFF_X1 port map( D => n10003, CK => clk, Q => 
                           registers_50_30_port, QN => n15788);
   registers_reg_51_30_inst : DFF_X1 port map( D => n10002, CK => clk, Q => 
                           registers_51_30_port, QN => n15272);
   registers_reg_52_30_inst : DFF_X1 port map( D => n10001, CK => clk, Q => 
                           net227444, QN => n14855);
   registers_reg_53_30_inst : DFF_X1 port map( D => n10000, CK => clk, Q => 
                           net227443, QN => n15782);
   registers_reg_54_30_inst : DFF_X1 port map( D => n9999, CK => clk, Q => 
                           registers_54_30_port, QN => n14534);
   registers_reg_55_30_inst : DFF_X1 port map( D => n9998, CK => clk, Q => 
                           registers_55_30_port, QN => n12048);
   registers_reg_56_30_inst : DFF_X1 port map( D => n9997, CK => clk, Q => 
                           registers_56_30_port, QN => n15789);
   registers_reg_57_30_inst : DFF_X1 port map( D => n9996, CK => clk, Q => 
                           net227442, QN => n15033);
   registers_reg_58_30_inst : DFF_X1 port map( D => n9995, CK => clk, Q => 
                           net227441, QN => n14858);
   registers_reg_59_30_inst : DFF_X1 port map( D => n9994, CK => clk, Q => 
                           registers_59_30_port, QN => n15315);
   registers_reg_60_30_inst : DFF_X1 port map( D => n9993, CK => clk, Q => 
                           registers_60_30_port, QN => n14633);
   registers_reg_61_30_inst : DFF_X1 port map( D => n9992, CK => clk, Q => 
                           net227440, QN => n15316);
   registers_reg_62_30_inst : DFF_X1 port map( D => n9991, CK => clk, Q => 
                           registers_62_30_port, QN => n14991);
   registers_reg_63_30_inst : DFF_X1 port map( D => n9990, CK => clk, Q => 
                           registers_63_30_port, QN => n14280);
   to_mem_reg_30_inst : DFF_X1 port map( D => n9989, CK => clk, Q => net271577,
                           QN => n7695);
   registers_reg_64_30_inst : DFF_X1 port map( D => n9988, CK => clk, Q => 
                           net227439, QN => n16031);
   registers_reg_65_30_inst : DFF_X1 port map( D => n9987, CK => clk, Q => 
                           net227438, QN => n16027);
   registers_reg_66_30_inst : DFF_X1 port map( D => n9986, CK => clk, Q => 
                           net227437, QN => n16026);
   registers_reg_67_30_inst : DFF_X1 port map( D => n9985, CK => clk, Q => 
                           net271576, QN => n14052);
   registers_reg_68_30_inst : DFF_X1 port map( D => n9984, CK => clk, Q => 
                           registers_68_30_port, QN => n16032);
   registers_reg_69_30_inst : DFF_X1 port map( D => n9983, CK => clk, Q => 
                           net227436, QN => n16030);
   registers_reg_70_30_inst : DFF_X1 port map( D => n9982, CK => clk, Q => 
                           net227435, QN => n16025);
   registers_reg_0_29_inst : DFF_X1 port map( D => n9981, CK => clk, Q => 
                           registers_0_29_port, QN => n15880);
   registers_reg_1_29_inst : DFF_X1 port map( D => n9980, CK => clk, Q => 
                           registers_1_29_port, QN => n15615);
   registers_reg_2_29_inst : DFF_X1 port map( D => n9979, CK => clk, Q => 
                           registers_2_29_port, QN => n14769);
   registers_reg_3_29_inst : DFF_X1 port map( D => n9978, CK => clk, Q => 
                           net227434, QN => n15735);
   registers_reg_4_29_inst : DFF_X1 port map( D => n9977, CK => clk, Q => 
                           registers_4_29_port, QN => n15457);
   registers_reg_5_29_inst : DFF_X1 port map( D => n9976, CK => clk, Q => 
                           registers_5_29_port, QN => n14709);
   registers_reg_6_29_inst : DFF_X1 port map( D => n9975, CK => clk, Q => 
                           net271575, QN => n12347);
   registers_reg_7_29_inst : DFF_X1 port map( D => n9974, CK => clk, Q => 
                           registers_7_29_port, QN => n15325);
   registers_reg_8_29_inst : DFF_X1 port map( D => n9973, CK => clk, Q => 
                           net227433, QN => n15238);
   registers_reg_9_29_inst : DFF_X1 port map( D => n9972, CK => clk, Q => 
                           registers_9_29_port, QN => n14357);
   registers_reg_10_29_inst : DFF_X1 port map( D => n9971, CK => clk, Q => 
                           registers_10_29_port, QN => n14710);
   registers_reg_11_29_inst : DFF_X1 port map( D => n9970, CK => clk, Q => 
                           registers_11_29_port, QN => n14424);
   registers_reg_12_29_inst : DFF_X1 port map( D => n9969, CK => clk, Q => 
                           registers_12_29_port, QN => n15668);
   registers_reg_13_29_inst : DFF_X1 port map( D => n9968, CK => clk, Q => 
                           net227432, QN => n15070);
   registers_reg_14_29_inst : DFF_X1 port map( D => n9967, CK => clk, Q => 
                           net271574, QN => n11880);
   registers_reg_15_29_inst : DFF_X1 port map( D => n9966, CK => clk, Q => 
                           registers_15_29_port, QN => n15291);
   registers_reg_16_29_inst : DFF_X1 port map( D => n9965, CK => clk, Q => 
                           registers_16_29_port, QN => n15698);
   registers_reg_17_29_inst : DFF_X1 port map( D => n9964, CK => clk, Q => 
                           registers_17_29_port, QN => n14604);
   registers_reg_18_29_inst : DFF_X1 port map( D => n9963, CK => clk, Q => 
                           registers_18_29_port, QN => n14397);
   registers_reg_19_29_inst : DFF_X1 port map( D => n9962, CK => clk, Q => 
                           registers_19_29_port, QN => n15840);
   registers_reg_20_29_inst : DFF_X1 port map( D => n9961, CK => clk, Q => 
                           net271573, QN => n14830);
   registers_reg_21_29_inst : DFF_X1 port map( D => n9960, CK => clk, Q => 
                           net271572, QN => n12204);
   registers_reg_22_29_inst : DFF_X1 port map( D => n9959, CK => clk, Q => 
                           registers_22_29_port, QN => n15390);
   registers_reg_23_29_inst : DFF_X1 port map( D => n9958, CK => clk, Q => 
                           registers_23_29_port, QN => n15902);
   registers_reg_24_29_inst : DFF_X1 port map( D => n9957, CK => clk, Q => 
                           net227431, QN => n15208);
   registers_reg_25_29_inst : DFF_X1 port map( D => n9956, CK => clk, Q => 
                           registers_25_29_port, QN => n14327);
   registers_reg_26_29_inst : DFF_X1 port map( D => n9955, CK => clk, Q => 
                           net271571, QN => n12354);
   registers_reg_27_29_inst : DFF_X1 port map( D => n9954, CK => clk, Q => 
                           net271570, QN => n12046);
   registers_reg_28_29_inst : DFF_X1 port map( D => n9953, CK => clk, Q => 
                           net227430, QN => n15031);
   registers_reg_29_29_inst : DFF_X1 port map( D => n9952, CK => clk, Q => 
                           registers_29_29_port, QN => n15839);
   registers_reg_30_29_inst : DFF_X1 port map( D => n9951, CK => clk, Q => 
                           registers_30_29_port, QN => n14677);
   registers_reg_31_29_inst : DFF_X1 port map( D => n9950, CK => clk, Q => 
                           net227429, QN => n15734);
   registers_reg_32_29_inst : DFF_X1 port map( D => n9949, CK => clk, Q => 
                           net271569, QN => n12339);
   registers_reg_33_29_inst : DFF_X1 port map( D => n9948, CK => clk, Q => 
                           net271568, QN => n11861);
   registers_reg_34_29_inst : DFF_X1 port map( D => n9947, CK => clk, Q => 
                           registers_34_29_port, QN => n15494);
   registers_reg_35_29_inst : DFF_X1 port map( D => n9946, CK => clk, Q => 
                           net227428, QN => n15614);
   registers_reg_36_29_inst : DFF_X1 port map( D => n9945, CK => clk, Q => 
                           registers_36_29_port, QN => n15169);
   registers_reg_37_29_inst : DFF_X1 port map( D => n9944, CK => clk, Q => 
                           registers_37_29_port, QN => n14396);
   registers_reg_38_29_inst : DFF_X1 port map( D => n9943, CK => clk, Q => 
                           registers_38_29_port, QN => n15054);
   registers_reg_39_29_inst : DFF_X1 port map( D => n9942, CK => clk, Q => 
                           net271567, QN => n12170);
   registers_reg_40_29_inst : DFF_X1 port map( D => n9941, CK => clk, Q => 
                           registers_40_29_port, QN => n15149);
   registers_reg_41_29_inst : DFF_X1 port map( D => n9940, CK => clk, Q => 
                           registers_41_29_port, QN => n14532);
   registers_reg_42_29_inst : DFF_X1 port map( D => n9939, CK => clk, Q => 
                           registers_42_29_port, QN => n15939);
   registers_reg_43_29_inst : DFF_X1 port map( D => n9938, CK => clk, Q => 
                           registers_43_29_port, QN => n14885);
   registers_reg_44_29_inst : DFF_X1 port map( D => n9937, CK => clk, Q => 
                           registers_44_29_port, QN => n15465);
   registers_reg_45_29_inst : DFF_X1 port map( D => n9936, CK => clk, Q => 
                           registers_45_29_port, QN => n14770);
   registers_reg_46_29_inst : DFF_X1 port map( D => n9935, CK => clk, Q => 
                           net227427, QN => n11949);
   registers_reg_47_29_inst : DFF_X1 port map( D => n9934, CK => clk, Q => 
                           registers_47_29_port, QN => n14545);
   registers_reg_48_29_inst : DFF_X1 port map( D => n9933, CK => clk, Q => 
                           registers_48_29_port, QN => n15550);
   registers_reg_49_29_inst : DFF_X1 port map( D => n9932, CK => clk, Q => 
                           registers_49_29_port, QN => n14476);
   registers_reg_50_29_inst : DFF_X1 port map( D => n9931, CK => clk, Q => 
                           registers_50_29_port, QN => n15988);
   registers_reg_51_29_inst : DFF_X1 port map( D => n9930, CK => clk, Q => 
                           registers_51_29_port, QN => n15426);
   registers_reg_52_29_inst : DFF_X1 port map( D => n9929, CK => clk, Q => 
                           net227426, QN => n14936);
   registers_reg_53_29_inst : DFF_X1 port map( D => n9928, CK => clk, Q => 
                           net227425, QN => n15968);
   registers_reg_54_29_inst : DFF_X1 port map( D => n9927, CK => clk, Q => 
                           registers_54_29_port, QN => n14597);
   registers_reg_55_29_inst : DFF_X1 port map( D => n9926_port, CK => clk, Q =>
                           registers_55_29_port, QN => n12159);
   registers_reg_56_29_inst : DFF_X1 port map( D => n9925_port, CK => clk, Q =>
                           registers_56_29_port, QN => n16012);
   registers_reg_57_29_inst : DFF_X1 port map( D => n9924_port, CK => clk, Q =>
                           net227424, QN => n15269);
   registers_reg_58_29_inst : DFF_X1 port map( D => n9923_port, CK => clk, Q =>
                           net227423, QN => n14886);
   registers_reg_59_29_inst : DFF_X1 port map( D => n9922_port, CK => clk, Q =>
                           registers_59_29_port, QN => n15431);
   registers_reg_60_29_inst : DFF_X1 port map( D => n9921_port, CK => clk, Q =>
                           registers_60_29_port, QN => n14644);
   registers_reg_61_29_inst : DFF_X1 port map( D => n9920, CK => clk, Q => 
                           net227422, QN => n15660);
   registers_reg_62_29_inst : DFF_X1 port map( D => n9919, CK => clk, Q => 
                           registers_62_29_port, QN => n15122);
   registers_reg_63_29_inst : DFF_X1 port map( D => n9918, CK => clk, Q => 
                           registers_63_29_port, QN => n14483);
   to_mem_reg_29_inst : DFF_X1 port map( D => n9917, CK => clk, Q => net271566,
                           QN => n7696);
   registers_reg_64_29_inst : DFF_X1 port map( D => n9916, CK => clk, Q => 
                           net227421, QN => n16148);
   registers_reg_65_29_inst : DFF_X1 port map( D => n9915, CK => clk, Q => 
                           net227420, QN => n16097);
   registers_reg_66_29_inst : DFF_X1 port map( D => n9914, CK => clk, Q => 
                           net227419, QN => n16059);
   registers_reg_67_29_inst : DFF_X1 port map( D => n9913, CK => clk, Q => 
                           net271565, QN => n14278);
   registers_reg_68_29_inst : DFF_X1 port map( D => n9912, CK => clk, Q => 
                           registers_68_29_port, QN => n16185);
   registers_reg_69_29_inst : DFF_X1 port map( D => n9911, CK => clk, Q => 
                           net227418, QN => n16137);
   registers_reg_70_29_inst : DFF_X1 port map( D => n9910_port, CK => clk, Q =>
                           net227417, QN => n16049);
   registers_reg_0_28_inst : DFF_X1 port map( D => n9909_port, CK => clk, Q => 
                           registers_0_28_port, QN => n15879);
   registers_reg_1_28_inst : DFF_X1 port map( D => n9908_port, CK => clk, Q => 
                           registers_1_28_port, QN => n15636);
   registers_reg_2_28_inst : DFF_X1 port map( D => n9907, CK => clk, Q => 
                           registers_2_28_port, QN => n14767);
   registers_reg_3_28_inst : DFF_X1 port map( D => n9906, CK => clk, Q => 
                           net227416, QN => n15733);
   registers_reg_4_28_inst : DFF_X1 port map( D => n9905, CK => clk, Q => 
                           registers_4_28_port, QN => n15456);
   registers_reg_5_28_inst : DFF_X1 port map( D => n9904, CK => clk, Q => 
                           registers_5_28_port, QN => n14707);
   registers_reg_6_28_inst : DFF_X1 port map( D => n9903, CK => clk, Q => 
                           net271564, QN => n12346);
   registers_reg_7_28_inst : DFF_X1 port map( D => n9902, CK => clk, Q => 
                           registers_7_28_port, QN => n15324);
   registers_reg_8_28_inst : DFF_X1 port map( D => n9901, CK => clk, Q => 
                           net227415, QN => n15237);
   registers_reg_9_28_inst : DFF_X1 port map( D => n9900, CK => clk, Q => 
                           registers_9_28_port, QN => n14356);
   registers_reg_10_28_inst : DFF_X1 port map( D => n9899, CK => clk, Q => 
                           registers_10_28_port, QN => n14708);
   registers_reg_11_28_inst : DFF_X1 port map( D => n9898, CK => clk, Q => 
                           registers_11_28_port, QN => n14423);
   registers_reg_12_28_inst : DFF_X1 port map( D => n9897, CK => clk, Q => 
                           registers_12_28_port, QN => n15667);
   registers_reg_13_28_inst : DFF_X1 port map( D => n9896, CK => clk, Q => 
                           net227414, QN => n15069);
   registers_reg_14_28_inst : DFF_X1 port map( D => n9895, CK => clk, Q => 
                           net271563, QN => n11879);
   registers_reg_15_28_inst : DFF_X1 port map( D => n9894, CK => clk, Q => 
                           registers_15_28_port, QN => n15290);
   registers_reg_16_28_inst : DFF_X1 port map( D => n9893, CK => clk, Q => 
                           registers_16_28_port, QN => n15697);
   registers_reg_17_28_inst : DFF_X1 port map( D => n9892, CK => clk, Q => 
                           registers_17_28_port, QN => n14603);
   registers_reg_18_28_inst : DFF_X1 port map( D => n9891, CK => clk, Q => 
                           registers_18_28_port, QN => n14418);
   registers_reg_19_28_inst : DFF_X1 port map( D => n9890, CK => clk, Q => 
                           registers_19_28_port, QN => n15857);
   registers_reg_20_28_inst : DFF_X1 port map( D => n9889, CK => clk, Q => 
                           net271562, QN => n14829);
   registers_reg_21_28_inst : DFF_X1 port map( D => n9888, CK => clk, Q => 
                           net271561, QN => n12203);
   registers_reg_22_28_inst : DFF_X1 port map( D => n9887, CK => clk, Q => 
                           registers_22_28_port, QN => n15400);
   registers_reg_23_28_inst : DFF_X1 port map( D => n9886, CK => clk, Q => 
                           registers_23_28_port, QN => n15910);
   registers_reg_24_28_inst : DFF_X1 port map( D => n9885, CK => clk, Q => 
                           net227413, QN => n15207);
   registers_reg_25_28_inst : DFF_X1 port map( D => n9884, CK => clk, Q => 
                           registers_25_28_port, QN => n14326);
   registers_reg_26_28_inst : DFF_X1 port map( D => n9883, CK => clk, Q => 
                           net271560, QN => n12353);
   registers_reg_27_28_inst : DFF_X1 port map( D => n9882, CK => clk, Q => 
                           net271559, QN => n12045);
   registers_reg_28_28_inst : DFF_X1 port map( D => n9881, CK => clk, Q => 
                           net227412, QN => n15030);
   registers_reg_29_28_inst : DFF_X1 port map( D => n9880, CK => clk, Q => 
                           registers_29_28_port, QN => n15848);
   registers_reg_30_28_inst : DFF_X1 port map( D => n9879, CK => clk, Q => 
                           registers_30_28_port, QN => n14676);
   registers_reg_31_28_inst : DFF_X1 port map( D => n9878, CK => clk, Q => 
                           net227411, QN => n15732);
   registers_reg_32_28_inst : DFF_X1 port map( D => n9877, CK => clk, Q => 
                           net271558, QN => n12337);
   registers_reg_33_28_inst : DFF_X1 port map( D => n9876, CK => clk, Q => 
                           net271557, QN => n11873);
   registers_reg_34_28_inst : DFF_X1 port map( D => n9875, CK => clk, Q => 
                           registers_34_28_port, QN => n15493);
   registers_reg_35_28_inst : DFF_X1 port map( D => n9874, CK => clk, Q => 
                           net227410, QN => n15625);
   registers_reg_36_28_inst : DFF_X1 port map( D => n9873, CK => clk, Q => 
                           registers_36_28_port, QN => n15180);
   registers_reg_37_28_inst : DFF_X1 port map( D => n9872, CK => clk, Q => 
                           registers_37_28_port, QN => n14407);
   registers_reg_38_28_inst : DFF_X1 port map( D => n9871, CK => clk, Q => 
                           registers_38_28_port, QN => n15064);
   registers_reg_39_28_inst : DFF_X1 port map( D => n9870, CK => clk, Q => 
                           net271556, QN => n12169);
   registers_reg_40_28_inst : DFF_X1 port map( D => n9869, CK => clk, Q => 
                           registers_40_28_port, QN => n15148);
   registers_reg_41_28_inst : DFF_X1 port map( D => n9868, CK => clk, Q => 
                           registers_41_28_port, QN => n14531);
   registers_reg_42_28_inst : DFF_X1 port map( D => n9867, CK => clk, Q => 
                           registers_42_28_port, QN => n15955);
   registers_reg_43_28_inst : DFF_X1 port map( D => n9866, CK => clk, Q => 
                           registers_43_28_port, QN => n14883);
   registers_reg_44_28_inst : DFF_X1 port map( D => n9865, CK => clk, Q => 
                           registers_44_28_port, QN => n15464);
   registers_reg_45_28_inst : DFF_X1 port map( D => n9864, CK => clk, Q => 
                           registers_45_28_port, QN => n14768);
   registers_reg_46_28_inst : DFF_X1 port map( D => n9863, CK => clk, Q => 
                           net227409, QN => n11948);
   registers_reg_47_28_inst : DFF_X1 port map( D => n9862, CK => clk, Q => 
                           registers_47_28_port, QN => n14544);
   registers_reg_48_28_inst : DFF_X1 port map( D => n9861, CK => clk, Q => 
                           registers_48_28_port, QN => n15549);
   registers_reg_49_28_inst : DFF_X1 port map( D => n9860, CK => clk, Q => 
                           registers_49_28_port, QN => n14475);
   registers_reg_50_28_inst : DFF_X1 port map( D => n9859, CK => clk, Q => 
                           registers_50_28_port, QN => n15997);
   registers_reg_51_28_inst : DFF_X1 port map( D => n9858, CK => clk, Q => 
                           registers_51_28_port, QN => n15425);
   registers_reg_52_28_inst : DFF_X1 port map( D => n9857, CK => clk, Q => 
                           net227408, QN => n14935);
   registers_reg_53_28_inst : DFF_X1 port map( D => n9856, CK => clk, Q => 
                           net227407, QN => n15946);
   registers_reg_54_28_inst : DFF_X1 port map( D => n9855, CK => clk, Q => 
                           registers_54_28_port, QN => n14596);
   registers_reg_55_28_inst : DFF_X1 port map( D => n9854, CK => clk, Q => 
                           registers_55_28_port, QN => n12158);
   registers_reg_56_28_inst : DFF_X1 port map( D => n9853, CK => clk, Q => 
                           registers_56_28_port, QN => n16011);
   registers_reg_57_28_inst : DFF_X1 port map( D => n9852, CK => clk, Q => 
                           net227406, QN => n15268);
   registers_reg_58_28_inst : DFF_X1 port map( D => n9851, CK => clk, Q => 
                           net227405, QN => n14884);
   registers_reg_59_28_inst : DFF_X1 port map( D => n9850, CK => clk, Q => 
                           registers_59_28_port, QN => n15430);
   registers_reg_60_28_inst : DFF_X1 port map( D => n9849, CK => clk, Q => 
                           registers_60_28_port, QN => n14668);
   registers_reg_61_28_inst : DFF_X1 port map( D => n9848, CK => clk, Q => 
                           net227404, QN => n15659);
   registers_reg_62_28_inst : DFF_X1 port map( D => n9847, CK => clk, Q => 
                           registers_62_28_port, QN => n15121);
   registers_reg_63_28_inst : DFF_X1 port map( D => n9846, CK => clk, Q => 
                           registers_63_28_port, QN => n14482);
   to_mem_reg_28_inst : DFF_X1 port map( D => n9845, CK => clk, Q => net271555,
                           QN => n7697);
   registers_reg_64_28_inst : DFF_X1 port map( D => n9844, CK => clk, Q => 
                           net227403, QN => n16147);
   registers_reg_65_28_inst : DFF_X1 port map( D => n9843, CK => clk, Q => 
                           net227402, QN => n16096);
   registers_reg_66_28_inst : DFF_X1 port map( D => n9842, CK => clk, Q => 
                           net227401, QN => n16058);
   registers_reg_67_28_inst : DFF_X1 port map( D => n9841, CK => clk, Q => 
                           net271554, QN => n14277);
   registers_reg_68_28_inst : DFF_X1 port map( D => n9840, CK => clk, Q => 
                           registers_68_28_port, QN => n16184);
   registers_reg_69_28_inst : DFF_X1 port map( D => n9839, CK => clk, Q => 
                           net227400, QN => n16136);
   registers_reg_70_28_inst : DFF_X1 port map( D => n9838, CK => clk, Q => 
                           net227399, QN => n16048);
   registers_reg_0_27_inst : DFF_X1 port map( D => n9837, CK => clk, Q => 
                           registers_0_27_port, QN => n15878);
   registers_reg_1_27_inst : DFF_X1 port map( D => n9836, CK => clk, Q => 
                           registers_1_27_port, QN => n15635);
   registers_reg_2_27_inst : DFF_X1 port map( D => n9835, CK => clk, Q => 
                           registers_2_27_port, QN => n14765);
   registers_reg_3_27_inst : DFF_X1 port map( D => n9834, CK => clk, Q => 
                           net227398, QN => n15731);
   registers_reg_4_27_inst : DFF_X1 port map( D => n9833, CK => clk, Q => 
                           registers_4_27_port, QN => n15455);
   registers_reg_5_27_inst : DFF_X1 port map( D => n9832, CK => clk, Q => 
                           registers_5_27_port, QN => n14705);
   registers_reg_6_27_inst : DFF_X1 port map( D => n9831, CK => clk, Q => 
                           net271553, QN => n12345);
   registers_reg_7_27_inst : DFF_X1 port map( D => n9830, CK => clk, Q => 
                           registers_7_27_port, QN => n15323);
   registers_reg_8_27_inst : DFF_X1 port map( D => n9829, CK => clk, Q => 
                           net227397, QN => n15236);
   registers_reg_9_27_inst : DFF_X1 port map( D => n9828, CK => clk, Q => 
                           registers_9_27_port, QN => n14355);
   registers_reg_10_27_inst : DFF_X1 port map( D => n9827, CK => clk, Q => 
                           registers_10_27_port, QN => n14706);
   registers_reg_11_27_inst : DFF_X1 port map( D => n9826, CK => clk, Q => 
                           registers_11_27_port, QN => n14422);
   registers_reg_12_27_inst : DFF_X1 port map( D => n9825, CK => clk, Q => 
                           registers_12_27_port, QN => n15666);
   registers_reg_13_27_inst : DFF_X1 port map( D => n9824, CK => clk, Q => 
                           net227396, QN => n15068);
   registers_reg_14_27_inst : DFF_X1 port map( D => n9823, CK => clk, Q => 
                           net271552, QN => n11878);
   registers_reg_15_27_inst : DFF_X1 port map( D => n9822, CK => clk, Q => 
                           registers_15_27_port, QN => n15289);
   registers_reg_16_27_inst : DFF_X1 port map( D => n9821, CK => clk, Q => 
                           registers_16_27_port, QN => n15696);
   registers_reg_17_27_inst : DFF_X1 port map( D => n9820, CK => clk, Q => 
                           registers_17_27_port, QN => n14602);
   registers_reg_18_27_inst : DFF_X1 port map( D => n9819, CK => clk, Q => 
                           registers_18_27_port, QN => n14417);
   registers_reg_19_27_inst : DFF_X1 port map( D => n9818, CK => clk, Q => 
                           registers_19_27_port, QN => n15856);
   registers_reg_20_27_inst : DFF_X1 port map( D => n9817, CK => clk, Q => 
                           net271551, QN => n14828);
   registers_reg_21_27_inst : DFF_X1 port map( D => n9816, CK => clk, Q => 
                           net271550, QN => n12202);
   registers_reg_22_27_inst : DFF_X1 port map( D => n9815, CK => clk, Q => 
                           registers_22_27_port, QN => n15399);
   registers_reg_23_27_inst : DFF_X1 port map( D => n9814, CK => clk, Q => 
                           registers_23_27_port, QN => n15909);
   registers_reg_24_27_inst : DFF_X1 port map( D => n9813, CK => clk, Q => 
                           net227395, QN => n15206);
   registers_reg_25_27_inst : DFF_X1 port map( D => n9812, CK => clk, Q => 
                           registers_25_27_port, QN => n14325);
   registers_reg_26_27_inst : DFF_X1 port map( D => n9811, CK => clk, Q => 
                           net271549, QN => n12352);
   registers_reg_27_27_inst : DFF_X1 port map( D => n9810, CK => clk, Q => 
                           net271548, QN => n12044);
   registers_reg_28_27_inst : DFF_X1 port map( D => n9809, CK => clk, Q => 
                           net227394, QN => n15029);
   registers_reg_29_27_inst : DFF_X1 port map( D => n9808, CK => clk, Q => 
                           registers_29_27_port, QN => n15847);
   registers_reg_30_27_inst : DFF_X1 port map( D => n9807, CK => clk, Q => 
                           registers_30_27_port, QN => n14675);
   registers_reg_31_27_inst : DFF_X1 port map( D => n9806, CK => clk, Q => 
                           net227393, QN => n15730);
   registers_reg_32_27_inst : DFF_X1 port map( D => n9805, CK => clk, Q => 
                           net271547, QN => n12336);
   registers_reg_33_27_inst : DFF_X1 port map( D => n9804, CK => clk, Q => 
                           net271546, QN => n11872);
   registers_reg_34_27_inst : DFF_X1 port map( D => n9803, CK => clk, Q => 
                           registers_34_27_port, QN => n15492);
   registers_reg_35_27_inst : DFF_X1 port map( D => n9802, CK => clk, Q => 
                           net227392, QN => n15624);
   registers_reg_36_27_inst : DFF_X1 port map( D => n9801, CK => clk, Q => 
                           registers_36_27_port, QN => n15179);
   registers_reg_37_27_inst : DFF_X1 port map( D => n9800, CK => clk, Q => 
                           registers_37_27_port, QN => n14406);
   registers_reg_38_27_inst : DFF_X1 port map( D => n9799, CK => clk, Q => 
                           registers_38_27_port, QN => n15063);
   registers_reg_39_27_inst : DFF_X1 port map( D => n9798, CK => clk, Q => 
                           net271545, QN => n12168);
   registers_reg_40_27_inst : DFF_X1 port map( D => n9797, CK => clk, Q => 
                           registers_40_27_port, QN => n15147);
   registers_reg_41_27_inst : DFF_X1 port map( D => n9796, CK => clk, Q => 
                           registers_41_27_port, QN => n14530);
   registers_reg_42_27_inst : DFF_X1 port map( D => n9795, CK => clk, Q => 
                           registers_42_27_port, QN => n15954);
   registers_reg_43_27_inst : DFF_X1 port map( D => n9794, CK => clk, Q => 
                           registers_43_27_port, QN => n14881);
   registers_reg_44_27_inst : DFF_X1 port map( D => n9793, CK => clk, Q => 
                           registers_44_27_port, QN => n15463);
   registers_reg_45_27_inst : DFF_X1 port map( D => n9792, CK => clk, Q => 
                           registers_45_27_port, QN => n14766);
   registers_reg_46_27_inst : DFF_X1 port map( D => n9791, CK => clk, Q => 
                           net227391, QN => n11947);
   registers_reg_47_27_inst : DFF_X1 port map( D => n9790, CK => clk, Q => 
                           registers_47_27_port, QN => n14543);
   registers_reg_48_27_inst : DFF_X1 port map( D => n9789, CK => clk, Q => 
                           registers_48_27_port, QN => n15548);
   registers_reg_49_27_inst : DFF_X1 port map( D => n9788, CK => clk, Q => 
                           registers_49_27_port, QN => n14474);
   registers_reg_50_27_inst : DFF_X1 port map( D => n9787, CK => clk, Q => 
                           registers_50_27_port, QN => n15996);
   registers_reg_51_27_inst : DFF_X1 port map( D => n9786, CK => clk, Q => 
                           registers_51_27_port, QN => n15424);
   registers_reg_52_27_inst : DFF_X1 port map( D => n9785, CK => clk, Q => 
                           net227390, QN => n14934);
   registers_reg_53_27_inst : DFF_X1 port map( D => n9784, CK => clk, Q => 
                           net227389, QN => n15945);
   registers_reg_54_27_inst : DFF_X1 port map( D => n9783, CK => clk, Q => 
                           registers_54_27_port, QN => n14595);
   registers_reg_55_27_inst : DFF_X1 port map( D => n9782, CK => clk, Q => 
                           registers_55_27_port, QN => n12157);
   registers_reg_56_27_inst : DFF_X1 port map( D => n9781, CK => clk, Q => 
                           registers_56_27_port, QN => n16010);
   registers_reg_57_27_inst : DFF_X1 port map( D => n9780, CK => clk, Q => 
                           net227388, QN => n15267);
   registers_reg_58_27_inst : DFF_X1 port map( D => n9779, CK => clk, Q => 
                           net227387, QN => n14882);
   registers_reg_59_27_inst : DFF_X1 port map( D => n9778, CK => clk, Q => 
                           registers_59_27_port, QN => n15429);
   registers_reg_60_27_inst : DFF_X1 port map( D => n9777, CK => clk, Q => 
                           registers_60_27_port, QN => n14667);
   registers_reg_61_27_inst : DFF_X1 port map( D => n9776, CK => clk, Q => 
                           net227386, QN => n15658);
   registers_reg_62_27_inst : DFF_X1 port map( D => n9775, CK => clk, Q => 
                           registers_62_27_port, QN => n15120);
   registers_reg_63_27_inst : DFF_X1 port map( D => n9774, CK => clk, Q => 
                           registers_63_27_port, QN => n14481);
   to_mem_reg_27_inst : DFF_X1 port map( D => n9773, CK => clk, Q => net271544,
                           QN => n7698);
   registers_reg_64_27_inst : DFF_X1 port map( D => n9772, CK => clk, Q => 
                           net227385, QN => n16146);
   registers_reg_65_27_inst : DFF_X1 port map( D => n9771, CK => clk, Q => 
                           net227384, QN => n16095);
   registers_reg_66_27_inst : DFF_X1 port map( D => n9770, CK => clk, Q => 
                           net227383, QN => n16057);
   registers_reg_67_27_inst : DFF_X1 port map( D => n9769, CK => clk, Q => 
                           net271543, QN => n14276);
   registers_reg_68_27_inst : DFF_X1 port map( D => n9768, CK => clk, Q => 
                           registers_68_27_port, QN => n16183);
   registers_reg_69_27_inst : DFF_X1 port map( D => n9767, CK => clk, Q => 
                           net227382, QN => n16135);
   registers_reg_70_27_inst : DFF_X1 port map( D => n9766, CK => clk, Q => 
                           net227381, QN => n16047);
   registers_reg_0_26_inst : DFF_X1 port map( D => n9765, CK => clk, Q => 
                           registers_0_26_port, QN => n15877);
   registers_reg_1_26_inst : DFF_X1 port map( D => n9764, CK => clk, Q => 
                           registers_1_26_port, QN => n15634);
   registers_reg_2_26_inst : DFF_X1 port map( D => n9763, CK => clk, Q => 
                           registers_2_26_port, QN => n14763);
   registers_reg_3_26_inst : DFF_X1 port map( D => n9762, CK => clk, Q => 
                           net227380, QN => n15729);
   registers_reg_4_26_inst : DFF_X1 port map( D => n9761, CK => clk, Q => 
                           registers_4_26_port, QN => n15454);
   registers_reg_5_26_inst : DFF_X1 port map( D => n9760, CK => clk, Q => 
                           registers_5_26_port, QN => n14703);
   registers_reg_6_26_inst : DFF_X1 port map( D => n9759, CK => clk, Q => 
                           net271542, QN => n12344);
   registers_reg_7_26_inst : DFF_X1 port map( D => n9758, CK => clk, Q => 
                           registers_7_26_port, QN => n15322);
   registers_reg_8_26_inst : DFF_X1 port map( D => n9757, CK => clk, Q => 
                           net227379, QN => n15235);
   registers_reg_9_26_inst : DFF_X1 port map( D => n9756, CK => clk, Q => 
                           registers_9_26_port, QN => n14354);
   registers_reg_10_26_inst : DFF_X1 port map( D => n9755, CK => clk, Q => 
                           registers_10_26_port, QN => n14704);
   registers_reg_11_26_inst : DFF_X1 port map( D => n9754, CK => clk, Q => 
                           registers_11_26_port, QN => n14421);
   registers_reg_12_26_inst : DFF_X1 port map( D => n9753, CK => clk, Q => 
                           registers_12_26_port, QN => n15665);
   registers_reg_13_26_inst : DFF_X1 port map( D => n9752, CK => clk, Q => 
                           net227378, QN => n15067);
   registers_reg_14_26_inst : DFF_X1 port map( D => n9751, CK => clk, Q => 
                           net271541, QN => n11877);
   registers_reg_15_26_inst : DFF_X1 port map( D => n9750, CK => clk, Q => 
                           registers_15_26_port, QN => n15288);
   registers_reg_16_26_inst : DFF_X1 port map( D => n9749, CK => clk, Q => 
                           registers_16_26_port, QN => n15695);
   registers_reg_17_26_inst : DFF_X1 port map( D => n9748, CK => clk, Q => 
                           registers_17_26_port, QN => n14601);
   registers_reg_18_26_inst : DFF_X1 port map( D => n9747, CK => clk, Q => 
                           registers_18_26_port, QN => n14416);
   registers_reg_19_26_inst : DFF_X1 port map( D => n9746, CK => clk, Q => 
                           registers_19_26_port, QN => n15855);
   registers_reg_20_26_inst : DFF_X1 port map( D => n9745, CK => clk, Q => 
                           net271540, QN => n14827);
   registers_reg_21_26_inst : DFF_X1 port map( D => n9744, CK => clk, Q => 
                           net271539, QN => n12201);
   registers_reg_22_26_inst : DFF_X1 port map( D => n9743, CK => clk, Q => 
                           registers_22_26_port, QN => n15398);
   registers_reg_23_26_inst : DFF_X1 port map( D => n9742, CK => clk, Q => 
                           registers_23_26_port, QN => n15908);
   registers_reg_24_26_inst : DFF_X1 port map( D => n9741, CK => clk, Q => 
                           net227377, QN => n15205);
   registers_reg_25_26_inst : DFF_X1 port map( D => n9740, CK => clk, Q => 
                           registers_25_26_port, QN => n14324);
   registers_reg_26_26_inst : DFF_X1 port map( D => n9739, CK => clk, Q => 
                           net271538, QN => n12351);
   registers_reg_27_26_inst : DFF_X1 port map( D => n9738, CK => clk, Q => 
                           net271537, QN => n12043);
   registers_reg_28_26_inst : DFF_X1 port map( D => n9737, CK => clk, Q => 
                           net227376, QN => n15028);
   registers_reg_29_26_inst : DFF_X1 port map( D => n9736, CK => clk, Q => 
                           registers_29_26_port, QN => n15846);
   registers_reg_30_26_inst : DFF_X1 port map( D => n9735, CK => clk, Q => 
                           registers_30_26_port, QN => n14674);
   registers_reg_31_26_inst : DFF_X1 port map( D => n9734, CK => clk, Q => 
                           net227375, QN => n15728);
   registers_reg_32_26_inst : DFF_X1 port map( D => n9733, CK => clk, Q => 
                           net271536, QN => n12335);
   registers_reg_33_26_inst : DFF_X1 port map( D => n9732, CK => clk, Q => 
                           net271535, QN => n11871);
   registers_reg_34_26_inst : DFF_X1 port map( D => n9731, CK => clk, Q => 
                           registers_34_26_port, QN => n15491);
   registers_reg_35_26_inst : DFF_X1 port map( D => n9730, CK => clk, Q => 
                           net227374, QN => n15623);
   registers_reg_36_26_inst : DFF_X1 port map( D => n9729, CK => clk, Q => 
                           registers_36_26_port, QN => n15178);
   registers_reg_37_26_inst : DFF_X1 port map( D => n9728, CK => clk, Q => 
                           registers_37_26_port, QN => n14405);
   registers_reg_38_26_inst : DFF_X1 port map( D => n9727, CK => clk, Q => 
                           registers_38_26_port, QN => n15062);
   registers_reg_39_26_inst : DFF_X1 port map( D => n9726, CK => clk, Q => 
                           net271534, QN => n12167);
   registers_reg_40_26_inst : DFF_X1 port map( D => n9725, CK => clk, Q => 
                           registers_40_26_port, QN => n15146);
   registers_reg_41_26_inst : DFF_X1 port map( D => n9724, CK => clk, Q => 
                           registers_41_26_port, QN => n14529);
   registers_reg_42_26_inst : DFF_X1 port map( D => n9723, CK => clk, Q => 
                           registers_42_26_port, QN => n15953);
   registers_reg_43_26_inst : DFF_X1 port map( D => n9722, CK => clk, Q => 
                           registers_43_26_port, QN => n14879);
   registers_reg_44_26_inst : DFF_X1 port map( D => n9721, CK => clk, Q => 
                           registers_44_26_port, QN => n15462);
   registers_reg_45_26_inst : DFF_X1 port map( D => n9720, CK => clk, Q => 
                           registers_45_26_port, QN => n14764);
   registers_reg_46_26_inst : DFF_X1 port map( D => n9719, CK => clk, Q => 
                           net227373, QN => n11946);
   registers_reg_47_26_inst : DFF_X1 port map( D => n9718, CK => clk, Q => 
                           registers_47_26_port, QN => n14542);
   registers_reg_48_26_inst : DFF_X1 port map( D => n9717, CK => clk, Q => 
                           registers_48_26_port, QN => n15547);
   registers_reg_49_26_inst : DFF_X1 port map( D => n9716, CK => clk, Q => 
                           registers_49_26_port, QN => n14473);
   registers_reg_50_26_inst : DFF_X1 port map( D => n9715, CK => clk, Q => 
                           registers_50_26_port, QN => n15995);
   registers_reg_51_26_inst : DFF_X1 port map( D => n9714, CK => clk, Q => 
                           registers_51_26_port, QN => n15423);
   registers_reg_52_26_inst : DFF_X1 port map( D => n9713, CK => clk, Q => 
                           net227372, QN => n14933);
   registers_reg_53_26_inst : DFF_X1 port map( D => n9712, CK => clk, Q => 
                           net227371, QN => n15944);
   registers_reg_54_26_inst : DFF_X1 port map( D => n9711, CK => clk, Q => 
                           registers_54_26_port, QN => n14594);
   registers_reg_55_26_inst : DFF_X1 port map( D => n9710, CK => clk, Q => 
                           registers_55_26_port, QN => n12156);
   registers_reg_56_26_inst : DFF_X1 port map( D => n9709, CK => clk, Q => 
                           registers_56_26_port, QN => n16009);
   registers_reg_57_26_inst : DFF_X1 port map( D => n9708, CK => clk, Q => 
                           net227370, QN => n15266);
   registers_reg_58_26_inst : DFF_X1 port map( D => n9707, CK => clk, Q => 
                           net227369, QN => n14880);
   registers_reg_59_26_inst : DFF_X1 port map( D => n9706, CK => clk, Q => 
                           registers_59_26_port, QN => n15428);
   registers_reg_60_26_inst : DFF_X1 port map( D => n9705, CK => clk, Q => 
                           registers_60_26_port, QN => n14666);
   registers_reg_61_26_inst : DFF_X1 port map( D => n9704, CK => clk, Q => 
                           net227368, QN => n15657);
   registers_reg_62_26_inst : DFF_X1 port map( D => n9703, CK => clk, Q => 
                           registers_62_26_port, QN => n15119);
   registers_reg_63_26_inst : DFF_X1 port map( D => n9702, CK => clk, Q => 
                           registers_63_26_port, QN => n14480);
   to_mem_reg_26_inst : DFF_X1 port map( D => n9701, CK => clk, Q => net271533,
                           QN => n7699);
   registers_reg_64_26_inst : DFF_X1 port map( D => n9700, CK => clk, Q => 
                           net227367, QN => n16145);
   registers_reg_65_26_inst : DFF_X1 port map( D => n9699, CK => clk, Q => 
                           net227366, QN => n16094);
   registers_reg_66_26_inst : DFF_X1 port map( D => n9698, CK => clk, Q => 
                           net227365, QN => n16056);
   registers_reg_67_26_inst : DFF_X1 port map( D => n9697, CK => clk, Q => 
                           net271532, QN => n14275);
   registers_reg_68_26_inst : DFF_X1 port map( D => n9696, CK => clk, Q => 
                           registers_68_26_port, QN => n16182);
   registers_reg_69_26_inst : DFF_X1 port map( D => n9695, CK => clk, Q => 
                           net227364, QN => n16134);
   registers_reg_70_26_inst : DFF_X1 port map( D => n9694, CK => clk, Q => 
                           net227363, QN => n16046);
   registers_reg_0_25_inst : DFF_X1 port map( D => n9693, CK => clk, Q => 
                           registers_0_25_port, QN => n15876);
   registers_reg_1_25_inst : DFF_X1 port map( D => n9692, CK => clk, Q => 
                           registers_1_25_port, QN => n15633);
   registers_reg_2_25_inst : DFF_X1 port map( D => n9691, CK => clk, Q => 
                           registers_2_25_port, QN => n14761);
   registers_reg_3_25_inst : DFF_X1 port map( D => n9690, CK => clk, Q => 
                           net227362, QN => n15727);
   registers_reg_4_25_inst : DFF_X1 port map( D => n9689, CK => clk, Q => 
                           registers_4_25_port, QN => n15453);
   registers_reg_5_25_inst : DFF_X1 port map( D => n9688, CK => clk, Q => 
                           registers_5_25_port, QN => n14819);
   registers_reg_6_25_inst : DFF_X1 port map( D => n9687, CK => clk, Q => 
                           net271531, QN => n12343);
   registers_reg_7_25_inst : DFF_X1 port map( D => n9686, CK => clk, Q => 
                           registers_7_25_port, QN => n15321);
   registers_reg_8_25_inst : DFF_X1 port map( D => n9685, CK => clk, Q => 
                           net227361, QN => n15234);
   registers_reg_9_25_inst : DFF_X1 port map( D => n9684, CK => clk, Q => 
                           registers_9_25_port, QN => n14353);
   registers_reg_10_25_inst : DFF_X1 port map( D => n9683, CK => clk, Q => 
                           registers_10_25_port, QN => n14702);
   registers_reg_11_25_inst : DFF_X1 port map( D => n9682, CK => clk, Q => 
                           registers_11_25_port, QN => n14420);
   registers_reg_12_25_inst : DFF_X1 port map( D => n9681, CK => clk, Q => 
                           registers_12_25_port, QN => n15664);
   registers_reg_13_25_inst : DFF_X1 port map( D => n9680, CK => clk, Q => 
                           net227360, QN => n15066);
   registers_reg_14_25_inst : DFF_X1 port map( D => n9679, CK => clk, Q => 
                           net271530, QN => n11876);
   registers_reg_15_25_inst : DFF_X1 port map( D => n9678, CK => clk, Q => 
                           registers_15_25_port, QN => n15287);
   registers_reg_16_25_inst : DFF_X1 port map( D => n9677, CK => clk, Q => 
                           registers_16_25_port, QN => n15694);
   registers_reg_17_25_inst : DFF_X1 port map( D => n9676, CK => clk, Q => 
                           registers_17_25_port, QN => n14600);
   registers_reg_18_25_inst : DFF_X1 port map( D => n9675, CK => clk, Q => 
                           registers_18_25_port, QN => n14415);
   registers_reg_19_25_inst : DFF_X1 port map( D => n9674, CK => clk, Q => 
                           registers_19_25_port, QN => n15854);
   registers_reg_20_25_inst : DFF_X1 port map( D => n9673, CK => clk, Q => 
                           net271529, QN => n14826);
   registers_reg_21_25_inst : DFF_X1 port map( D => n9672, CK => clk, Q => 
                           net271528, QN => n12200);
   registers_reg_22_25_inst : DFF_X1 port map( D => n9671, CK => clk, Q => 
                           registers_22_25_port, QN => n15397);
   registers_reg_23_25_inst : DFF_X1 port map( D => n9670, CK => clk, Q => 
                           registers_23_25_port, QN => n15907);
   registers_reg_24_25_inst : DFF_X1 port map( D => n9669, CK => clk, Q => 
                           net227359, QN => n15204);
   registers_reg_25_25_inst : DFF_X1 port map( D => n9668, CK => clk, Q => 
                           registers_25_25_port, QN => n14323);
   registers_reg_26_25_inst : DFF_X1 port map( D => n9667, CK => clk, Q => 
                           net271527, QN => n12350);
   registers_reg_27_25_inst : DFF_X1 port map( D => n9666, CK => clk, Q => 
                           net271526, QN => n12042);
   registers_reg_28_25_inst : DFF_X1 port map( D => n9665, CK => clk, Q => 
                           net227358, QN => n15027);
   registers_reg_29_25_inst : DFF_X1 port map( D => n9664, CK => clk, Q => 
                           registers_29_25_port, QN => n15845);
   registers_reg_30_25_inst : DFF_X1 port map( D => n9663, CK => clk, Q => 
                           registers_30_25_port, QN => n14673);
   registers_reg_31_25_inst : DFF_X1 port map( D => n9662, CK => clk, Q => 
                           net227357, QN => n15726);
   registers_reg_32_25_inst : DFF_X1 port map( D => n9661, CK => clk, Q => 
                           net271525, QN => n12334);
   registers_reg_33_25_inst : DFF_X1 port map( D => n9660, CK => clk, Q => 
                           net271524, QN => n11870);
   registers_reg_34_25_inst : DFF_X1 port map( D => n9659, CK => clk, Q => 
                           registers_34_25_port, QN => n15490);
   registers_reg_35_25_inst : DFF_X1 port map( D => n9658, CK => clk, Q => 
                           net227356, QN => n15622);
   registers_reg_36_25_inst : DFF_X1 port map( D => n9657, CK => clk, Q => 
                           registers_36_25_port, QN => n15177);
   registers_reg_37_25_inst : DFF_X1 port map( D => n9656, CK => clk, Q => 
                           registers_37_25_port, QN => n14404);
   registers_reg_38_25_inst : DFF_X1 port map( D => n9655, CK => clk, Q => 
                           registers_38_25_port, QN => n15061);
   registers_reg_39_25_inst : DFF_X1 port map( D => n9654, CK => clk, Q => 
                           net271523, QN => n12166);
   registers_reg_40_25_inst : DFF_X1 port map( D => n9653, CK => clk, Q => 
                           registers_40_25_port, QN => n15145);
   registers_reg_41_25_inst : DFF_X1 port map( D => n9652, CK => clk, Q => 
                           registers_41_25_port, QN => n14528);
   registers_reg_42_25_inst : DFF_X1 port map( D => n9651, CK => clk, Q => 
                           registers_42_25_port, QN => n15952);
   registers_reg_43_25_inst : DFF_X1 port map( D => n9650, CK => clk, Q => 
                           registers_43_25_port, QN => n14877);
   registers_reg_44_25_inst : DFF_X1 port map( D => n9649, CK => clk, Q => 
                           registers_44_25_port, QN => n15461);
   registers_reg_45_25_inst : DFF_X1 port map( D => n9648, CK => clk, Q => 
                           registers_45_25_port, QN => n14762);
   registers_reg_46_25_inst : DFF_X1 port map( D => n9647, CK => clk, Q => 
                           net227355, QN => n11945);
   registers_reg_47_25_inst : DFF_X1 port map( D => n9646, CK => clk, Q => 
                           registers_47_25_port, QN => n14541);
   registers_reg_48_25_inst : DFF_X1 port map( D => n9645, CK => clk, Q => 
                           registers_48_25_port, QN => n15546);
   registers_reg_49_25_inst : DFF_X1 port map( D => n9644, CK => clk, Q => 
                           registers_49_25_port, QN => n14472);
   registers_reg_50_25_inst : DFF_X1 port map( D => n9643, CK => clk, Q => 
                           registers_50_25_port, QN => n15994);
   registers_reg_51_25_inst : DFF_X1 port map( D => n9642, CK => clk, Q => 
                           registers_51_25_port, QN => n15422);
   registers_reg_52_25_inst : DFF_X1 port map( D => n9641_port, CK => clk, Q =>
                           net227354, QN => n14932);
   registers_reg_53_25_inst : DFF_X1 port map( D => n9640, CK => clk, Q => 
                           net227353, QN => n15943);
   registers_reg_54_25_inst : DFF_X1 port map( D => n9639, CK => clk, Q => 
                           registers_54_25_port, QN => n14593);
   registers_reg_55_25_inst : DFF_X1 port map( D => n9638, CK => clk, Q => 
                           registers_55_25_port, QN => n12155);
   registers_reg_56_25_inst : DFF_X1 port map( D => n9637, CK => clk, Q => 
                           registers_56_25_port, QN => n16008);
   registers_reg_57_25_inst : DFF_X1 port map( D => n9636, CK => clk, Q => 
                           net227352, QN => n15265);
   registers_reg_58_25_inst : DFF_X1 port map( D => n9635, CK => clk, Q => 
                           net227351, QN => n14878);
   registers_reg_59_25_inst : DFF_X1 port map( D => n9634, CK => clk, Q => 
                           registers_59_25_port, QN => n15520);
   registers_reg_60_25_inst : DFF_X1 port map( D => n9633, CK => clk, Q => 
                           registers_60_25_port, QN => n14665);
   registers_reg_61_25_inst : DFF_X1 port map( D => n9632, CK => clk, Q => 
                           net227350, QN => n15656);
   registers_reg_62_25_inst : DFF_X1 port map( D => n9631, CK => clk, Q => 
                           registers_62_25_port, QN => n15118);
   registers_reg_63_25_inst : DFF_X1 port map( D => n9630, CK => clk, Q => 
                           registers_63_25_port, QN => n14479);
   to_mem_reg_25_inst : DFF_X1 port map( D => n9629, CK => clk, Q => net271522,
                           QN => n7700);
   registers_reg_64_25_inst : DFF_X1 port map( D => n9628, CK => clk, Q => 
                           net227349, QN => n16144);
   registers_reg_65_25_inst : DFF_X1 port map( D => n9627, CK => clk, Q => 
                           net227348, QN => n16093);
   registers_reg_66_25_inst : DFF_X1 port map( D => n9626, CK => clk, Q => 
                           net227347, QN => n16055);
   registers_reg_67_25_inst : DFF_X1 port map( D => n9625, CK => clk, Q => 
                           net271521, QN => n14274);
   registers_reg_68_25_inst : DFF_X1 port map( D => n9624, CK => clk, Q => 
                           registers_68_25_port, QN => n16181);
   registers_reg_69_25_inst : DFF_X1 port map( D => n9623, CK => clk, Q => 
                           net227346, QN => n16133);
   registers_reg_70_25_inst : DFF_X1 port map( D => n9622, CK => clk, Q => 
                           net227345, QN => n16045);
   registers_reg_0_24_inst : DFF_X1 port map( D => n9621, CK => clk, Q => 
                           registers_0_24_port, QN => n15875);
   registers_reg_1_24_inst : DFF_X1 port map( D => n9620, CK => clk, Q => 
                           registers_1_24_port, QN => n15632);
   registers_reg_2_24_inst : DFF_X1 port map( D => n9619, CK => clk, Q => 
                           registers_2_24_port, QN => n14759);
   registers_reg_3_24_inst : DFF_X1 port map( D => n9618, CK => clk, Q => 
                           net227344, QN => n15725);
   registers_reg_4_24_inst : DFF_X1 port map( D => n9617, CK => clk, Q => 
                           registers_4_24_port, QN => n15452);
   registers_reg_5_24_inst : DFF_X1 port map( D => n9616, CK => clk, Q => 
                           registers_5_24_port, QN => n14818);
   registers_reg_6_24_inst : DFF_X1 port map( D => n9615, CK => clk, Q => 
                           net271520, QN => n12342);
   registers_reg_7_24_inst : DFF_X1 port map( D => n9614, CK => clk, Q => 
                           registers_7_24_port, QN => n15320);
   registers_reg_8_24_inst : DFF_X1 port map( D => n9613, CK => clk, Q => 
                           net227343, QN => n15233);
   registers_reg_9_24_inst : DFF_X1 port map( D => n9612, CK => clk, Q => 
                           registers_9_24_port, QN => n14352);
   registers_reg_10_24_inst : DFF_X1 port map( D => n9611, CK => clk, Q => 
                           registers_10_24_port, QN => n14701);
   registers_reg_11_24_inst : DFF_X1 port map( D => n9610, CK => clk, Q => 
                           registers_11_24_port, QN => n14419);
   registers_reg_12_24_inst : DFF_X1 port map( D => n9609, CK => clk, Q => 
                           registers_12_24_port, QN => n15663);
   registers_reg_13_24_inst : DFF_X1 port map( D => n9608, CK => clk, Q => 
                           net227342, QN => n15065);
   registers_reg_14_24_inst : DFF_X1 port map( D => n9607, CK => clk, Q => 
                           net271519, QN => n11875);
   registers_reg_15_24_inst : DFF_X1 port map( D => n9606, CK => clk, Q => 
                           registers_15_24_port, QN => n15286);
   registers_reg_16_24_inst : DFF_X1 port map( D => n9605, CK => clk, Q => 
                           registers_16_24_port, QN => n15693);
   registers_reg_17_24_inst : DFF_X1 port map( D => n9604, CK => clk, Q => 
                           registers_17_24_port, QN => n14599);
   registers_reg_18_24_inst : DFF_X1 port map( D => n9603, CK => clk, Q => 
                           registers_18_24_port, QN => n14414);
   registers_reg_19_24_inst : DFF_X1 port map( D => n9602, CK => clk, Q => 
                           registers_19_24_port, QN => n15853);
   registers_reg_20_24_inst : DFF_X1 port map( D => n9601, CK => clk, Q => 
                           net271518, QN => n14825);
   registers_reg_21_24_inst : DFF_X1 port map( D => n9600, CK => clk, Q => 
                           net271517, QN => n12199);
   registers_reg_22_24_inst : DFF_X1 port map( D => n9599, CK => clk, Q => 
                           registers_22_24_port, QN => n15396);
   registers_reg_23_24_inst : DFF_X1 port map( D => n9598, CK => clk, Q => 
                           registers_23_24_port, QN => n15906);
   registers_reg_24_24_inst : DFF_X1 port map( D => n9597, CK => clk, Q => 
                           net227341, QN => n15203);
   registers_reg_25_24_inst : DFF_X1 port map( D => n9596, CK => clk, Q => 
                           registers_25_24_port, QN => n14322);
   registers_reg_26_24_inst : DFF_X1 port map( D => n9595, CK => clk, Q => 
                           net271516, QN => n12349);
   registers_reg_27_24_inst : DFF_X1 port map( D => n9594, CK => clk, Q => 
                           net271515, QN => n12041);
   registers_reg_28_24_inst : DFF_X1 port map( D => n9593, CK => clk, Q => 
                           net227340, QN => n15026);
   registers_reg_29_24_inst : DFF_X1 port map( D => n9592, CK => clk, Q => 
                           registers_29_24_port, QN => n15844);
   registers_reg_30_24_inst : DFF_X1 port map( D => n9591, CK => clk, Q => 
                           registers_30_24_port, QN => n14672);
   registers_reg_31_24_inst : DFF_X1 port map( D => n9590, CK => clk, Q => 
                           net227339, QN => n15724);
   registers_reg_32_24_inst : DFF_X1 port map( D => n9589, CK => clk, Q => 
                           net271514, QN => n12333);
   registers_reg_33_24_inst : DFF_X1 port map( D => n9588, CK => clk, Q => 
                           net271513, QN => n11869);
   registers_reg_34_24_inst : DFF_X1 port map( D => n9587, CK => clk, Q => 
                           registers_34_24_port, QN => n15489);
   registers_reg_35_24_inst : DFF_X1 port map( D => n9586, CK => clk, Q => 
                           net227338, QN => n15621);
   registers_reg_36_24_inst : DFF_X1 port map( D => n9585, CK => clk, Q => 
                           registers_36_24_port, QN => n15176);
   registers_reg_37_24_inst : DFF_X1 port map( D => n9584, CK => clk, Q => 
                           registers_37_24_port, QN => n14403);
   registers_reg_38_24_inst : DFF_X1 port map( D => n9583, CK => clk, Q => 
                           registers_38_24_port, QN => n15060);
   registers_reg_39_24_inst : DFF_X1 port map( D => n9582, CK => clk, Q => 
                           net271512, QN => n12165);
   registers_reg_40_24_inst : DFF_X1 port map( D => n9581, CK => clk, Q => 
                           registers_40_24_port, QN => n15144);
   registers_reg_41_24_inst : DFF_X1 port map( D => n9580, CK => clk, Q => 
                           registers_41_24_port, QN => n14527);
   registers_reg_42_24_inst : DFF_X1 port map( D => n9579, CK => clk, Q => 
                           registers_42_24_port, QN => n15951);
   registers_reg_43_24_inst : DFF_X1 port map( D => n9578, CK => clk, Q => 
                           registers_43_24_port, QN => n14875);
   registers_reg_44_24_inst : DFF_X1 port map( D => n9577, CK => clk, Q => 
                           registers_44_24_port, QN => n15460);
   registers_reg_45_24_inst : DFF_X1 port map( D => n9576, CK => clk, Q => 
                           registers_45_24_port, QN => n14760);
   registers_reg_46_24_inst : DFF_X1 port map( D => n9575, CK => clk, Q => 
                           net227337, QN => n11907);
   registers_reg_47_24_inst : DFF_X1 port map( D => n9574, CK => clk, Q => 
                           registers_47_24_port, QN => n14540);
   registers_reg_48_24_inst : DFF_X1 port map( D => n9573, CK => clk, Q => 
                           registers_48_24_port, QN => n15545);
   registers_reg_49_24_inst : DFF_X1 port map( D => n9572, CK => clk, Q => 
                           registers_49_24_port, QN => n14471);
   registers_reg_50_24_inst : DFF_X1 port map( D => n9571, CK => clk, Q => 
                           registers_50_24_port, QN => n15993);
   registers_reg_51_24_inst : DFF_X1 port map( D => n9570, CK => clk, Q => 
                           registers_51_24_port, QN => n15421);
   registers_reg_52_24_inst : DFF_X1 port map( D => n9569, CK => clk, Q => 
                           net227336, QN => n14931);
   registers_reg_53_24_inst : DFF_X1 port map( D => n9568, CK => clk, Q => 
                           net227335, QN => n15942);
   registers_reg_54_24_inst : DFF_X1 port map( D => n9567, CK => clk, Q => 
                           registers_54_24_port, QN => n14592);
   registers_reg_55_24_inst : DFF_X1 port map( D => n9566, CK => clk, Q => 
                           registers_55_24_port, QN => n12154);
   registers_reg_56_24_inst : DFF_X1 port map( D => n9565, CK => clk, Q => 
                           registers_56_24_port, QN => n16007);
   registers_reg_57_24_inst : DFF_X1 port map( D => n9564, CK => clk, Q => 
                           net227334, QN => n15264);
   registers_reg_58_24_inst : DFF_X1 port map( D => n9563, CK => clk, Q => 
                           net227333, QN => n14876);
   registers_reg_59_24_inst : DFF_X1 port map( D => n9562, CK => clk, Q => 
                           registers_59_24_port, QN => n15519);
   registers_reg_60_24_inst : DFF_X1 port map( D => n9561, CK => clk, Q => 
                           registers_60_24_port, QN => n14664);
   registers_reg_61_24_inst : DFF_X1 port map( D => n9560, CK => clk, Q => 
                           net227332, QN => n15655);
   registers_reg_62_24_inst : DFF_X1 port map( D => n9559, CK => clk, Q => 
                           registers_62_24_port, QN => n15117);
   registers_reg_63_24_inst : DFF_X1 port map( D => n9558, CK => clk, Q => 
                           registers_63_24_port, QN => n14478);
   to_mem_reg_24_inst : DFF_X1 port map( D => n9557, CK => clk, Q => net271511,
                           QN => n7701);
   registers_reg_64_24_inst : DFF_X1 port map( D => n9556, CK => clk, Q => 
                           net227331, QN => n16143);
   registers_reg_65_24_inst : DFF_X1 port map( D => n9555, CK => clk, Q => 
                           net227330, QN => n16092);
   registers_reg_66_24_inst : DFF_X1 port map( D => n9554, CK => clk, Q => 
                           net227329, QN => n16054);
   registers_reg_67_24_inst : DFF_X1 port map( D => n9553, CK => clk, Q => 
                           net271510, QN => n14273);
   registers_reg_68_24_inst : DFF_X1 port map( D => n9552, CK => clk, Q => 
                           registers_68_24_port, QN => n16180);
   registers_reg_69_24_inst : DFF_X1 port map( D => n9551, CK => clk, Q => 
                           net227328, QN => n16132);
   registers_reg_70_24_inst : DFF_X1 port map( D => n9550, CK => clk, Q => 
                           net227327, QN => n16044);
   registers_reg_0_23_inst : DFF_X1 port map( D => n9549, CK => clk, Q => 
                           registers_0_23_port, QN => n15874);
   registers_reg_1_23_inst : DFF_X1 port map( D => n9548, CK => clk, Q => 
                           registers_1_23_port, QN => n15631);
   registers_reg_2_23_inst : DFF_X1 port map( D => n9547, CK => clk, Q => 
                           registers_2_23_port, QN => n14757);
   registers_reg_3_23_inst : DFF_X1 port map( D => n9546, CK => clk, Q => 
                           net227326, QN => n15723);
   registers_reg_4_23_inst : DFF_X1 port map( D => n9545, CK => clk, Q => 
                           registers_4_23_port, QN => n15544);
   registers_reg_5_23_inst : DFF_X1 port map( D => n9544, CK => clk, Q => 
                           registers_5_23_port, QN => n14817);
   registers_reg_6_23_inst : DFF_X1 port map( D => n9543, CK => clk, Q => 
                           net271509, QN => n14050);
   registers_reg_7_23_inst : DFF_X1 port map( D => n9542, CK => clk, Q => 
                           registers_7_23_port, QN => n15319);
   registers_reg_8_23_inst : DFF_X1 port map( D => n9541, CK => clk, Q => 
                           net227325, QN => n15232);
   registers_reg_9_23_inst : DFF_X1 port map( D => n9540, CK => clk, Q => 
                           registers_9_23_port, QN => n14351);
   registers_reg_10_23_inst : DFF_X1 port map( D => n9539, CK => clk, Q => 
                           registers_10_23_port, QN => n14700);
   registers_reg_11_23_inst : DFF_X1 port map( D => n9538, CK => clk, Q => 
                           registers_11_23_port, QN => n14469);
   registers_reg_12_23_inst : DFF_X1 port map( D => n9537, CK => clk, Q => 
                           registers_12_23_port, QN => n15662);
   registers_reg_13_23_inst : DFF_X1 port map( D => n9536, CK => clk, Q => 
                           net227324, QN => n15115);
   registers_reg_14_23_inst : DFF_X1 port map( D => n9535, CK => clk, Q => 
                           net271508, QN => n11874);
   registers_reg_15_23_inst : DFF_X1 port map( D => n9534, CK => clk, Q => 
                           registers_15_23_port, QN => n15285);
   registers_reg_16_23_inst : DFF_X1 port map( D => n9533, CK => clk, Q => 
                           registers_16_23_port, QN => n15692);
   registers_reg_17_23_inst : DFF_X1 port map( D => n9532, CK => clk, Q => 
                           registers_17_23_port, QN => n14598);
   registers_reg_18_23_inst : DFF_X1 port map( D => n9531, CK => clk, Q => 
                           registers_18_23_port, QN => n14413);
   registers_reg_19_23_inst : DFF_X1 port map( D => n9530, CK => clk, Q => 
                           registers_19_23_port, QN => n15852);
   registers_reg_20_23_inst : DFF_X1 port map( D => n9529, CK => clk, Q => 
                           net271507, QN => n14824);
   registers_reg_21_23_inst : DFF_X1 port map( D => n9528, CK => clk, Q => 
                           net271506, QN => n12198);
   registers_reg_22_23_inst : DFF_X1 port map( D => n9527, CK => clk, Q => 
                           registers_22_23_port, QN => n15395);
   registers_reg_23_23_inst : DFF_X1 port map( D => n9526, CK => clk, Q => 
                           registers_23_23_port, QN => n15905);
   registers_reg_24_23_inst : DFF_X1 port map( D => n9525, CK => clk, Q => 
                           net227323, QN => n15202);
   registers_reg_25_23_inst : DFF_X1 port map( D => n9524, CK => clk, Q => 
                           registers_25_23_port, QN => n14321);
   registers_reg_26_23_inst : DFF_X1 port map( D => n9523, CK => clk, Q => 
                           net271505, QN => n14049);
   registers_reg_27_23_inst : DFF_X1 port map( D => n9522, CK => clk, Q => 
                           net271504, QN => n12040);
   registers_reg_28_23_inst : DFF_X1 port map( D => n9521, CK => clk, Q => 
                           net227322, QN => n15025);
   registers_reg_29_23_inst : DFF_X1 port map( D => n9520, CK => clk, Q => 
                           registers_29_23_port, QN => n15843);
   registers_reg_30_23_inst : DFF_X1 port map( D => n9519, CK => clk, Q => 
                           registers_30_23_port, QN => n14671);
   registers_reg_31_23_inst : DFF_X1 port map( D => n9518, CK => clk, Q => 
                           net227321, QN => n15722);
   registers_reg_32_23_inst : DFF_X1 port map( D => n9517, CK => clk, Q => 
                           net271503, QN => n12332);
   registers_reg_33_23_inst : DFF_X1 port map( D => n9516, CK => clk, Q => 
                           net271502, QN => n11867);
   registers_reg_34_23_inst : DFF_X1 port map( D => n9515, CK => clk, Q => 
                           registers_34_23_port, QN => n15488);
   registers_reg_35_23_inst : DFF_X1 port map( D => n9514, CK => clk, Q => 
                           net227320, QN => n15620);
   registers_reg_36_23_inst : DFF_X1 port map( D => n9513, CK => clk, Q => 
                           registers_36_23_port, QN => n15175);
   registers_reg_37_23_inst : DFF_X1 port map( D => n9512, CK => clk, Q => 
                           registers_37_23_port, QN => n14402);
   registers_reg_38_23_inst : DFF_X1 port map( D => n9511, CK => clk, Q => 
                           registers_38_23_port, QN => n15059);
   registers_reg_39_23_inst : DFF_X1 port map( D => n9510, CK => clk, Q => 
                           net271501, QN => n12164);
   registers_reg_40_23_inst : DFF_X1 port map( D => n9509, CK => clk, Q => 
                           registers_40_23_port, QN => n15116);
   registers_reg_41_23_inst : DFF_X1 port map( D => n9508, CK => clk, Q => 
                           registers_41_23_port, QN => n14470);
   registers_reg_42_23_inst : DFF_X1 port map( D => n9507, CK => clk, Q => 
                           registers_42_23_port, QN => n15950);
   registers_reg_43_23_inst : DFF_X1 port map( D => n9506, CK => clk, Q => 
                           registers_43_23_port, QN => n14909);
   registers_reg_44_23_inst : DFF_X1 port map( D => n9505, CK => clk, Q => 
                           registers_44_23_port, QN => n15459);
   registers_reg_45_23_inst : DFF_X1 port map( D => n9504, CK => clk, Q => 
                           registers_45_23_port, QN => n14758);
   registers_reg_46_23_inst : DFF_X1 port map( D => n9503, CK => clk, Q => 
                           net227319, QN => n12015);
   registers_reg_47_23_inst : DFF_X1 port map( D => n9502, CK => clk, Q => 
                           registers_47_23_port, QN => n14568);
   registers_reg_48_23_inst : DFF_X1 port map( D => n9501, CK => clk, Q => 
                           registers_48_23_port, QN => n15573);
   registers_reg_49_23_inst : DFF_X1 port map( D => n9500, CK => clk, Q => 
                           registers_49_23_port, QN => n14505);
   registers_reg_50_23_inst : DFF_X1 port map( D => n9499, CK => clk, Q => 
                           registers_50_23_port, QN => n15992);
   registers_reg_51_23_inst : DFF_X1 port map( D => n9498, CK => clk, Q => 
                           registers_51_23_port, QN => n15420);
   registers_reg_52_23_inst : DFF_X1 port map( D => n9497, CK => clk, Q => 
                           net227318, QN => n14959);
   registers_reg_53_23_inst : DFF_X1 port map( D => n9496, CK => clk, Q => 
                           net227317, QN => n15941);
   registers_reg_54_23_inst : DFF_X1 port map( D => n9495, CK => clk, Q => 
                           registers_54_23_port, QN => n14591);
   registers_reg_55_23_inst : DFF_X1 port map( D => n9494, CK => clk, Q => 
                           registers_55_23_port, QN => n12153);
   registers_reg_56_23_inst : DFF_X1 port map( D => n9493, CK => clk, Q => 
                           registers_56_23_port, QN => n16006);
   registers_reg_57_23_inst : DFF_X1 port map( D => n9492, CK => clk, Q => 
                           net227316, QN => n15263);
   registers_reg_58_23_inst : DFF_X1 port map( D => n9491, CK => clk, Q => 
                           net227315, QN => n14930);
   registers_reg_59_23_inst : DFF_X1 port map( D => n9490, CK => clk, Q => 
                           registers_59_23_port, QN => n15518);
   registers_reg_60_23_inst : DFF_X1 port map( D => n9489, CK => clk, Q => 
                           registers_60_23_port, QN => n14663);
   registers_reg_61_23_inst : DFF_X1 port map( D => n9488, CK => clk, Q => 
                           net227314, QN => n15654);
   registers_reg_62_23_inst : DFF_X1 port map( D => n9487, CK => clk, Q => 
                           registers_62_23_port, QN => n15143);
   registers_reg_63_23_inst : DFF_X1 port map( D => n9486, CK => clk, Q => 
                           registers_63_23_port, QN => n14526);
   to_mem_reg_23_inst : DFF_X1 port map( D => n9485, CK => clk, Q => net271500,
                           QN => n7702);
   registers_reg_64_23_inst : DFF_X1 port map( D => n9484, CK => clk, Q => 
                           net227313, QN => n16142);
   registers_reg_65_23_inst : DFF_X1 port map( D => n9483, CK => clk, Q => 
                           net227312, QN => n16091);
   registers_reg_66_23_inst : DFF_X1 port map( D => n9482, CK => clk, Q => 
                           net227311, QN => n16053);
   registers_reg_67_23_inst : DFF_X1 port map( D => n9481, CK => clk, Q => 
                           net271499, QN => n14272);
   registers_reg_68_23_inst : DFF_X1 port map( D => n9480, CK => clk, Q => 
                           registers_68_23_port, QN => n16179);
   registers_reg_69_23_inst : DFF_X1 port map( D => n9479, CK => clk, Q => 
                           net227310, QN => n16131);
   registers_reg_70_23_inst : DFF_X1 port map( D => n9478, CK => clk, Q => 
                           net227309, QN => n16043);
   registers_reg_0_22_inst : DFF_X1 port map( D => n9477, CK => clk, Q => 
                           registers_0_22_port, QN => n15873);
   registers_reg_1_22_inst : DFF_X1 port map( D => n9476, CK => clk, Q => 
                           registers_1_22_port, QN => n15630);
   registers_reg_2_22_inst : DFF_X1 port map( D => n9475, CK => clk, Q => 
                           registers_2_22_port, QN => n14813);
   registers_reg_3_22_inst : DFF_X1 port map( D => n9474, CK => clk, Q => 
                           net227308, QN => n15780);
   registers_reg_4_22_inst : DFF_X1 port map( D => n9473, CK => clk, Q => 
                           registers_4_22_port, QN => n15543);
   registers_reg_5_22_inst : DFF_X1 port map( D => n9472, CK => clk, Q => 
                           registers_5_22_port, QN => n14754);
   registers_reg_6_22_inst : DFF_X1 port map( D => n9471, CK => clk, Q => 
                           net271498, QN => n14048);
   registers_reg_7_22_inst : DFF_X1 port map( D => n9470, CK => clk, Q => 
                           registers_7_22_port, QN => n15348);
   registers_reg_8_22_inst : DFF_X1 port map( D => n9469, CK => clk, Q => 
                           net227307, QN => n15231);
   registers_reg_9_22_inst : DFF_X1 port map( D => n9468, CK => clk, Q => 
                           registers_9_22_port, QN => n14350);
   registers_reg_10_22_inst : DFF_X1 port map( D => n9467, CK => clk, Q => 
                           registers_10_22_port, QN => n14755);
   registers_reg_11_22_inst : DFF_X1 port map( D => n9466, CK => clk, Q => 
                           registers_11_22_port, QN => n14467);
   registers_reg_12_22_inst : DFF_X1 port map( D => n9465, CK => clk, Q => 
                           registers_12_22_port, QN => n15690);
   registers_reg_13_22_inst : DFF_X1 port map( D => n9464, CK => clk, Q => 
                           net227306, QN => n15113);
   registers_reg_14_22_inst : DFF_X1 port map( D => n9463, CK => clk, Q => 
                           net271497, QN => n11902);
   registers_reg_15_22_inst : DFF_X1 port map( D => n9462, CK => clk, Q => 
                           registers_15_22_port, QN => n15313);
   registers_reg_16_22_inst : DFF_X1 port map( D => n9461, CK => clk, Q => 
                           registers_16_22_port, QN => n15720);
   registers_reg_17_22_inst : DFF_X1 port map( D => n9460, CK => clk, Q => 
                           registers_17_22_port, QN => n14626);
   registers_reg_18_22_inst : DFF_X1 port map( D => n9459, CK => clk, Q => 
                           registers_18_22_port, QN => n14412);
   registers_reg_19_22_inst : DFF_X1 port map( D => n9458, CK => clk, Q => 
                           registers_19_22_port, QN => n15851);
   registers_reg_20_22_inst : DFF_X1 port map( D => n9457, CK => clk, Q => 
                           net271496, QN => n14852);
   registers_reg_21_22_inst : DFF_X1 port map( D => n9456, CK => clk, Q => 
                           net271495, QN => n12306);
   registers_reg_22_22_inst : DFF_X1 port map( D => n9455, CK => clk, Q => 
                           registers_22_22_port, QN => n15394);
   registers_reg_23_22_inst : DFF_X1 port map( D => n9454, CK => clk, Q => 
                           registers_23_22_port, QN => n15904);
   registers_reg_24_22_inst : DFF_X1 port map( D => n9453, CK => clk, Q => 
                           net227305, QN => n15201);
   registers_reg_25_22_inst : DFF_X1 port map( D => n9452, CK => clk, Q => 
                           registers_25_22_port, QN => n14320);
   registers_reg_26_22_inst : DFF_X1 port map( D => n9451, CK => clk, Q => 
                           net271494, QN => n14047);
   registers_reg_27_22_inst : DFF_X1 port map( D => n9450, CK => clk, Q => 
                           net271493, QN => n12039);
   registers_reg_28_22_inst : DFF_X1 port map( D => n9449, CK => clk, Q => 
                           net227304, QN => n15024);
   registers_reg_29_22_inst : DFF_X1 port map( D => n9448, CK => clk, Q => 
                           registers_29_22_port, QN => n15842);
   registers_reg_30_22_inst : DFF_X1 port map( D => n9447, CK => clk, Q => 
                           registers_30_22_port, QN => n14698);
   registers_reg_31_22_inst : DFF_X1 port map( D => n9446, CK => clk, Q => 
                           net227303, QN => n15756);
   registers_reg_32_22_inst : DFF_X1 port map( D => n9445, CK => clk, Q => 
                           net271492, QN => n12331);
   registers_reg_33_22_inst : DFF_X1 port map( D => n9444, CK => clk, Q => 
                           net271491, QN => n11866);
   registers_reg_34_22_inst : DFF_X1 port map( D => n9443, CK => clk, Q => 
                           registers_34_22_port, QN => n15516);
   registers_reg_35_22_inst : DFF_X1 port map( D => n9442, CK => clk, Q => 
                           net227302, QN => n15619);
   registers_reg_36_22_inst : DFF_X1 port map( D => n9441, CK => clk, Q => 
                           registers_36_22_port, QN => n15174);
   registers_reg_37_22_inst : DFF_X1 port map( D => n9440, CK => clk, Q => 
                           registers_37_22_port, QN => n14401);
   registers_reg_38_22_inst : DFF_X1 port map( D => n9439, CK => clk, Q => 
                           registers_38_22_port, QN => n15058);
   registers_reg_39_22_inst : DFF_X1 port map( D => n9438, CK => clk, Q => 
                           net271490, QN => n12193);
   registers_reg_40_22_inst : DFF_X1 port map( D => n9437, CK => clk, Q => 
                           registers_40_22_port, QN => n15114);
   registers_reg_41_22_inst : DFF_X1 port map( D => n9436, CK => clk, Q => 
                           registers_41_22_port, QN => n14468);
   registers_reg_42_22_inst : DFF_X1 port map( D => n9435, CK => clk, Q => 
                           registers_42_22_port, QN => n15949);
   registers_reg_43_22_inst : DFF_X1 port map( D => n9434, CK => clk, Q => 
                           registers_43_22_port, QN => n14908);
   registers_reg_44_22_inst : DFF_X1 port map( D => n9433, CK => clk, Q => 
                           registers_44_22_port, QN => n15486);
   registers_reg_45_22_inst : DFF_X1 port map( D => n9432, CK => clk, Q => 
                           registers_45_22_port, QN => n14814);
   registers_reg_46_22_inst : DFF_X1 port map( D => n9431, CK => clk, Q => 
                           net227301, QN => n12014);
   registers_reg_47_22_inst : DFF_X1 port map( D => n9430, CK => clk, Q => 
                           registers_47_22_port, QN => n14567);
   registers_reg_48_22_inst : DFF_X1 port map( D => n9429, CK => clk, Q => 
                           registers_48_22_port, QN => n15572);
   registers_reg_49_22_inst : DFF_X1 port map( D => n9428, CK => clk, Q => 
                           registers_49_22_port, QN => n14504);
   registers_reg_50_22_inst : DFF_X1 port map( D => n9427, CK => clk, Q => 
                           registers_50_22_port, QN => n15991);
   registers_reg_51_22_inst : DFF_X1 port map( D => n9426, CK => clk, Q => 
                           registers_51_22_port, QN => n15419);
   registers_reg_52_22_inst : DFF_X1 port map( D => n9425, CK => clk, Q => 
                           net227300, QN => n14958);
   registers_reg_53_22_inst : DFF_X1 port map( D => n9424, CK => clk, Q => 
                           net227299, QN => n15940);
   registers_reg_54_22_inst : DFF_X1 port map( D => n9423, CK => clk, Q => 
                           registers_54_22_port, QN => n14590);
   registers_reg_55_22_inst : DFF_X1 port map( D => n9422, CK => clk, Q => 
                           registers_55_22_port, QN => n12152);
   registers_reg_56_22_inst : DFF_X1 port map( D => n9421, CK => clk, Q => 
                           registers_56_22_port, QN => n16024);
   registers_reg_57_22_inst : DFF_X1 port map( D => n9420, CK => clk, Q => 
                           net227298, QN => n15262);
   registers_reg_58_22_inst : DFF_X1 port map( D => n9419, CK => clk, Q => 
                           net227297, QN => n14929);
   registers_reg_59_22_inst : DFF_X1 port map( D => n9418, CK => clk, Q => 
                           registers_59_22_port, QN => n15451);
   registers_reg_60_22_inst : DFF_X1 port map( D => n9417, CK => clk, Q => 
                           registers_60_22_port, QN => n14662);
   registers_reg_61_22_inst : DFF_X1 port map( D => n9416, CK => clk, Q => 
                           net227296, QN => n15653);
   registers_reg_62_22_inst : DFF_X1 port map( D => n9415, CK => clk, Q => 
                           registers_62_22_port, QN => n15142);
   registers_reg_63_22_inst : DFF_X1 port map( D => n9414, CK => clk, Q => 
                           registers_63_22_port, QN => n14525);
   to_mem_reg_22_inst : DFF_X1 port map( D => n9413, CK => clk, Q => net271489,
                           QN => n7703);
   registers_reg_64_22_inst : DFF_X1 port map( D => n9412, CK => clk, Q => 
                           net227295, QN => n16160);
   registers_reg_65_22_inst : DFF_X1 port map( D => n9411, CK => clk, Q => 
                           net227294, QN => n16110);
   registers_reg_66_22_inst : DFF_X1 port map( D => n9410, CK => clk, Q => 
                           net227293, QN => n16084);
   registers_reg_67_22_inst : DFF_X1 port map( D => n9409, CK => clk, Q => 
                           net271488, QN => n14268);
   registers_reg_68_22_inst : DFF_X1 port map( D => n9408, CK => clk, Q => 
                           registers_68_22_port, QN => n16198);
   registers_reg_69_22_inst : DFF_X1 port map( D => n9407, CK => clk, Q => 
                           net227292, QN => n16173);
   registers_reg_70_22_inst : DFF_X1 port map( D => n9406, CK => clk, Q => 
                           net227291, QN => n16083);
   registers_reg_0_21_inst : DFF_X1 port map( D => n9405, CK => clk, Q => 
                           registers_0_21_port, QN => n15872);
   registers_reg_1_21_inst : DFF_X1 port map( D => n9404, CK => clk, Q => 
                           registers_1_21_port, QN => n15629);
   registers_reg_2_21_inst : DFF_X1 port map( D => n9403, CK => clk, Q => 
                           registers_2_21_port, QN => n14811);
   registers_reg_3_21_inst : DFF_X1 port map( D => n9402, CK => clk, Q => 
                           net227290, QN => n15779);
   registers_reg_4_21_inst : DFF_X1 port map( D => n9401, CK => clk, Q => 
                           registers_4_21_port, QN => n15542);
   registers_reg_5_21_inst : DFF_X1 port map( D => n9400, CK => clk, Q => 
                           registers_5_21_port, QN => n14752);
   registers_reg_6_21_inst : DFF_X1 port map( D => n9399, CK => clk, Q => 
                           net271487, QN => n14046);
   registers_reg_7_21_inst : DFF_X1 port map( D => n9398, CK => clk, Q => 
                           registers_7_21_port, QN => n15347);
   registers_reg_8_21_inst : DFF_X1 port map( D => n9397, CK => clk, Q => 
                           net227289, QN => n15230);
   registers_reg_9_21_inst : DFF_X1 port map( D => n9396, CK => clk, Q => 
                           registers_9_21_port, QN => n14349);
   registers_reg_10_21_inst : DFF_X1 port map( D => n9395, CK => clk, Q => 
                           registers_10_21_port, QN => n14753);
   registers_reg_11_21_inst : DFF_X1 port map( D => n9394, CK => clk, Q => 
                           registers_11_21_port, QN => n14465);
   registers_reg_12_21_inst : DFF_X1 port map( D => n9393, CK => clk, Q => 
                           registers_12_21_port, QN => n15689);
   registers_reg_13_21_inst : DFF_X1 port map( D => n9392, CK => clk, Q => 
                           net227288, QN => n15111);
   registers_reg_14_21_inst : DFF_X1 port map( D => n9391, CK => clk, Q => 
                           net271486, QN => n11901);
   registers_reg_15_21_inst : DFF_X1 port map( D => n9390, CK => clk, Q => 
                           registers_15_21_port, QN => n15312);
   registers_reg_16_21_inst : DFF_X1 port map( D => n9389, CK => clk, Q => 
                           registers_16_21_port, QN => n15719);
   registers_reg_17_21_inst : DFF_X1 port map( D => n9388, CK => clk, Q => 
                           registers_17_21_port, QN => n14625);
   registers_reg_18_21_inst : DFF_X1 port map( D => n9387, CK => clk, Q => 
                           registers_18_21_port, QN => n14411);
   registers_reg_19_21_inst : DFF_X1 port map( D => n9386, CK => clk, Q => 
                           registers_19_21_port, QN => n15850);
   registers_reg_20_21_inst : DFF_X1 port map( D => n9385, CK => clk, Q => 
                           net271485, QN => n14851);
   registers_reg_21_21_inst : DFF_X1 port map( D => n9384, CK => clk, Q => 
                           net271484, QN => n12305);
   registers_reg_22_21_inst : DFF_X1 port map( D => n9383, CK => clk, Q => 
                           registers_22_21_port, QN => n15393);
   registers_reg_23_21_inst : DFF_X1 port map( D => n9382, CK => clk, Q => 
                           registers_23_21_port, QN => n15903);
   registers_reg_24_21_inst : DFF_X1 port map( D => n9381, CK => clk, Q => 
                           net227287, QN => n15200);
   registers_reg_25_21_inst : DFF_X1 port map( D => n9380, CK => clk, Q => 
                           registers_25_21_port, QN => n14319);
   registers_reg_26_21_inst : DFF_X1 port map( D => n9379, CK => clk, Q => 
                           net271483, QN => n14045);
   registers_reg_27_21_inst : DFF_X1 port map( D => n9378, CK => clk, Q => 
                           net271482, QN => n12038);
   registers_reg_28_21_inst : DFF_X1 port map( D => n9377, CK => clk, Q => 
                           net227286, QN => n15023);
   registers_reg_29_21_inst : DFF_X1 port map( D => n9376, CK => clk, Q => 
                           registers_29_21_port, QN => n15841);
   registers_reg_30_21_inst : DFF_X1 port map( D => n9375, CK => clk, Q => 
                           registers_30_21_port, QN => n14697);
   registers_reg_31_21_inst : DFF_X1 port map( D => n9374, CK => clk, Q => 
                           net227285, QN => n15755);
   registers_reg_32_21_inst : DFF_X1 port map( D => n9373, CK => clk, Q => 
                           net271481, QN => n12330);
   registers_reg_33_21_inst : DFF_X1 port map( D => n9372, CK => clk, Q => 
                           net271480, QN => n11865);
   registers_reg_34_21_inst : DFF_X1 port map( D => n9371, CK => clk, Q => 
                           registers_34_21_port, QN => n15515);
   registers_reg_35_21_inst : DFF_X1 port map( D => n9370, CK => clk, Q => 
                           net227284, QN => n15618);
   registers_reg_36_21_inst : DFF_X1 port map( D => n9369, CK => clk, Q => 
                           registers_36_21_port, QN => n15173);
   registers_reg_37_21_inst : DFF_X1 port map( D => n9368, CK => clk, Q => 
                           registers_37_21_port, QN => n14400);
   registers_reg_38_21_inst : DFF_X1 port map( D => n9367, CK => clk, Q => 
                           registers_38_21_port, QN => n15057);
   registers_reg_39_21_inst : DFF_X1 port map( D => n9366, CK => clk, Q => 
                           net271479, QN => n12192);
   registers_reg_40_21_inst : DFF_X1 port map( D => n9365, CK => clk, Q => 
                           registers_40_21_port, QN => n15112);
   registers_reg_41_21_inst : DFF_X1 port map( D => n9364, CK => clk, Q => 
                           registers_41_21_port, QN => n14466);
   registers_reg_42_21_inst : DFF_X1 port map( D => n9363, CK => clk, Q => 
                           registers_42_21_port, QN => n15948);
   registers_reg_43_21_inst : DFF_X1 port map( D => n9362, CK => clk, Q => 
                           registers_43_21_port, QN => n14907);
   registers_reg_44_21_inst : DFF_X1 port map( D => n9361, CK => clk, Q => 
                           registers_44_21_port, QN => n15485);
   registers_reg_45_21_inst : DFF_X1 port map( D => n9360, CK => clk, Q => 
                           registers_45_21_port, QN => n14812);
   registers_reg_46_21_inst : DFF_X1 port map( D => n9359, CK => clk, Q => 
                           net227283, QN => n12013);
   registers_reg_47_21_inst : DFF_X1 port map( D => n9358, CK => clk, Q => 
                           registers_47_21_port, QN => n14566);
   registers_reg_48_21_inst : DFF_X1 port map( D => n9357, CK => clk, Q => 
                           registers_48_21_port, QN => n15571);
   registers_reg_49_21_inst : DFF_X1 port map( D => n9356, CK => clk, Q => 
                           registers_49_21_port, QN => n14503);
   registers_reg_50_21_inst : DFF_X1 port map( D => n9355, CK => clk, Q => 
                           registers_50_21_port, QN => n15990);
   registers_reg_51_21_inst : DFF_X1 port map( D => n9354, CK => clk, Q => 
                           registers_51_21_port, QN => n15418);
   registers_reg_52_21_inst : DFF_X1 port map( D => n9353, CK => clk, Q => 
                           net227282, QN => n14957);
   registers_reg_53_21_inst : DFF_X1 port map( D => n9352, CK => clk, Q => 
                           net227281, QN => n15967);
   registers_reg_54_21_inst : DFF_X1 port map( D => n9351, CK => clk, Q => 
                           registers_54_21_port, QN => n14589);
   registers_reg_55_21_inst : DFF_X1 port map( D => n9350, CK => clk, Q => 
                           registers_55_21_port, QN => n12151);
   registers_reg_56_21_inst : DFF_X1 port map( D => n9349, CK => clk, Q => 
                           registers_56_21_port, QN => n16005);
   registers_reg_57_21_inst : DFF_X1 port map( D => n9348, CK => clk, Q => 
                           net227280, QN => n15261);
   registers_reg_58_21_inst : DFF_X1 port map( D => n9347, CK => clk, Q => 
                           net227279, QN => n14928);
   registers_reg_59_21_inst : DFF_X1 port map( D => n9346, CK => clk, Q => 
                           registers_59_21_port, QN => n15450);
   registers_reg_60_21_inst : DFF_X1 port map( D => n9345, CK => clk, Q => 
                           registers_60_21_port, QN => n14661);
   registers_reg_61_21_inst : DFF_X1 port map( D => n9344, CK => clk, Q => 
                           net227278, QN => n15652);
   registers_reg_62_21_inst : DFF_X1 port map( D => n9343, CK => clk, Q => 
                           registers_62_21_port, QN => n15141);
   registers_reg_63_21_inst : DFF_X1 port map( D => n9342, CK => clk, Q => 
                           registers_63_21_port, QN => n14524);
   to_mem_reg_21_inst : DFF_X1 port map( D => n9341, CK => clk, Q => net271478,
                           QN => n7704);
   registers_reg_64_21_inst : DFF_X1 port map( D => n9340, CK => clk, Q => 
                           net227277, QN => n16141);
   registers_reg_65_21_inst : DFF_X1 port map( D => n9339, CK => clk, Q => 
                           net227276, QN => n16090);
   registers_reg_66_21_inst : DFF_X1 port map( D => n9338, CK => clk, Q => 
                           net227275, QN => n16052);
   registers_reg_67_21_inst : DFF_X1 port map( D => n9337, CK => clk, Q => 
                           net271477, QN => n14271);
   registers_reg_68_21_inst : DFF_X1 port map( D => n9336, CK => clk, Q => 
                           registers_68_21_port, QN => n16178);
   registers_reg_69_21_inst : DFF_X1 port map( D => n9335, CK => clk, Q => 
                           net227274, QN => n16130);
   registers_reg_70_21_inst : DFF_X1 port map( D => n9334, CK => clk, Q => 
                           net227273, QN => n16042);
   registers_reg_0_20_inst : DFF_X1 port map( D => n9333, CK => clk, Q => 
                           registers_0_20_port, QN => n15871);
   registers_reg_1_20_inst : DFF_X1 port map( D => n9332, CK => clk, Q => 
                           registers_1_20_port, QN => n15628);
   registers_reg_2_20_inst : DFF_X1 port map( D => n9331, CK => clk, Q => 
                           registers_2_20_port, QN => n14809);
   registers_reg_3_20_inst : DFF_X1 port map( D => n9330, CK => clk, Q => 
                           net227272, QN => n15778);
   registers_reg_4_20_inst : DFF_X1 port map( D => n9329, CK => clk, Q => 
                           registers_4_20_port, QN => n15541);
   registers_reg_5_20_inst : DFF_X1 port map( D => n9328, CK => clk, Q => 
                           registers_5_20_port, QN => n14750);
   registers_reg_6_20_inst : DFF_X1 port map( D => n9327, CK => clk, Q => 
                           net271476, QN => n14044);
   registers_reg_7_20_inst : DFF_X1 port map( D => n9326, CK => clk, Q => 
                           registers_7_20_port, QN => n15346);
   registers_reg_8_20_inst : DFF_X1 port map( D => n9325, CK => clk, Q => 
                           net227271, QN => n15229);
   registers_reg_9_20_inst : DFF_X1 port map( D => n9324, CK => clk, Q => 
                           registers_9_20_port, QN => n14348);
   registers_reg_10_20_inst : DFF_X1 port map( D => n9323, CK => clk, Q => 
                           registers_10_20_port, QN => n14751);
   registers_reg_11_20_inst : DFF_X1 port map( D => n9322, CK => clk, Q => 
                           registers_11_20_port, QN => n14463);
   registers_reg_12_20_inst : DFF_X1 port map( D => n9321, CK => clk, Q => 
                           registers_12_20_port, QN => n15688);
   registers_reg_13_20_inst : DFF_X1 port map( D => n9320, CK => clk, Q => 
                           net227270, QN => n15109);
   registers_reg_14_20_inst : DFF_X1 port map( D => n9319, CK => clk, Q => 
                           net271475, QN => n11900);
   registers_reg_15_20_inst : DFF_X1 port map( D => n9318, CK => clk, Q => 
                           registers_15_20_port, QN => n15311);
   registers_reg_16_20_inst : DFF_X1 port map( D => n9317, CK => clk, Q => 
                           registers_16_20_port, QN => n15718);
   registers_reg_17_20_inst : DFF_X1 port map( D => n9316, CK => clk, Q => 
                           registers_17_20_port, QN => n14624);
   registers_reg_18_20_inst : DFF_X1 port map( D => n9315, CK => clk, Q => 
                           registers_18_20_port, QN => n14410);
   registers_reg_19_20_inst : DFF_X1 port map( D => n9314, CK => clk, Q => 
                           registers_19_20_port, QN => n15849);
   registers_reg_20_20_inst : DFF_X1 port map( D => n9313, CK => clk, Q => 
                           net271474, QN => n14850);
   registers_reg_21_20_inst : DFF_X1 port map( D => n9312, CK => clk, Q => 
                           net271473, QN => n12304);
   registers_reg_22_20_inst : DFF_X1 port map( D => n9311, CK => clk, Q => 
                           registers_22_20_port, QN => n15392);
   registers_reg_23_20_inst : DFF_X1 port map( D => n9310, CK => clk, Q => 
                           registers_23_20_port, QN => n15901);
   registers_reg_24_20_inst : DFF_X1 port map( D => n9309, CK => clk, Q => 
                           net227269, QN => n15199);
   registers_reg_25_20_inst : DFF_X1 port map( D => n9308, CK => clk, Q => 
                           registers_25_20_port, QN => n14318);
   registers_reg_26_20_inst : DFF_X1 port map( D => n9307, CK => clk, Q => 
                           net271472, QN => n14043);
   registers_reg_27_20_inst : DFF_X1 port map( D => n9306, CK => clk, Q => 
                           net271471, QN => n12037);
   registers_reg_28_20_inst : DFF_X1 port map( D => n9305, CK => clk, Q => 
                           net227268, QN => n15022);
   registers_reg_29_20_inst : DFF_X1 port map( D => n9304, CK => clk, Q => 
                           registers_29_20_port, QN => n15838);
   registers_reg_30_20_inst : DFF_X1 port map( D => n9303, CK => clk, Q => 
                           registers_30_20_port, QN => n14696);
   registers_reg_31_20_inst : DFF_X1 port map( D => n9302, CK => clk, Q => 
                           net227267, QN => n15754);
   registers_reg_32_20_inst : DFF_X1 port map( D => n9301, CK => clk, Q => 
                           net271470, QN => n12329);
   registers_reg_33_20_inst : DFF_X1 port map( D => n9300, CK => clk, Q => 
                           net271469, QN => n11864);
   registers_reg_34_20_inst : DFF_X1 port map( D => n9299, CK => clk, Q => 
                           registers_34_20_port, QN => n15514);
   registers_reg_35_20_inst : DFF_X1 port map( D => n9298, CK => clk, Q => 
                           net227266, QN => n15617);
   registers_reg_36_20_inst : DFF_X1 port map( D => n9297, CK => clk, Q => 
                           registers_36_20_port, QN => n15172);
   registers_reg_37_20_inst : DFF_X1 port map( D => n9296, CK => clk, Q => 
                           registers_37_20_port, QN => n14399);
   registers_reg_38_20_inst : DFF_X1 port map( D => n9295, CK => clk, Q => 
                           registers_38_20_port, QN => n15056);
   registers_reg_39_20_inst : DFF_X1 port map( D => n9294, CK => clk, Q => 
                           net271468, QN => n12191);
   registers_reg_40_20_inst : DFF_X1 port map( D => n9293, CK => clk, Q => 
                           registers_40_20_port, QN => n15110);
   registers_reg_41_20_inst : DFF_X1 port map( D => n9292, CK => clk, Q => 
                           registers_41_20_port, QN => n14464);
   registers_reg_42_20_inst : DFF_X1 port map( D => n9291, CK => clk, Q => 
                           registers_42_20_port, QN => n15947);
   registers_reg_43_20_inst : DFF_X1 port map( D => n9290, CK => clk, Q => 
                           registers_43_20_port, QN => n14906);
   registers_reg_44_20_inst : DFF_X1 port map( D => n9289, CK => clk, Q => 
                           registers_44_20_port, QN => n15484);
   registers_reg_45_20_inst : DFF_X1 port map( D => n9288, CK => clk, Q => 
                           registers_45_20_port, QN => n14810);
   registers_reg_46_20_inst : DFF_X1 port map( D => n9287, CK => clk, Q => 
                           net227265, QN => n12012);
   registers_reg_47_20_inst : DFF_X1 port map( D => n9286, CK => clk, Q => 
                           registers_47_20_port, QN => n14565);
   registers_reg_48_20_inst : DFF_X1 port map( D => n9285, CK => clk, Q => 
                           registers_48_20_port, QN => n15570);
   registers_reg_49_20_inst : DFF_X1 port map( D => n9284, CK => clk, Q => 
                           registers_49_20_port, QN => n14502);
   registers_reg_50_20_inst : DFF_X1 port map( D => n9283, CK => clk, Q => 
                           registers_50_20_port, QN => n15989);
   registers_reg_51_20_inst : DFF_X1 port map( D => n9282, CK => clk, Q => 
                           registers_51_20_port, QN => n15417);
   registers_reg_52_20_inst : DFF_X1 port map( D => n9281, CK => clk, Q => 
                           net227264, QN => n14956);
   registers_reg_53_20_inst : DFF_X1 port map( D => n9280, CK => clk, Q => 
                           net227263, QN => n15966);
   registers_reg_54_20_inst : DFF_X1 port map( D => n9279, CK => clk, Q => 
                           registers_54_20_port, QN => n14588);
   registers_reg_55_20_inst : DFF_X1 port map( D => n9278, CK => clk, Q => 
                           registers_55_20_port, QN => n12150);
   registers_reg_56_20_inst : DFF_X1 port map( D => n9277, CK => clk, Q => 
                           registers_56_20_port, QN => n16004);
   registers_reg_57_20_inst : DFF_X1 port map( D => n9276, CK => clk, Q => 
                           net227262, QN => n15260);
   registers_reg_58_20_inst : DFF_X1 port map( D => n9275, CK => clk, Q => 
                           net227261, QN => n14927);
   registers_reg_59_20_inst : DFF_X1 port map( D => n9274, CK => clk, Q => 
                           registers_59_20_port, QN => n15449);
   registers_reg_60_20_inst : DFF_X1 port map( D => n9273, CK => clk, Q => 
                           registers_60_20_port, QN => n14660);
   registers_reg_61_20_inst : DFF_X1 port map( D => n9272, CK => clk, Q => 
                           net227260, QN => n15651);
   registers_reg_62_20_inst : DFF_X1 port map( D => n9271, CK => clk, Q => 
                           registers_62_20_port, QN => n15140);
   registers_reg_63_20_inst : DFF_X1 port map( D => n9270, CK => clk, Q => 
                           registers_63_20_port, QN => n14523);
   to_mem_reg_20_inst : DFF_X1 port map( D => n9269, CK => clk, Q => net271467,
                           QN => n7705);
   registers_reg_64_20_inst : DFF_X1 port map( D => n9268, CK => clk, Q => 
                           net227259, QN => n16140);
   registers_reg_65_20_inst : DFF_X1 port map( D => n9267, CK => clk, Q => 
                           net227258, QN => n16089);
   registers_reg_66_20_inst : DFF_X1 port map( D => n9266, CK => clk, Q => 
                           net227257, QN => n16051);
   registers_reg_67_20_inst : DFF_X1 port map( D => n9265, CK => clk, Q => 
                           net271466, QN => n14270);
   registers_reg_68_20_inst : DFF_X1 port map( D => n9264, CK => clk, Q => 
                           registers_68_20_port, QN => n16177);
   registers_reg_69_20_inst : DFF_X1 port map( D => n9263, CK => clk, Q => 
                           net227256, QN => n16129);
   registers_reg_70_20_inst : DFF_X1 port map( D => n9262, CK => clk, Q => 
                           net227255, QN => n16082);
   registers_reg_0_19_inst : DFF_X1 port map( D => n9261, CK => clk, Q => 
                           registers_0_19_port, QN => n15870);
   registers_reg_1_19_inst : DFF_X1 port map( D => n9260, CK => clk, Q => 
                           registers_1_19_port, QN => n15627);
   registers_reg_2_19_inst : DFF_X1 port map( D => n9259, CK => clk, Q => 
                           registers_2_19_port, QN => n14807);
   registers_reg_3_19_inst : DFF_X1 port map( D => n9258, CK => clk, Q => 
                           net227254, QN => n15777);
   registers_reg_4_19_inst : DFF_X1 port map( D => n9257, CK => clk, Q => 
                           registers_4_19_port, QN => n15540);
   registers_reg_5_19_inst : DFF_X1 port map( D => n9256, CK => clk, Q => 
                           registers_5_19_port, QN => n14748);
   registers_reg_6_19_inst : DFF_X1 port map( D => n9255, CK => clk, Q => 
                           net271465, QN => n14042);
   registers_reg_7_19_inst : DFF_X1 port map( D => n9254, CK => clk, Q => 
                           registers_7_19_port, QN => n15345);
   registers_reg_8_19_inst : DFF_X1 port map( D => n9253, CK => clk, Q => 
                           net227253, QN => n15228);
   registers_reg_9_19_inst : DFF_X1 port map( D => n9252, CK => clk, Q => 
                           registers_9_19_port, QN => n14347);
   registers_reg_10_19_inst : DFF_X1 port map( D => n9251, CK => clk, Q => 
                           registers_10_19_port, QN => n14749);
   registers_reg_11_19_inst : DFF_X1 port map( D => n9250, CK => clk, Q => 
                           registers_11_19_port, QN => n14461);
   registers_reg_12_19_inst : DFF_X1 port map( D => n9249, CK => clk, Q => 
                           registers_12_19_port, QN => n15687);
   registers_reg_13_19_inst : DFF_X1 port map( D => n9248, CK => clk, Q => 
                           net227252, QN => n15107);
   registers_reg_14_19_inst : DFF_X1 port map( D => n9247, CK => clk, Q => 
                           net271464, QN => n11899);
   registers_reg_15_19_inst : DFF_X1 port map( D => n9246, CK => clk, Q => 
                           registers_15_19_port, QN => n15310);
   registers_reg_16_19_inst : DFF_X1 port map( D => n9245, CK => clk, Q => 
                           registers_16_19_port, QN => n15717);
   registers_reg_17_19_inst : DFF_X1 port map( D => n9244, CK => clk, Q => 
                           registers_17_19_port, QN => n14623);
   registers_reg_18_19_inst : DFF_X1 port map( D => n9243, CK => clk, Q => 
                           registers_18_19_port, QN => n14409);
   registers_reg_19_19_inst : DFF_X1 port map( D => n9242, CK => clk, Q => 
                           registers_19_19_port, QN => n15837);
   registers_reg_20_19_inst : DFF_X1 port map( D => n9241, CK => clk, Q => 
                           net271463, QN => n14849);
   registers_reg_21_19_inst : DFF_X1 port map( D => n9240, CK => clk, Q => 
                           net271462, QN => n12303);
   registers_reg_22_19_inst : DFF_X1 port map( D => n9239, CK => clk, Q => 
                           registers_22_19_port, QN => n15391);
   registers_reg_23_19_inst : DFF_X1 port map( D => n9238, CK => clk, Q => 
                           registers_23_19_port, QN => n15900);
   registers_reg_24_19_inst : DFF_X1 port map( D => n9237, CK => clk, Q => 
                           net227251, QN => n15198);
   registers_reg_25_19_inst : DFF_X1 port map( D => n9236, CK => clk, Q => 
                           registers_25_19_port, QN => n14317);
   registers_reg_26_19_inst : DFF_X1 port map( D => n9235, CK => clk, Q => 
                           net271461, QN => n14041);
   registers_reg_27_19_inst : DFF_X1 port map( D => n9234, CK => clk, Q => 
                           net271460, QN => n12036);
   registers_reg_28_19_inst : DFF_X1 port map( D => n9233, CK => clk, Q => 
                           net227250, QN => n15021);
   registers_reg_29_19_inst : DFF_X1 port map( D => n9232, CK => clk, Q => 
                           registers_29_19_port, QN => n15836);
   registers_reg_30_19_inst : DFF_X1 port map( D => n9231, CK => clk, Q => 
                           registers_30_19_port, QN => n14695);
   registers_reg_31_19_inst : DFF_X1 port map( D => n9230, CK => clk, Q => 
                           net227249, QN => n15753);
   registers_reg_32_19_inst : DFF_X1 port map( D => n9229, CK => clk, Q => 
                           net271459, QN => n12328);
   registers_reg_33_19_inst : DFF_X1 port map( D => n9228, CK => clk, Q => 
                           net271458, QN => n11863);
   registers_reg_34_19_inst : DFF_X1 port map( D => n9227, CK => clk, Q => 
                           registers_34_19_port, QN => n15513);
   registers_reg_35_19_inst : DFF_X1 port map( D => n9226, CK => clk, Q => 
                           net227248, QN => n15616);
   registers_reg_36_19_inst : DFF_X1 port map( D => n9225, CK => clk, Q => 
                           registers_36_19_port, QN => n15171);
   registers_reg_37_19_inst : DFF_X1 port map( D => n9224, CK => clk, Q => 
                           registers_37_19_port, QN => n14398);
   registers_reg_38_19_inst : DFF_X1 port map( D => n9223, CK => clk, Q => 
                           registers_38_19_port, QN => n15055);
   registers_reg_39_19_inst : DFF_X1 port map( D => n9222, CK => clk, Q => 
                           net271457, QN => n12190);
   registers_reg_40_19_inst : DFF_X1 port map( D => n9221, CK => clk, Q => 
                           registers_40_19_port, QN => n15108);
   registers_reg_41_19_inst : DFF_X1 port map( D => n9220, CK => clk, Q => 
                           registers_41_19_port, QN => n14462);
   registers_reg_42_19_inst : DFF_X1 port map( D => n9219, CK => clk, Q => 
                           registers_42_19_port, QN => n15938);
   registers_reg_43_19_inst : DFF_X1 port map( D => n9218, CK => clk, Q => 
                           registers_43_19_port, QN => n14905);
   registers_reg_44_19_inst : DFF_X1 port map( D => n9217, CK => clk, Q => 
                           registers_44_19_port, QN => n15483);
   registers_reg_45_19_inst : DFF_X1 port map( D => n9216, CK => clk, Q => 
                           registers_45_19_port, QN => n14808);
   registers_reg_46_19_inst : DFF_X1 port map( D => n9215, CK => clk, Q => 
                           net227247, QN => n12011);
   registers_reg_47_19_inst : DFF_X1 port map( D => n9214, CK => clk, Q => 
                           registers_47_19_port, QN => n14564);
   registers_reg_48_19_inst : DFF_X1 port map( D => n9213, CK => clk, Q => 
                           registers_48_19_port, QN => n15569);
   registers_reg_49_19_inst : DFF_X1 port map( D => n9212, CK => clk, Q => 
                           registers_49_19_port, QN => n14501);
   registers_reg_50_19_inst : DFF_X1 port map( D => n9211, CK => clk, Q => 
                           registers_50_19_port, QN => n15987);
   registers_reg_51_19_inst : DFF_X1 port map( D => n9210, CK => clk, Q => 
                           registers_51_19_port, QN => n15416);
   registers_reg_52_19_inst : DFF_X1 port map( D => n9209, CK => clk, Q => 
                           net227246, QN => n14955);
   registers_reg_53_19_inst : DFF_X1 port map( D => n9208, CK => clk, Q => 
                           net227245, QN => n15965);
   registers_reg_54_19_inst : DFF_X1 port map( D => n9207, CK => clk, Q => 
                           registers_54_19_port, QN => n14587);
   registers_reg_55_19_inst : DFF_X1 port map( D => n9206, CK => clk, Q => 
                           registers_55_19_port, QN => n12148);
   registers_reg_56_19_inst : DFF_X1 port map( D => n9205, CK => clk, Q => 
                           registers_56_19_port, QN => n16023);
   registers_reg_57_19_inst : DFF_X1 port map( D => n9204, CK => clk, Q => 
                           net227244, QN => n15259);
   registers_reg_58_19_inst : DFF_X1 port map( D => n9203, CK => clk, Q => 
                           net227243, QN => n14926);
   registers_reg_59_19_inst : DFF_X1 port map( D => n9202, CK => clk, Q => 
                           registers_59_19_port, QN => n15448);
   registers_reg_60_19_inst : DFF_X1 port map( D => n9201, CK => clk, Q => 
                           registers_60_19_port, QN => n14659);
   registers_reg_61_19_inst : DFF_X1 port map( D => n9200, CK => clk, Q => 
                           net227242, QN => n15650);
   registers_reg_62_19_inst : DFF_X1 port map( D => n9199, CK => clk, Q => 
                           registers_62_19_port, QN => n15139);
   registers_reg_63_19_inst : DFF_X1 port map( D => n9198, CK => clk, Q => 
                           registers_63_19_port, QN => n14522);
   to_mem_reg_19_inst : DFF_X1 port map( D => n9197, CK => clk, Q => net271456,
                           QN => n7706);
   registers_reg_64_19_inst : DFF_X1 port map( D => n9196, CK => clk, Q => 
                           net227241, QN => n16139);
   registers_reg_65_19_inst : DFF_X1 port map( D => n9195, CK => clk, Q => 
                           net227240, QN => n16088);
   registers_reg_66_19_inst : DFF_X1 port map( D => n9194, CK => clk, Q => 
                           net227239, QN => n16050);
   registers_reg_67_19_inst : DFF_X1 port map( D => n9193, CK => clk, Q => 
                           net271455, QN => n14269);
   registers_reg_68_19_inst : DFF_X1 port map( D => n9192, CK => clk, Q => 
                           registers_68_19_port, QN => n16176);
   registers_reg_69_19_inst : DFF_X1 port map( D => n9191, CK => clk, Q => 
                           net227238, QN => n16172);
   registers_reg_70_19_inst : DFF_X1 port map( D => n9190, CK => clk, Q => 
                           net227237, QN => n16085);
   registers_reg_0_18_inst : DFF_X1 port map( D => n9189, CK => clk, Q => 
                           registers_0_18_port, QN => n15869);
   registers_reg_1_18_inst : DFF_X1 port map( D => n9188, CK => clk, Q => 
                           registers_1_18_port, QN => n15626);
   registers_reg_2_18_inst : DFF_X1 port map( D => n9187, CK => clk, Q => 
                           registers_2_18_port, QN => n14805);
   registers_reg_3_18_inst : DFF_X1 port map( D => n9186, CK => clk, Q => 
                           net227236, QN => n15776);
   registers_reg_4_18_inst : DFF_X1 port map( D => n9185, CK => clk, Q => 
                           registers_4_18_port, QN => n15539);
   registers_reg_5_18_inst : DFF_X1 port map( D => n9184, CK => clk, Q => 
                           registers_5_18_port, QN => n14746);
   registers_reg_6_18_inst : DFF_X1 port map( D => n9183, CK => clk, Q => 
                           net271454, QN => n14040);
   registers_reg_7_18_inst : DFF_X1 port map( D => n9182, CK => clk, Q => 
                           registers_7_18_port, QN => n15344);
   registers_reg_8_18_inst : DFF_X1 port map( D => n9181, CK => clk, Q => 
                           net227235, QN => n15227);
   registers_reg_9_18_inst : DFF_X1 port map( D => n9180, CK => clk, Q => 
                           registers_9_18_port, QN => n14346);
   registers_reg_10_18_inst : DFF_X1 port map( D => n9179, CK => clk, Q => 
                           registers_10_18_port, QN => n14747);
   registers_reg_11_18_inst : DFF_X1 port map( D => n9178, CK => clk, Q => 
                           registers_11_18_port, QN => n14459);
   registers_reg_12_18_inst : DFF_X1 port map( D => n9177, CK => clk, Q => 
                           registers_12_18_port, QN => n15686);
   registers_reg_13_18_inst : DFF_X1 port map( D => n9176, CK => clk, Q => 
                           net227234, QN => n15105);
   registers_reg_14_18_inst : DFF_X1 port map( D => n9175, CK => clk, Q => 
                           net271453, QN => n11898);
   registers_reg_15_18_inst : DFF_X1 port map( D => n9174, CK => clk, Q => 
                           registers_15_18_port, QN => n15309);
   registers_reg_16_18_inst : DFF_X1 port map( D => n9173, CK => clk, Q => 
                           registers_16_18_port, QN => n15716);
   registers_reg_17_18_inst : DFF_X1 port map( D => n9172, CK => clk, Q => 
                           registers_17_18_port, QN => n14622);
   registers_reg_18_18_inst : DFF_X1 port map( D => n9171, CK => clk, Q => 
                           registers_18_18_port, QN => n14408);
   registers_reg_19_18_inst : DFF_X1 port map( D => n9170, CK => clk, Q => 
                           registers_19_18_port, QN => n15835);
   registers_reg_20_18_inst : DFF_X1 port map( D => n9169, CK => clk, Q => 
                           net271452, QN => n14848);
   registers_reg_21_18_inst : DFF_X1 port map( D => n9168, CK => clk, Q => 
                           net271451, QN => n12301);
   registers_reg_22_18_inst : DFF_X1 port map( D => n9167, CK => clk, Q => 
                           registers_22_18_port, QN => n15389);
   registers_reg_23_18_inst : DFF_X1 port map( D => n9166, CK => clk, Q => 
                           registers_23_18_port, QN => n15899);
   registers_reg_24_18_inst : DFF_X1 port map( D => n9165, CK => clk, Q => 
                           net227233, QN => n15197);
   registers_reg_25_18_inst : DFF_X1 port map( D => n9164, CK => clk, Q => 
                           registers_25_18_port, QN => n14316);
   registers_reg_26_18_inst : DFF_X1 port map( D => n9163, CK => clk, Q => 
                           net271450, QN => n14039);
   registers_reg_27_18_inst : DFF_X1 port map( D => n9162, CK => clk, Q => 
                           net271449, QN => n12035);
   registers_reg_28_18_inst : DFF_X1 port map( D => n9161, CK => clk, Q => 
                           net227232, QN => n15020);
   registers_reg_29_18_inst : DFF_X1 port map( D => n9160, CK => clk, Q => 
                           registers_29_18_port, QN => n15834);
   registers_reg_30_18_inst : DFF_X1 port map( D => n9159, CK => clk, Q => 
                           registers_30_18_port, QN => n14694);
   registers_reg_31_18_inst : DFF_X1 port map( D => n9158, CK => clk, Q => 
                           net227231, QN => n15752);
   registers_reg_32_18_inst : DFF_X1 port map( D => n9157, CK => clk, Q => 
                           net271448, QN => n12327);
   registers_reg_33_18_inst : DFF_X1 port map( D => n9156, CK => clk, Q => 
                           net271447, QN => n11862);
   registers_reg_34_18_inst : DFF_X1 port map( D => n9155, CK => clk, Q => 
                           registers_34_18_port, QN => n15512);
   registers_reg_35_18_inst : DFF_X1 port map( D => n9154, CK => clk, Q => 
                           net227230, QN => n15613);
   registers_reg_36_18_inst : DFF_X1 port map( D => n9153, CK => clk, Q => 
                           registers_36_18_port, QN => n15170);
   registers_reg_37_18_inst : DFF_X1 port map( D => n9152, CK => clk, Q => 
                           registers_37_18_port, QN => n14395);
   registers_reg_38_18_inst : DFF_X1 port map( D => n9151, CK => clk, Q => 
                           registers_38_18_port, QN => n15053);
   registers_reg_39_18_inst : DFF_X1 port map( D => n9150, CK => clk, Q => 
                           net271446, QN => n12189);
   registers_reg_40_18_inst : DFF_X1 port map( D => n9149, CK => clk, Q => 
                           registers_40_18_port, QN => n15106);
   registers_reg_41_18_inst : DFF_X1 port map( D => n9148, CK => clk, Q => 
                           registers_41_18_port, QN => n14460);
   registers_reg_42_18_inst : DFF_X1 port map( D => n9147, CK => clk, Q => 
                           registers_42_18_port, QN => n15937);
   registers_reg_43_18_inst : DFF_X1 port map( D => n9146, CK => clk, Q => 
                           registers_43_18_port, QN => n14904);
   registers_reg_44_18_inst : DFF_X1 port map( D => n9145, CK => clk, Q => 
                           registers_44_18_port, QN => n15482);
   registers_reg_45_18_inst : DFF_X1 port map( D => n9144, CK => clk, Q => 
                           registers_45_18_port, QN => n14806);
   registers_reg_46_18_inst : DFF_X1 port map( D => n9143, CK => clk, Q => 
                           net227229, QN => n12010);
   registers_reg_47_18_inst : DFF_X1 port map( D => n9142, CK => clk, Q => 
                           registers_47_18_port, QN => n14563);
   registers_reg_48_18_inst : DFF_X1 port map( D => n9141, CK => clk, Q => 
                           registers_48_18_port, QN => n15568);
   registers_reg_49_18_inst : DFF_X1 port map( D => n9140, CK => clk, Q => 
                           registers_49_18_port, QN => n14500);
   registers_reg_50_18_inst : DFF_X1 port map( D => n9139, CK => clk, Q => 
                           registers_50_18_port, QN => n15986);
   registers_reg_51_18_inst : DFF_X1 port map( D => n9138, CK => clk, Q => 
                           registers_51_18_port, QN => n15415);
   registers_reg_52_18_inst : DFF_X1 port map( D => n9137, CK => clk, Q => 
                           net227228, QN => n14954);
   registers_reg_53_18_inst : DFF_X1 port map( D => n9136, CK => clk, Q => 
                           net227227, QN => n15964);
   registers_reg_54_18_inst : DFF_X1 port map( D => n9135, CK => clk, Q => 
                           registers_54_18_port, QN => n14586);
   registers_reg_55_18_inst : DFF_X1 port map( D => n9134, CK => clk, Q => 
                           registers_55_18_port, QN => n12105);
   registers_reg_56_18_inst : DFF_X1 port map( D => n9133, CK => clk, Q => 
                           registers_56_18_port, QN => n16022);
   registers_reg_57_18_inst : DFF_X1 port map( D => n9132, CK => clk, Q => 
                           net227226, QN => n15258);
   registers_reg_58_18_inst : DFF_X1 port map( D => n9131, CK => clk, Q => 
                           net227225, QN => n14925);
   registers_reg_59_18_inst : DFF_X1 port map( D => n9130, CK => clk, Q => 
                           registers_59_18_port, QN => n15447);
   registers_reg_60_18_inst : DFF_X1 port map( D => n9129, CK => clk, Q => 
                           registers_60_18_port, QN => n14658);
   registers_reg_61_18_inst : DFF_X1 port map( D => n9128, CK => clk, Q => 
                           net227224, QN => n15649);
   registers_reg_62_18_inst : DFF_X1 port map( D => n9127, CK => clk, Q => 
                           registers_62_18_port, QN => n15138);
   registers_reg_63_18_inst : DFF_X1 port map( D => n9126, CK => clk, Q => 
                           registers_63_18_port, QN => n14521);
   to_mem_reg_18_inst : DFF_X1 port map( D => n9125, CK => clk, Q => net271445,
                           QN => n7707);
   registers_reg_64_18_inst : DFF_X1 port map( D => n9124, CK => clk, Q => 
                           net227223, QN => n16138);
   registers_reg_65_18_inst : DFF_X1 port map( D => n9123, CK => clk, Q => 
                           net227222, QN => n16109);
   registers_reg_66_18_inst : DFF_X1 port map( D => n9122, CK => clk, Q => 
                           net227221, QN => n16081);
   registers_reg_67_18_inst : DFF_X1 port map( D => n9121, CK => clk, Q => 
                           net271444, QN => n14264);
   registers_reg_68_18_inst : DFF_X1 port map( D => n9120, CK => clk, Q => 
                           registers_68_18_port, QN => n16197);
   registers_reg_69_18_inst : DFF_X1 port map( D => n9119, CK => clk, Q => 
                           net227220, QN => n16171);
   registers_reg_70_18_inst : DFF_X1 port map( D => n9118, CK => clk, Q => 
                           net227219, QN => n16080);
   registers_reg_0_17_inst : DFF_X1 port map( D => n9117, CK => clk, Q => 
                           registers_0_17_port, QN => n15868);
   registers_reg_1_17_inst : DFF_X1 port map( D => n9116, CK => clk, Q => 
                           registers_1_17_port, QN => n15612);
   registers_reg_2_17_inst : DFF_X1 port map( D => n9115, CK => clk, Q => 
                           registers_2_17_port, QN => n14803);
   registers_reg_3_17_inst : DFF_X1 port map( D => n9114, CK => clk, Q => 
                           net227218, QN => n15775);
   registers_reg_4_17_inst : DFF_X1 port map( D => n9113, CK => clk, Q => 
                           registers_4_17_port, QN => n15538);
   registers_reg_5_17_inst : DFF_X1 port map( D => n9112, CK => clk, Q => 
                           registers_5_17_port, QN => n14744);
   registers_reg_6_17_inst : DFF_X1 port map( D => n9111, CK => clk, Q => 
                           net271443, QN => n14038);
   registers_reg_7_17_inst : DFF_X1 port map( D => n9110, CK => clk, Q => 
                           registers_7_17_port, QN => n15343);
   registers_reg_8_17_inst : DFF_X1 port map( D => n9109, CK => clk, Q => 
                           net227217, QN => n15226);
   registers_reg_9_17_inst : DFF_X1 port map( D => n9108, CK => clk, Q => 
                           registers_9_17_port, QN => n14345);
   registers_reg_10_17_inst : DFF_X1 port map( D => n9107, CK => clk, Q => 
                           registers_10_17_port, QN => n14745);
   registers_reg_11_17_inst : DFF_X1 port map( D => n9106, CK => clk, Q => 
                           registers_11_17_port, QN => n14457);
   registers_reg_12_17_inst : DFF_X1 port map( D => n9105, CK => clk, Q => 
                           registers_12_17_port, QN => n15685);
   registers_reg_13_17_inst : DFF_X1 port map( D => n9104, CK => clk, Q => 
                           net227216, QN => n15103);
   registers_reg_14_17_inst : DFF_X1 port map( D => n9103, CK => clk, Q => 
                           net271442, QN => n11897);
   registers_reg_15_17_inst : DFF_X1 port map( D => n9102, CK => clk, Q => 
                           registers_15_17_port, QN => n15308);
   registers_reg_16_17_inst : DFF_X1 port map( D => n9101, CK => clk, Q => 
                           registers_16_17_port, QN => n15715);
   registers_reg_17_17_inst : DFF_X1 port map( D => n9100, CK => clk, Q => 
                           registers_17_17_port, QN => n14621);
   registers_reg_18_17_inst : DFF_X1 port map( D => n9099, CK => clk, Q => 
                           registers_18_17_port, QN => n14394);
   registers_reg_19_17_inst : DFF_X1 port map( D => n9098, CK => clk, Q => 
                           registers_19_17_port, QN => n15833);
   registers_reg_20_17_inst : DFF_X1 port map( D => n9097, CK => clk, Q => 
                           net271441, QN => n14847);
   registers_reg_21_17_inst : DFF_X1 port map( D => n9096, CK => clk, Q => 
                           net271440, QN => n12258);
   registers_reg_22_17_inst : DFF_X1 port map( D => n9095, CK => clk, Q => 
                           registers_22_17_port, QN => n15388);
   registers_reg_23_17_inst : DFF_X1 port map( D => n9094, CK => clk, Q => 
                           registers_23_17_port, QN => n15898);
   registers_reg_24_17_inst : DFF_X1 port map( D => n9093, CK => clk, Q => 
                           net227215, QN => n15196);
   registers_reg_25_17_inst : DFF_X1 port map( D => n9092, CK => clk, Q => 
                           registers_25_17_port, QN => n14315);
   registers_reg_26_17_inst : DFF_X1 port map( D => n9091, CK => clk, Q => 
                           net271439, QN => n14037);
   registers_reg_27_17_inst : DFF_X1 port map( D => n9090, CK => clk, Q => 
                           net271438, QN => n12034);
   registers_reg_28_17_inst : DFF_X1 port map( D => n9089, CK => clk, Q => 
                           net227214, QN => n15019);
   registers_reg_29_17_inst : DFF_X1 port map( D => n9088, CK => clk, Q => 
                           registers_29_17_port, QN => n15832);
   registers_reg_30_17_inst : DFF_X1 port map( D => n9087, CK => clk, Q => 
                           registers_30_17_port, QN => n14693);
   registers_reg_31_17_inst : DFF_X1 port map( D => n9086, CK => clk, Q => 
                           net227213, QN => n15751);
   registers_reg_32_17_inst : DFF_X1 port map( D => n9085, CK => clk, Q => 
                           net271437, QN => n12326);
   registers_reg_33_17_inst : DFF_X1 port map( D => n9084, CK => clk, Q => 
                           net271436, QN => n11860);
   registers_reg_34_17_inst : DFF_X1 port map( D => n9083, CK => clk, Q => 
                           registers_34_17_port, QN => n15511);
   registers_reg_35_17_inst : DFF_X1 port map( D => n9082, CK => clk, Q => 
                           net227212, QN => n15611);
   registers_reg_36_17_inst : DFF_X1 port map( D => n9081, CK => clk, Q => 
                           registers_36_17_port, QN => n15168);
   registers_reg_37_17_inst : DFF_X1 port map( D => n9080, CK => clk, Q => 
                           registers_37_17_port, QN => n14393);
   registers_reg_38_17_inst : DFF_X1 port map( D => n9079, CK => clk, Q => 
                           registers_38_17_port, QN => n15052);
   registers_reg_39_17_inst : DFF_X1 port map( D => n9078, CK => clk, Q => 
                           net271435, QN => n12188);
   registers_reg_40_17_inst : DFF_X1 port map( D => n9077, CK => clk, Q => 
                           registers_40_17_port, QN => n15104);
   registers_reg_41_17_inst : DFF_X1 port map( D => n9076, CK => clk, Q => 
                           registers_41_17_port, QN => n14458);
   registers_reg_42_17_inst : DFF_X1 port map( D => n9075, CK => clk, Q => 
                           registers_42_17_port, QN => n15936);
   registers_reg_43_17_inst : DFF_X1 port map( D => n9074, CK => clk, Q => 
                           registers_43_17_port, QN => n14903);
   registers_reg_44_17_inst : DFF_X1 port map( D => n9073, CK => clk, Q => 
                           registers_44_17_port, QN => n15481);
   registers_reg_45_17_inst : DFF_X1 port map( D => n9072, CK => clk, Q => 
                           registers_45_17_port, QN => n14804);
   registers_reg_46_17_inst : DFF_X1 port map( D => n9071, CK => clk, Q => 
                           net227211, QN => n12009);
   registers_reg_47_17_inst : DFF_X1 port map( D => n9070, CK => clk, Q => 
                           registers_47_17_port, QN => n14562);
   registers_reg_48_17_inst : DFF_X1 port map( D => n9069, CK => clk, Q => 
                           registers_48_17_port, QN => n15567);
   registers_reg_49_17_inst : DFF_X1 port map( D => n9068, CK => clk, Q => 
                           registers_49_17_port, QN => n14499);
   registers_reg_50_17_inst : DFF_X1 port map( D => n9067, CK => clk, Q => 
                           registers_50_17_port, QN => n15985);
   registers_reg_51_17_inst : DFF_X1 port map( D => n9066, CK => clk, Q => 
                           registers_51_17_port, QN => n15414);
   registers_reg_52_17_inst : DFF_X1 port map( D => n9065, CK => clk, Q => 
                           net227210, QN => n14953);
   registers_reg_53_17_inst : DFF_X1 port map( D => n9064, CK => clk, Q => 
                           net227209, QN => n15963);
   registers_reg_54_17_inst : DFF_X1 port map( D => n9063, CK => clk, Q => 
                           registers_54_17_port, QN => n14585);
   registers_reg_55_17_inst : DFF_X1 port map( D => n9062, CK => clk, Q => 
                           registers_55_17_port, QN => n12104);
   registers_reg_56_17_inst : DFF_X1 port map( D => n9061, CK => clk, Q => 
                           registers_56_17_port, QN => n16021);
   registers_reg_57_17_inst : DFF_X1 port map( D => n9060, CK => clk, Q => 
                           net227208, QN => n15257);
   registers_reg_58_17_inst : DFF_X1 port map( D => n9059, CK => clk, Q => 
                           net227207, QN => n14924);
   registers_reg_59_17_inst : DFF_X1 port map( D => n9058, CK => clk, Q => 
                           registers_59_17_port, QN => n15446);
   registers_reg_60_17_inst : DFF_X1 port map( D => n9057, CK => clk, Q => 
                           registers_60_17_port, QN => n14657);
   registers_reg_61_17_inst : DFF_X1 port map( D => n9056, CK => clk, Q => 
                           net227206, QN => n15648);
   registers_reg_62_17_inst : DFF_X1 port map( D => n9055, CK => clk, Q => 
                           registers_62_17_port, QN => n15137);
   registers_reg_63_17_inst : DFF_X1 port map( D => n9054, CK => clk, Q => 
                           registers_63_17_port, QN => n14520);
   to_mem_reg_17_inst : DFF_X1 port map( D => n9053, CK => clk, Q => net271434,
                           QN => n7708);
   registers_reg_64_17_inst : DFF_X1 port map( D => n9052, CK => clk, Q => 
                           net227205, QN => n16159);
   registers_reg_65_17_inst : DFF_X1 port map( D => n9051, CK => clk, Q => 
                           net227204, QN => n16108);
   registers_reg_66_17_inst : DFF_X1 port map( D => n9050, CK => clk, Q => 
                           net227203, QN => n16079);
   registers_reg_67_17_inst : DFF_X1 port map( D => n9049, CK => clk, Q => 
                           net271433, QN => n14261);
   registers_reg_68_17_inst : DFF_X1 port map( D => n9048, CK => clk, Q => 
                           registers_68_17_port, QN => n16196);
   registers_reg_69_17_inst : DFF_X1 port map( D => n9047, CK => clk, Q => 
                           net227202, QN => n16170);
   registers_reg_70_17_inst : DFF_X1 port map( D => n9046, CK => clk, Q => 
                           net227201, QN => n16078);
   registers_reg_0_16_inst : DFF_X1 port map( D => n9045, CK => clk, Q => 
                           registers_0_16_port, QN => n15867);
   registers_reg_1_16_inst : DFF_X1 port map( D => n9044, CK => clk, Q => 
                           registers_1_16_port, QN => n15610);
   registers_reg_2_16_inst : DFF_X1 port map( D => n9043, CK => clk, Q => 
                           registers_2_16_port, QN => n14801);
   registers_reg_3_16_inst : DFF_X1 port map( D => n9042, CK => clk, Q => 
                           net227200, QN => n15774);
   registers_reg_4_16_inst : DFF_X1 port map( D => n9041, CK => clk, Q => 
                           registers_4_16_port, QN => n15537);
   registers_reg_5_16_inst : DFF_X1 port map( D => n9040, CK => clk, Q => 
                           registers_5_16_port, QN => n14742);
   registers_reg_6_16_inst : DFF_X1 port map( D => n9039, CK => clk, Q => 
                           net271432, QN => n14036);
   registers_reg_7_16_inst : DFF_X1 port map( D => n9038, CK => clk, Q => 
                           registers_7_16_port, QN => n15342);
   registers_reg_8_16_inst : DFF_X1 port map( D => n9037, CK => clk, Q => 
                           net227199, QN => n15225);
   registers_reg_9_16_inst : DFF_X1 port map( D => n9036, CK => clk, Q => 
                           registers_9_16_port, QN => n14344);
   registers_reg_10_16_inst : DFF_X1 port map( D => n9035, CK => clk, Q => 
                           registers_10_16_port, QN => n14743);
   registers_reg_11_16_inst : DFF_X1 port map( D => n9034, CK => clk, Q => 
                           registers_11_16_port, QN => n14455);
   registers_reg_12_16_inst : DFF_X1 port map( D => n9033, CK => clk, Q => 
                           registers_12_16_port, QN => n15684);
   registers_reg_13_16_inst : DFF_X1 port map( D => n9032, CK => clk, Q => 
                           net227198, QN => n15101);
   registers_reg_14_16_inst : DFF_X1 port map( D => n9031, CK => clk, Q => 
                           net271431, QN => n11896);
   registers_reg_15_16_inst : DFF_X1 port map( D => n9030, CK => clk, Q => 
                           registers_15_16_port, QN => n15307);
   registers_reg_16_16_inst : DFF_X1 port map( D => n9029, CK => clk, Q => 
                           registers_16_16_port, QN => n15714);
   registers_reg_17_16_inst : DFF_X1 port map( D => n9028, CK => clk, Q => 
                           registers_17_16_port, QN => n14620);
   registers_reg_18_16_inst : DFF_X1 port map( D => n9027, CK => clk, Q => 
                           registers_18_16_port, QN => n14392);
   registers_reg_19_16_inst : DFF_X1 port map( D => n9026, CK => clk, Q => 
                           registers_19_16_port, QN => n15831);
   registers_reg_20_16_inst : DFF_X1 port map( D => n9025, CK => clk, Q => 
                           net271430, QN => n14846);
   registers_reg_21_16_inst : DFF_X1 port map( D => n9024, CK => clk, Q => 
                           net271429, QN => n12257);
   registers_reg_22_16_inst : DFF_X1 port map( D => n9023, CK => clk, Q => 
                           registers_22_16_port, QN => n15387);
   registers_reg_23_16_inst : DFF_X1 port map( D => n9022, CK => clk, Q => 
                           registers_23_16_port, QN => n15897);
   registers_reg_24_16_inst : DFF_X1 port map( D => n9021, CK => clk, Q => 
                           net227197, QN => n15195);
   registers_reg_25_16_inst : DFF_X1 port map( D => n9020, CK => clk, Q => 
                           registers_25_16_port, QN => n14314);
   registers_reg_26_16_inst : DFF_X1 port map( D => n9019, CK => clk, Q => 
                           net271428, QN => n14035);
   registers_reg_27_16_inst : DFF_X1 port map( D => n9018, CK => clk, Q => 
                           net271427, QN => n12033);
   registers_reg_28_16_inst : DFF_X1 port map( D => n9017, CK => clk, Q => 
                           net227196, QN => n15018);
   registers_reg_29_16_inst : DFF_X1 port map( D => n9016, CK => clk, Q => 
                           registers_29_16_port, QN => n15830);
   registers_reg_30_16_inst : DFF_X1 port map( D => n9015, CK => clk, Q => 
                           registers_30_16_port, QN => n14692);
   registers_reg_31_16_inst : DFF_X1 port map( D => n9014, CK => clk, Q => 
                           net227195, QN => n15750);
   registers_reg_32_16_inst : DFF_X1 port map( D => n9013, CK => clk, Q => 
                           net271426, QN => n12325);
   registers_reg_33_16_inst : DFF_X1 port map( D => n9012, CK => clk, Q => 
                           net271425, QN => n11858);
   registers_reg_34_16_inst : DFF_X1 port map( D => n9011, CK => clk, Q => 
                           registers_34_16_port, QN => n15510);
   registers_reg_35_16_inst : DFF_X1 port map( D => n9010, CK => clk, Q => 
                           net227194, QN => n15609);
   registers_reg_36_16_inst : DFF_X1 port map( D => n9009, CK => clk, Q => 
                           registers_36_16_port, QN => n15167);
   registers_reg_37_16_inst : DFF_X1 port map( D => n9008, CK => clk, Q => 
                           registers_37_16_port, QN => n14391);
   registers_reg_38_16_inst : DFF_X1 port map( D => n9007, CK => clk, Q => 
                           registers_38_16_port, QN => n15051);
   registers_reg_39_16_inst : DFF_X1 port map( D => n9006, CK => clk, Q => 
                           net271424, QN => n12187);
   registers_reg_40_16_inst : DFF_X1 port map( D => n9005, CK => clk, Q => 
                           registers_40_16_port, QN => n15102);
   registers_reg_41_16_inst : DFF_X1 port map( D => n9004, CK => clk, Q => 
                           registers_41_16_port, QN => n14456);
   registers_reg_42_16_inst : DFF_X1 port map( D => n9003, CK => clk, Q => 
                           registers_42_16_port, QN => n15935);
   registers_reg_43_16_inst : DFF_X1 port map( D => n9002, CK => clk, Q => 
                           registers_43_16_port, QN => n14902);
   registers_reg_44_16_inst : DFF_X1 port map( D => n9001, CK => clk, Q => 
                           registers_44_16_port, QN => n15480);
   registers_reg_45_16_inst : DFF_X1 port map( D => n9000, CK => clk, Q => 
                           registers_45_16_port, QN => n14802);
   registers_reg_46_16_inst : DFF_X1 port map( D => n8999, CK => clk, Q => 
                           net227193, QN => n12008);
   registers_reg_47_16_inst : DFF_X1 port map( D => n8998, CK => clk, Q => 
                           registers_47_16_port, QN => n14561);
   registers_reg_48_16_inst : DFF_X1 port map( D => n8997, CK => clk, Q => 
                           registers_48_16_port, QN => n15566);
   registers_reg_49_16_inst : DFF_X1 port map( D => n8996, CK => clk, Q => 
                           registers_49_16_port, QN => n14498);
   registers_reg_50_16_inst : DFF_X1 port map( D => n8995, CK => clk, Q => 
                           registers_50_16_port, QN => n15984);
   registers_reg_51_16_inst : DFF_X1 port map( D => n8994, CK => clk, Q => 
                           registers_51_16_port, QN => n15413);
   registers_reg_52_16_inst : DFF_X1 port map( D => n8993, CK => clk, Q => 
                           net227192, QN => n14952);
   registers_reg_53_16_inst : DFF_X1 port map( D => n8992, CK => clk, Q => 
                           net227191, QN => n15962);
   registers_reg_54_16_inst : DFF_X1 port map( D => n8991, CK => clk, Q => 
                           registers_54_16_port, QN => n14584);
   registers_reg_55_16_inst : DFF_X1 port map( D => n8990, CK => clk, Q => 
                           registers_55_16_port, QN => n12103);
   registers_reg_56_16_inst : DFF_X1 port map( D => n8989, CK => clk, Q => 
                           registers_56_16_port, QN => n16020);
   registers_reg_57_16_inst : DFF_X1 port map( D => n8988, CK => clk, Q => 
                           net227190, QN => n15256);
   registers_reg_58_16_inst : DFF_X1 port map( D => n8987, CK => clk, Q => 
                           net227189, QN => n14923);
   registers_reg_59_16_inst : DFF_X1 port map( D => n8986, CK => clk, Q => 
                           registers_59_16_port, QN => n15445);
   registers_reg_60_16_inst : DFF_X1 port map( D => n8985, CK => clk, Q => 
                           registers_60_16_port, QN => n14656);
   registers_reg_61_16_inst : DFF_X1 port map( D => n8984, CK => clk, Q => 
                           net227188, QN => n15647);
   registers_reg_62_16_inst : DFF_X1 port map( D => n8983, CK => clk, Q => 
                           registers_62_16_port, QN => n15136);
   registers_reg_63_16_inst : DFF_X1 port map( D => n8982, CK => clk, Q => 
                           registers_63_16_port, QN => n14519);
   to_mem_reg_16_inst : DFF_X1 port map( D => n8981, CK => clk, Q => net271423,
                           QN => n7709);
   registers_reg_64_16_inst : DFF_X1 port map( D => n8980, CK => clk, Q => 
                           net227187, QN => n16158);
   registers_reg_65_16_inst : DFF_X1 port map( D => n8979, CK => clk, Q => 
                           net227186, QN => n16107);
   registers_reg_66_16_inst : DFF_X1 port map( D => n8978, CK => clk, Q => 
                           net227185, QN => n16077);
   registers_reg_67_16_inst : DFF_X1 port map( D => n8977, CK => clk, Q => 
                           net271422, QN => n14255);
   registers_reg_68_16_inst : DFF_X1 port map( D => n8976, CK => clk, Q => 
                           registers_68_16_port, QN => n16195);
   registers_reg_69_16_inst : DFF_X1 port map( D => n8975, CK => clk, Q => 
                           net227184, QN => n16169);
   registers_reg_70_16_inst : DFF_X1 port map( D => n8974, CK => clk, Q => 
                           net227183, QN => n16076);
   registers_reg_0_15_inst : DFF_X1 port map( D => n8973, CK => clk, Q => 
                           registers_0_15_port, QN => n15866);
   registers_reg_1_15_inst : DFF_X1 port map( D => n8972, CK => clk, Q => 
                           registers_1_15_port, QN => n15608);
   registers_reg_2_15_inst : DFF_X1 port map( D => n8971, CK => clk, Q => 
                           registers_2_15_port, QN => n14799);
   registers_reg_3_15_inst : DFF_X1 port map( D => n8970, CK => clk, Q => 
                           net227182, QN => n15773);
   registers_reg_4_15_inst : DFF_X1 port map( D => n8969, CK => clk, Q => 
                           registers_4_15_port, QN => n15536);
   registers_reg_5_15_inst : DFF_X1 port map( D => n8968, CK => clk, Q => 
                           registers_5_15_port, QN => n14740);
   registers_reg_6_15_inst : DFF_X1 port map( D => n8967, CK => clk, Q => 
                           net271421, QN => n14032);
   registers_reg_7_15_inst : DFF_X1 port map( D => n8966, CK => clk, Q => 
                           registers_7_15_port, QN => n15341);
   registers_reg_8_15_inst : DFF_X1 port map( D => n8965, CK => clk, Q => 
                           net227181, QN => n15224);
   registers_reg_9_15_inst : DFF_X1 port map( D => n8964, CK => clk, Q => 
                           registers_9_15_port, QN => n14343);
   registers_reg_10_15_inst : DFF_X1 port map( D => n8963, CK => clk, Q => 
                           registers_10_15_port, QN => n14741);
   registers_reg_11_15_inst : DFF_X1 port map( D => n8962, CK => clk, Q => 
                           registers_11_15_port, QN => n14453);
   registers_reg_12_15_inst : DFF_X1 port map( D => n8961, CK => clk, Q => 
                           registers_12_15_port, QN => n15683);
   registers_reg_13_15_inst : DFF_X1 port map( D => n8960, CK => clk, Q => 
                           net227180, QN => n15099);
   registers_reg_14_15_inst : DFF_X1 port map( D => n8959, CK => clk, Q => 
                           net271420, QN => n11895);
   registers_reg_15_15_inst : DFF_X1 port map( D => n8958, CK => clk, Q => 
                           registers_15_15_port, QN => n15306);
   registers_reg_16_15_inst : DFF_X1 port map( D => n8957, CK => clk, Q => 
                           registers_16_15_port, QN => n15713);
   registers_reg_17_15_inst : DFF_X1 port map( D => n8956, CK => clk, Q => 
                           registers_17_15_port, QN => n14619);
   registers_reg_18_15_inst : DFF_X1 port map( D => n8955, CK => clk, Q => 
                           registers_18_15_port, QN => n14390);
   registers_reg_19_15_inst : DFF_X1 port map( D => n8954, CK => clk, Q => 
                           registers_19_15_port, QN => n15829);
   registers_reg_20_15_inst : DFF_X1 port map( D => n8953, CK => clk, Q => 
                           net271419, QN => n14845);
   registers_reg_21_15_inst : DFF_X1 port map( D => n8952, CK => clk, Q => 
                           net271418, QN => n12256);
   registers_reg_22_15_inst : DFF_X1 port map( D => n8951, CK => clk, Q => 
                           registers_22_15_port, QN => n15386);
   registers_reg_23_15_inst : DFF_X1 port map( D => n8950, CK => clk, Q => 
                           registers_23_15_port, QN => n15896);
   registers_reg_24_15_inst : DFF_X1 port map( D => n8949, CK => clk, Q => 
                           net227179, QN => n15194);
   registers_reg_25_15_inst : DFF_X1 port map( D => n8948, CK => clk, Q => 
                           registers_25_15_port, QN => n14313);
   registers_reg_26_15_inst : DFF_X1 port map( D => n8947, CK => clk, Q => 
                           net271417, QN => n14015);
   registers_reg_27_15_inst : DFF_X1 port map( D => n8946, CK => clk, Q => 
                           net271416, QN => n12032);
   registers_reg_28_15_inst : DFF_X1 port map( D => n8945, CK => clk, Q => 
                           net227178, QN => n15017);
   registers_reg_29_15_inst : DFF_X1 port map( D => n8944, CK => clk, Q => 
                           registers_29_15_port, QN => n15828);
   registers_reg_30_15_inst : DFF_X1 port map( D => n8943, CK => clk, Q => 
                           registers_30_15_port, QN => n14691);
   registers_reg_31_15_inst : DFF_X1 port map( D => n8942, CK => clk, Q => 
                           net227177, QN => n15749);
   registers_reg_32_15_inst : DFF_X1 port map( D => n8941, CK => clk, Q => 
                           net271415, QN => n12324);
   registers_reg_33_15_inst : DFF_X1 port map( D => n8940, CK => clk, Q => 
                           net271414, QN => n11857);
   registers_reg_34_15_inst : DFF_X1 port map( D => n8939, CK => clk, Q => 
                           registers_34_15_port, QN => n15509);
   registers_reg_35_15_inst : DFF_X1 port map( D => n8938, CK => clk, Q => 
                           net227176, QN => n15607);
   registers_reg_36_15_inst : DFF_X1 port map( D => n8937, CK => clk, Q => 
                           registers_36_15_port, QN => n15166);
   registers_reg_37_15_inst : DFF_X1 port map( D => n8936, CK => clk, Q => 
                           registers_37_15_port, QN => n14389);
   registers_reg_38_15_inst : DFF_X1 port map( D => n8935, CK => clk, Q => 
                           registers_38_15_port, QN => n15050);
   registers_reg_39_15_inst : DFF_X1 port map( D => n8934, CK => clk, Q => 
                           net271413, QN => n12186);
   registers_reg_40_15_inst : DFF_X1 port map( D => n8933, CK => clk, Q => 
                           registers_40_15_port, QN => n15100);
   registers_reg_41_15_inst : DFF_X1 port map( D => n8932, CK => clk, Q => 
                           registers_41_15_port, QN => n14454);
   registers_reg_42_15_inst : DFF_X1 port map( D => n8931, CK => clk, Q => 
                           registers_42_15_port, QN => n15934);
   registers_reg_43_15_inst : DFF_X1 port map( D => n8930, CK => clk, Q => 
                           registers_43_15_port, QN => n14901);
   registers_reg_44_15_inst : DFF_X1 port map( D => n8929, CK => clk, Q => 
                           registers_44_15_port, QN => n15479);
   registers_reg_45_15_inst : DFF_X1 port map( D => n8928, CK => clk, Q => 
                           registers_45_15_port, QN => n14800);
   registers_reg_46_15_inst : DFF_X1 port map( D => n8927, CK => clk, Q => 
                           net227175, QN => n12007);
   registers_reg_47_15_inst : DFF_X1 port map( D => n8926, CK => clk, Q => 
                           registers_47_15_port, QN => n14560);
   registers_reg_48_15_inst : DFF_X1 port map( D => n8925, CK => clk, Q => 
                           registers_48_15_port, QN => n15565);
   registers_reg_49_15_inst : DFF_X1 port map( D => n8924, CK => clk, Q => 
                           registers_49_15_port, QN => n14497);
   registers_reg_50_15_inst : DFF_X1 port map( D => n8923, CK => clk, Q => 
                           registers_50_15_port, QN => n15983);
   registers_reg_51_15_inst : DFF_X1 port map( D => n8922, CK => clk, Q => 
                           registers_51_15_port, QN => n15412);
   registers_reg_52_15_inst : DFF_X1 port map( D => n8921, CK => clk, Q => 
                           net227174, QN => n14951);
   registers_reg_53_15_inst : DFF_X1 port map( D => n8920, CK => clk, Q => 
                           net227173, QN => n15961);
   registers_reg_54_15_inst : DFF_X1 port map( D => n8919, CK => clk, Q => 
                           registers_54_15_port, QN => n14583);
   registers_reg_55_15_inst : DFF_X1 port map( D => n8918, CK => clk, Q => 
                           registers_55_15_port, QN => n12102);
   registers_reg_56_15_inst : DFF_X1 port map( D => n8917, CK => clk, Q => 
                           registers_56_15_port, QN => n16019);
   registers_reg_57_15_inst : DFF_X1 port map( D => n8916, CK => clk, Q => 
                           net227172, QN => n15255);
   registers_reg_58_15_inst : DFF_X1 port map( D => n8915, CK => clk, Q => 
                           net227171, QN => n14922);
   registers_reg_59_15_inst : DFF_X1 port map( D => n8914, CK => clk, Q => 
                           registers_59_15_port, QN => n15444);
   registers_reg_60_15_inst : DFF_X1 port map( D => n8913, CK => clk, Q => 
                           registers_60_15_port, QN => n14655);
   registers_reg_61_15_inst : DFF_X1 port map( D => n8912, CK => clk, Q => 
                           net227170, QN => n15646);
   registers_reg_62_15_inst : DFF_X1 port map( D => n8911, CK => clk, Q => 
                           registers_62_15_port, QN => n15135);
   registers_reg_63_15_inst : DFF_X1 port map( D => n8910, CK => clk, Q => 
                           registers_63_15_port, QN => n14518);
   to_mem_reg_15_inst : DFF_X1 port map( D => n8909, CK => clk, Q => net271412,
                           QN => n7710);
   registers_reg_64_15_inst : DFF_X1 port map( D => n8908, CK => clk, Q => 
                           net227169, QN => n16157);
   registers_reg_65_15_inst : DFF_X1 port map( D => n8907, CK => clk, Q => 
                           net227168, QN => n16106);
   registers_reg_66_15_inst : DFF_X1 port map( D => n8906, CK => clk, Q => 
                           net227167, QN => n16075);
   registers_reg_67_15_inst : DFF_X1 port map( D => n8905, CK => clk, Q => 
                           net271411, QN => n14246);
   registers_reg_68_15_inst : DFF_X1 port map( D => n8904, CK => clk, Q => 
                           registers_68_15_port, QN => n16194);
   registers_reg_69_15_inst : DFF_X1 port map( D => n8903, CK => clk, Q => 
                           net227166, QN => n16168);
   registers_reg_70_15_inst : DFF_X1 port map( D => n8902, CK => clk, Q => 
                           net227165, QN => n16074);
   registers_reg_0_14_inst : DFF_X1 port map( D => n8901, CK => clk, Q => 
                           registers_0_14_port, QN => n15865);
   registers_reg_1_14_inst : DFF_X1 port map( D => n8900, CK => clk, Q => 
                           registers_1_14_port, QN => n15606);
   registers_reg_2_14_inst : DFF_X1 port map( D => n8899, CK => clk, Q => 
                           registers_2_14_port, QN => n14797);
   registers_reg_3_14_inst : DFF_X1 port map( D => n8898, CK => clk, Q => 
                           net227164, QN => n15772);
   registers_reg_4_14_inst : DFF_X1 port map( D => n8897, CK => clk, Q => 
                           registers_4_14_port, QN => n15535);
   registers_reg_5_14_inst : DFF_X1 port map( D => n8896, CK => clk, Q => 
                           registers_5_14_port, QN => n14738);
   registers_reg_6_14_inst : DFF_X1 port map( D => n8895, CK => clk, Q => 
                           net271410, QN => n14014);
   registers_reg_7_14_inst : DFF_X1 port map( D => n8894, CK => clk, Q => 
                           registers_7_14_port, QN => n15340);
   registers_reg_8_14_inst : DFF_X1 port map( D => n8893, CK => clk, Q => 
                           net227163, QN => n15223);
   registers_reg_9_14_inst : DFF_X1 port map( D => n8892, CK => clk, Q => 
                           registers_9_14_port, QN => n14342);
   registers_reg_10_14_inst : DFF_X1 port map( D => n8891, CK => clk, Q => 
                           registers_10_14_port, QN => n14739);
   registers_reg_11_14_inst : DFF_X1 port map( D => n8890, CK => clk, Q => 
                           registers_11_14_port, QN => n14451);
   registers_reg_12_14_inst : DFF_X1 port map( D => n8889, CK => clk, Q => 
                           registers_12_14_port, QN => n15682);
   registers_reg_13_14_inst : DFF_X1 port map( D => n8888, CK => clk, Q => 
                           net227162, QN => n15097);
   registers_reg_14_14_inst : DFF_X1 port map( D => n8887, CK => clk, Q => 
                           net271409, QN => n11894);
   registers_reg_15_14_inst : DFF_X1 port map( D => n8886, CK => clk, Q => 
                           registers_15_14_port, QN => n15305);
   registers_reg_16_14_inst : DFF_X1 port map( D => n8885, CK => clk, Q => 
                           registers_16_14_port, QN => n15712);
   registers_reg_17_14_inst : DFF_X1 port map( D => n8884, CK => clk, Q => 
                           registers_17_14_port, QN => n14618);
   registers_reg_18_14_inst : DFF_X1 port map( D => n8883, CK => clk, Q => 
                           registers_18_14_port, QN => n14388);
   registers_reg_19_14_inst : DFF_X1 port map( D => n8882, CK => clk, Q => 
                           registers_19_14_port, QN => n15827);
   registers_reg_20_14_inst : DFF_X1 port map( D => n8881, CK => clk, Q => 
                           net271408, QN => n14844);
   registers_reg_21_14_inst : DFF_X1 port map( D => n8880, CK => clk, Q => 
                           net271407, QN => n12255);
   registers_reg_22_14_inst : DFF_X1 port map( D => n8879, CK => clk, Q => 
                           registers_22_14_port, QN => n15385);
   registers_reg_23_14_inst : DFF_X1 port map( D => n8878, CK => clk, Q => 
                           registers_23_14_port, QN => n15895);
   registers_reg_24_14_inst : DFF_X1 port map( D => n8877, CK => clk, Q => 
                           net227161, QN => n15193);
   registers_reg_25_14_inst : DFF_X1 port map( D => n8876, CK => clk, Q => 
                           registers_25_14_port, QN => n14312);
   registers_reg_26_14_inst : DFF_X1 port map( D => n8875, CK => clk, Q => 
                           net271406, QN => n14008);
   registers_reg_27_14_inst : DFF_X1 port map( D => n8874, CK => clk, Q => 
                           net271405, QN => n12031);
   registers_reg_28_14_inst : DFF_X1 port map( D => n8873, CK => clk, Q => 
                           net227160, QN => n15016);
   registers_reg_29_14_inst : DFF_X1 port map( D => n8872, CK => clk, Q => 
                           registers_29_14_port, QN => n15826);
   registers_reg_30_14_inst : DFF_X1 port map( D => n8871, CK => clk, Q => 
                           registers_30_14_port, QN => n14690);
   registers_reg_31_14_inst : DFF_X1 port map( D => n8870, CK => clk, Q => 
                           net227159, QN => n15748);
   registers_reg_32_14_inst : DFF_X1 port map( D => n8869, CK => clk, Q => 
                           net271404, QN => n12323);
   registers_reg_33_14_inst : DFF_X1 port map( D => n8868, CK => clk, Q => 
                           net271403, QN => n11856);
   registers_reg_34_14_inst : DFF_X1 port map( D => n8867, CK => clk, Q => 
                           registers_34_14_port, QN => n15508);
   registers_reg_35_14_inst : DFF_X1 port map( D => n8866, CK => clk, Q => 
                           net227158, QN => n15605);
   registers_reg_36_14_inst : DFF_X1 port map( D => n8865, CK => clk, Q => 
                           registers_36_14_port, QN => n15165);
   registers_reg_37_14_inst : DFF_X1 port map( D => n8864, CK => clk, Q => 
                           registers_37_14_port, QN => n14387);
   registers_reg_38_14_inst : DFF_X1 port map( D => n8863, CK => clk, Q => 
                           registers_38_14_port, QN => n15049);
   registers_reg_39_14_inst : DFF_X1 port map( D => n8862, CK => clk, Q => 
                           net271402, QN => n12185);
   registers_reg_40_14_inst : DFF_X1 port map( D => n8861, CK => clk, Q => 
                           registers_40_14_port, QN => n15098);
   registers_reg_41_14_inst : DFF_X1 port map( D => n8860, CK => clk, Q => 
                           registers_41_14_port, QN => n14452);
   registers_reg_42_14_inst : DFF_X1 port map( D => n8859, CK => clk, Q => 
                           registers_42_14_port, QN => n15933);
   registers_reg_43_14_inst : DFF_X1 port map( D => n8858, CK => clk, Q => 
                           registers_43_14_port, QN => n14900);
   registers_reg_44_14_inst : DFF_X1 port map( D => n8857, CK => clk, Q => 
                           registers_44_14_port, QN => n15478);
   registers_reg_45_14_inst : DFF_X1 port map( D => n8856, CK => clk, Q => 
                           registers_45_14_port, QN => n14798);
   registers_reg_46_14_inst : DFF_X1 port map( D => n8855, CK => clk, Q => 
                           net227157, QN => n12006);
   registers_reg_47_14_inst : DFF_X1 port map( D => n8854, CK => clk, Q => 
                           registers_47_14_port, QN => n14559);
   registers_reg_48_14_inst : DFF_X1 port map( D => n8853, CK => clk, Q => 
                           registers_48_14_port, QN => n15564);
   registers_reg_49_14_inst : DFF_X1 port map( D => n8852, CK => clk, Q => 
                           registers_49_14_port, QN => n14496);
   registers_reg_50_14_inst : DFF_X1 port map( D => n8851, CK => clk, Q => 
                           registers_50_14_port, QN => n15982);
   registers_reg_51_14_inst : DFF_X1 port map( D => n8850, CK => clk, Q => 
                           registers_51_14_port, QN => n15411);
   registers_reg_52_14_inst : DFF_X1 port map( D => n8849, CK => clk, Q => 
                           net227156, QN => n14950);
   registers_reg_53_14_inst : DFF_X1 port map( D => n8848, CK => clk, Q => 
                           net227155, QN => n15960);
   registers_reg_54_14_inst : DFF_X1 port map( D => n8847, CK => clk, Q => 
                           registers_54_14_port, QN => n14582);
   registers_reg_55_14_inst : DFF_X1 port map( D => n8846, CK => clk, Q => 
                           registers_55_14_port, QN => n12101);
   registers_reg_56_14_inst : DFF_X1 port map( D => n8845, CK => clk, Q => 
                           registers_56_14_port, QN => n16018);
   registers_reg_57_14_inst : DFF_X1 port map( D => n8844, CK => clk, Q => 
                           net227154, QN => n15254);
   registers_reg_58_14_inst : DFF_X1 port map( D => n8843, CK => clk, Q => 
                           net227153, QN => n14921);
   registers_reg_59_14_inst : DFF_X1 port map( D => n8842, CK => clk, Q => 
                           registers_59_14_port, QN => n15443);
   registers_reg_60_14_inst : DFF_X1 port map( D => n8841, CK => clk, Q => 
                           registers_60_14_port, QN => n14654);
   registers_reg_61_14_inst : DFF_X1 port map( D => n8840, CK => clk, Q => 
                           net227152, QN => n15645);
   registers_reg_62_14_inst : DFF_X1 port map( D => n8839, CK => clk, Q => 
                           registers_62_14_port, QN => n15134);
   registers_reg_63_14_inst : DFF_X1 port map( D => n8838, CK => clk, Q => 
                           registers_63_14_port, QN => n14517);
   to_mem_reg_14_inst : DFF_X1 port map( D => n8837, CK => clk, Q => net271401,
                           QN => n7711);
   registers_reg_64_14_inst : DFF_X1 port map( D => n8836, CK => clk, Q => 
                           net227151, QN => n16156);
   registers_reg_65_14_inst : DFF_X1 port map( D => n8835, CK => clk, Q => 
                           net227150, QN => n16105);
   registers_reg_66_14_inst : DFF_X1 port map( D => n8834, CK => clk, Q => 
                           net227149, QN => n16073);
   registers_reg_67_14_inst : DFF_X1 port map( D => n8833, CK => clk, Q => 
                           net271400, QN => n14243);
   registers_reg_68_14_inst : DFF_X1 port map( D => n8832, CK => clk, Q => 
                           registers_68_14_port, QN => n16193);
   registers_reg_69_14_inst : DFF_X1 port map( D => n8831, CK => clk, Q => 
                           net227148, QN => n16167);
   registers_reg_70_14_inst : DFF_X1 port map( D => n8830, CK => clk, Q => 
                           net227147, QN => n16072);
   registers_reg_0_13_inst : DFF_X1 port map( D => n8829, CK => clk, Q => 
                           registers_0_13_port, QN => n15864);
   registers_reg_1_13_inst : DFF_X1 port map( D => n8828, CK => clk, Q => 
                           registers_1_13_port, QN => n15604);
   registers_reg_2_13_inst : DFF_X1 port map( D => n8827, CK => clk, Q => 
                           registers_2_13_port, QN => n14795);
   registers_reg_3_13_inst : DFF_X1 port map( D => n8826, CK => clk, Q => 
                           net227146, QN => n15771);
   registers_reg_4_13_inst : DFF_X1 port map( D => n8825, CK => clk, Q => 
                           registers_4_13_port, QN => n15534);
   registers_reg_5_13_inst : DFF_X1 port map( D => n8824, CK => clk, Q => 
                           registers_5_13_port, QN => n14736);
   registers_reg_6_13_inst : DFF_X1 port map( D => n8823, CK => clk, Q => 
                           net271399, QN => n13999);
   registers_reg_7_13_inst : DFF_X1 port map( D => n8822, CK => clk, Q => 
                           registers_7_13_port, QN => n15339);
   registers_reg_8_13_inst : DFF_X1 port map( D => n8821, CK => clk, Q => 
                           net227145, QN => n15222);
   registers_reg_9_13_inst : DFF_X1 port map( D => n8820, CK => clk, Q => 
                           registers_9_13_port, QN => n14341);
   registers_reg_10_13_inst : DFF_X1 port map( D => n8819, CK => clk, Q => 
                           registers_10_13_port, QN => n14737);
   registers_reg_11_13_inst : DFF_X1 port map( D => n8818, CK => clk, Q => 
                           registers_11_13_port, QN => n14449);
   registers_reg_12_13_inst : DFF_X1 port map( D => n8817, CK => clk, Q => 
                           registers_12_13_port, QN => n15681);
   registers_reg_13_13_inst : DFF_X1 port map( D => n8816, CK => clk, Q => 
                           net227144, QN => n15095);
   registers_reg_14_13_inst : DFF_X1 port map( D => n8815, CK => clk, Q => 
                           net271398, QN => n11893);
   registers_reg_15_13_inst : DFF_X1 port map( D => n8814, CK => clk, Q => 
                           registers_15_13_port, QN => n15304);
   registers_reg_16_13_inst : DFF_X1 port map( D => n8813, CK => clk, Q => 
                           registers_16_13_port, QN => n15711);
   registers_reg_17_13_inst : DFF_X1 port map( D => n8812, CK => clk, Q => 
                           registers_17_13_port, QN => n14617);
   registers_reg_18_13_inst : DFF_X1 port map( D => n8811, CK => clk, Q => 
                           registers_18_13_port, QN => n14386);
   registers_reg_19_13_inst : DFF_X1 port map( D => n8810, CK => clk, Q => 
                           registers_19_13_port, QN => n15825);
   registers_reg_20_13_inst : DFF_X1 port map( D => n8809, CK => clk, Q => 
                           net271397, QN => n14843);
   registers_reg_21_13_inst : DFF_X1 port map( D => n8808, CK => clk, Q => 
                           net271396, QN => n12254);
   registers_reg_22_13_inst : DFF_X1 port map( D => n8807, CK => clk, Q => 
                           registers_22_13_port, QN => n15384);
   registers_reg_23_13_inst : DFF_X1 port map( D => n8806, CK => clk, Q => 
                           registers_23_13_port, QN => n15894);
   registers_reg_24_13_inst : DFF_X1 port map( D => n8805, CK => clk, Q => 
                           net227143, QN => n15192);
   registers_reg_25_13_inst : DFF_X1 port map( D => n8804, CK => clk, Q => 
                           registers_25_13_port, QN => n14311);
   registers_reg_26_13_inst : DFF_X1 port map( D => n8803, CK => clk, Q => 
                           net271395, QN => n13996);
   registers_reg_27_13_inst : DFF_X1 port map( D => n8802, CK => clk, Q => 
                           net271394, QN => n12030);
   registers_reg_28_13_inst : DFF_X1 port map( D => n8801, CK => clk, Q => 
                           net227142, QN => n15015);
   registers_reg_29_13_inst : DFF_X1 port map( D => n8800, CK => clk, Q => 
                           registers_29_13_port, QN => n15824);
   registers_reg_30_13_inst : DFF_X1 port map( D => n8799, CK => clk, Q => 
                           registers_30_13_port, QN => n14689);
   registers_reg_31_13_inst : DFF_X1 port map( D => n8798, CK => clk, Q => 
                           net227141, QN => n15747);
   registers_reg_32_13_inst : DFF_X1 port map( D => n8797, CK => clk, Q => 
                           net271393, QN => n12322);
   registers_reg_33_13_inst : DFF_X1 port map( D => n8796, CK => clk, Q => 
                           net271392, QN => n11855);
   registers_reg_34_13_inst : DFF_X1 port map( D => n8795, CK => clk, Q => 
                           registers_34_13_port, QN => n15507);
   registers_reg_35_13_inst : DFF_X1 port map( D => n8794, CK => clk, Q => 
                           net227140, QN => n15603);
   registers_reg_36_13_inst : DFF_X1 port map( D => n8793, CK => clk, Q => 
                           registers_36_13_port, QN => n15164);
   registers_reg_37_13_inst : DFF_X1 port map( D => n8792, CK => clk, Q => 
                           registers_37_13_port, QN => n14385);
   registers_reg_38_13_inst : DFF_X1 port map( D => n8791, CK => clk, Q => 
                           registers_38_13_port, QN => n15048);
   registers_reg_39_13_inst : DFF_X1 port map( D => n8790, CK => clk, Q => 
                           net271391, QN => n12183);
   registers_reg_40_13_inst : DFF_X1 port map( D => n8789, CK => clk, Q => 
                           registers_40_13_port, QN => n15096);
   registers_reg_41_13_inst : DFF_X1 port map( D => n8788, CK => clk, Q => 
                           registers_41_13_port, QN => n14450);
   registers_reg_42_13_inst : DFF_X1 port map( D => n8787, CK => clk, Q => 
                           registers_42_13_port, QN => n15932);
   registers_reg_43_13_inst : DFF_X1 port map( D => n8786, CK => clk, Q => 
                           registers_43_13_port, QN => n14899);
   registers_reg_44_13_inst : DFF_X1 port map( D => n8785, CK => clk, Q => 
                           registers_44_13_port, QN => n15477);
   registers_reg_45_13_inst : DFF_X1 port map( D => n8784, CK => clk, Q => 
                           registers_45_13_port, QN => n14796);
   registers_reg_46_13_inst : DFF_X1 port map( D => n8783, CK => clk, Q => 
                           net227139, QN => n12005);
   registers_reg_47_13_inst : DFF_X1 port map( D => n8782, CK => clk, Q => 
                           registers_47_13_port, QN => n14558);
   registers_reg_48_13_inst : DFF_X1 port map( D => n8781, CK => clk, Q => 
                           registers_48_13_port, QN => n15563);
   registers_reg_49_13_inst : DFF_X1 port map( D => n8780, CK => clk, Q => 
                           registers_49_13_port, QN => n14495);
   registers_reg_50_13_inst : DFF_X1 port map( D => n8779, CK => clk, Q => 
                           registers_50_13_port, QN => n15981);
   registers_reg_51_13_inst : DFF_X1 port map( D => n8778, CK => clk, Q => 
                           registers_51_13_port, QN => n15410);
   registers_reg_52_13_inst : DFF_X1 port map( D => n8777, CK => clk, Q => 
                           net227138, QN => n14949);
   registers_reg_53_13_inst : DFF_X1 port map( D => n8776, CK => clk, Q => 
                           net227137, QN => n15959);
   registers_reg_54_13_inst : DFF_X1 port map( D => n8775, CK => clk, Q => 
                           registers_54_13_port, QN => n14581);
   registers_reg_55_13_inst : DFF_X1 port map( D => n8774, CK => clk, Q => 
                           registers_55_13_port, QN => n12100);
   registers_reg_56_13_inst : DFF_X1 port map( D => n8773, CK => clk, Q => 
                           registers_56_13_port, QN => n16017);
   registers_reg_57_13_inst : DFF_X1 port map( D => n8772, CK => clk, Q => 
                           net227136, QN => n15253);
   registers_reg_58_13_inst : DFF_X1 port map( D => n8771, CK => clk, Q => 
                           net227135, QN => n14920);
   registers_reg_59_13_inst : DFF_X1 port map( D => n8770, CK => clk, Q => 
                           registers_59_13_port, QN => n15442);
   registers_reg_60_13_inst : DFF_X1 port map( D => n8769, CK => clk, Q => 
                           registers_60_13_port, QN => n14653);
   registers_reg_61_13_inst : DFF_X1 port map( D => n8768, CK => clk, Q => 
                           net227134, QN => n15644);
   registers_reg_62_13_inst : DFF_X1 port map( D => n8767, CK => clk, Q => 
                           registers_62_13_port, QN => n15133);
   registers_reg_63_13_inst : DFF_X1 port map( D => n8766, CK => clk, Q => 
                           registers_63_13_port, QN => n14516);
   to_mem_reg_13_inst : DFF_X1 port map( D => n8765, CK => clk, Q => net271390,
                           QN => n7712);
   registers_reg_64_13_inst : DFF_X1 port map( D => n8764, CK => clk, Q => 
                           net227133, QN => n16155);
   registers_reg_65_13_inst : DFF_X1 port map( D => n8763, CK => clk, Q => 
                           net227132, QN => n16104);
   registers_reg_66_13_inst : DFF_X1 port map( D => n8762, CK => clk, Q => 
                           net227131, QN => n16071);
   registers_reg_67_13_inst : DFF_X1 port map( D => n8761, CK => clk, Q => 
                           net271389, QN => n14242);
   registers_reg_68_13_inst : DFF_X1 port map( D => n8760, CK => clk, Q => 
                           registers_68_13_port, QN => n16192);
   registers_reg_69_13_inst : DFF_X1 port map( D => n8759, CK => clk, Q => 
                           net227130, QN => n16166);
   registers_reg_70_13_inst : DFF_X1 port map( D => n8758, CK => clk, Q => 
                           net227129, QN => n16070);
   registers_reg_0_12_inst : DFF_X1 port map( D => n8757, CK => clk, Q => 
                           registers_0_12_port, QN => n15863);
   registers_reg_1_12_inst : DFF_X1 port map( D => n8756, CK => clk, Q => 
                           registers_1_12_port, QN => n15602);
   registers_reg_2_12_inst : DFF_X1 port map( D => n8755, CK => clk, Q => 
                           registers_2_12_port, QN => n14793);
   registers_reg_3_12_inst : DFF_X1 port map( D => n8754, CK => clk, Q => 
                           net227128, QN => n15770);
   registers_reg_4_12_inst : DFF_X1 port map( D => n8753, CK => clk, Q => 
                           registers_4_12_port, QN => n15533);
   registers_reg_5_12_inst : DFF_X1 port map( D => n8752, CK => clk, Q => 
                           registers_5_12_port, QN => n14734);
   registers_reg_6_12_inst : DFF_X1 port map( D => n8751, CK => clk, Q => 
                           net271388, QN => n12669);
   registers_reg_7_12_inst : DFF_X1 port map( D => n8750, CK => clk, Q => 
                           registers_7_12_port, QN => n15338);
   registers_reg_8_12_inst : DFF_X1 port map( D => n8749, CK => clk, Q => 
                           net227127, QN => n15221);
   registers_reg_9_12_inst : DFF_X1 port map( D => n8748, CK => clk, Q => 
                           registers_9_12_port, QN => n14340);
   registers_reg_10_12_inst : DFF_X1 port map( D => n8747, CK => clk, Q => 
                           registers_10_12_port, QN => n14735);
   registers_reg_11_12_inst : DFF_X1 port map( D => n8746, CK => clk, Q => 
                           registers_11_12_port, QN => n14447);
   registers_reg_12_12_inst : DFF_X1 port map( D => n8745, CK => clk, Q => 
                           registers_12_12_port, QN => n15680);
   registers_reg_13_12_inst : DFF_X1 port map( D => n8744, CK => clk, Q => 
                           net227126, QN => n15093);
   registers_reg_14_12_inst : DFF_X1 port map( D => n8743, CK => clk, Q => 
                           net271387, QN => n11892);
   registers_reg_15_12_inst : DFF_X1 port map( D => n8742, CK => clk, Q => 
                           registers_15_12_port, QN => n15303);
   registers_reg_16_12_inst : DFF_X1 port map( D => n8741, CK => clk, Q => 
                           registers_16_12_port, QN => n15710);
   registers_reg_17_12_inst : DFF_X1 port map( D => n8740, CK => clk, Q => 
                           registers_17_12_port, QN => n14616);
   registers_reg_18_12_inst : DFF_X1 port map( D => n8739, CK => clk, Q => 
                           registers_18_12_port, QN => n14384);
   registers_reg_19_12_inst : DFF_X1 port map( D => n8738, CK => clk, Q => 
                           registers_19_12_port, QN => n15823);
   registers_reg_20_12_inst : DFF_X1 port map( D => n8737, CK => clk, Q => 
                           net271386, QN => n14842);
   registers_reg_21_12_inst : DFF_X1 port map( D => n8736, CK => clk, Q => 
                           net271385, QN => n12253);
   registers_reg_22_12_inst : DFF_X1 port map( D => n8735, CK => clk, Q => 
                           registers_22_12_port, QN => n15383);
   registers_reg_23_12_inst : DFF_X1 port map( D => n8734, CK => clk, Q => 
                           registers_23_12_port, QN => n15893);
   registers_reg_24_12_inst : DFF_X1 port map( D => n8733, CK => clk, Q => 
                           net227125, QN => n15191);
   registers_reg_25_12_inst : DFF_X1 port map( D => n8732, CK => clk, Q => 
                           registers_25_12_port, QN => n14310);
   registers_reg_26_12_inst : DFF_X1 port map( D => n8731, CK => clk, Q => 
                           net271384, QN => n12652);
   registers_reg_27_12_inst : DFF_X1 port map( D => n8730, CK => clk, Q => 
                           net271383, QN => n12028);
   registers_reg_28_12_inst : DFF_X1 port map( D => n8729, CK => clk, Q => 
                           net227124, QN => n15014);
   registers_reg_29_12_inst : DFF_X1 port map( D => n8728, CK => clk, Q => 
                           registers_29_12_port, QN => n15822);
   registers_reg_30_12_inst : DFF_X1 port map( D => n8727, CK => clk, Q => 
                           registers_30_12_port, QN => n14688);
   registers_reg_31_12_inst : DFF_X1 port map( D => n8726, CK => clk, Q => 
                           net227123, QN => n15746);
   registers_reg_32_12_inst : DFF_X1 port map( D => n8725, CK => clk, Q => 
                           net271382, QN => n12321);
   registers_reg_33_12_inst : DFF_X1 port map( D => n8724, CK => clk, Q => 
                           net271381, QN => n11854);
   registers_reg_34_12_inst : DFF_X1 port map( D => n8723, CK => clk, Q => 
                           registers_34_12_port, QN => n15506);
   registers_reg_35_12_inst : DFF_X1 port map( D => n8722, CK => clk, Q => 
                           net227122, QN => n15601);
   registers_reg_36_12_inst : DFF_X1 port map( D => n8721, CK => clk, Q => 
                           registers_36_12_port, QN => n15163);
   registers_reg_37_12_inst : DFF_X1 port map( D => n8720, CK => clk, Q => 
                           registers_37_12_port, QN => n14383);
   registers_reg_38_12_inst : DFF_X1 port map( D => n8719, CK => clk, Q => 
                           registers_38_12_port, QN => n15047);
   registers_reg_39_12_inst : DFF_X1 port map( D => n8718, CK => clk, Q => 
                           net271380, QN => n12182);
   registers_reg_40_12_inst : DFF_X1 port map( D => n8717, CK => clk, Q => 
                           registers_40_12_port, QN => n15094);
   registers_reg_41_12_inst : DFF_X1 port map( D => n8716, CK => clk, Q => 
                           registers_41_12_port, QN => n14448);
   registers_reg_42_12_inst : DFF_X1 port map( D => n8715, CK => clk, Q => 
                           registers_42_12_port, QN => n15931);
   registers_reg_43_12_inst : DFF_X1 port map( D => n8714, CK => clk, Q => 
                           registers_43_12_port, QN => n14898);
   registers_reg_44_12_inst : DFF_X1 port map( D => n8713, CK => clk, Q => 
                           registers_44_12_port, QN => n15476);
   registers_reg_45_12_inst : DFF_X1 port map( D => n8712, CK => clk, Q => 
                           registers_45_12_port, QN => n14794);
   registers_reg_46_12_inst : DFF_X1 port map( D => n8711, CK => clk, Q => 
                           net227121, QN => n12004);
   registers_reg_47_12_inst : DFF_X1 port map( D => n8710, CK => clk, Q => 
                           registers_47_12_port, QN => n14557);
   registers_reg_48_12_inst : DFF_X1 port map( D => n8709, CK => clk, Q => 
                           registers_48_12_port, QN => n15562);
   registers_reg_49_12_inst : DFF_X1 port map( D => n8708, CK => clk, Q => 
                           registers_49_12_port, QN => n14494);
   registers_reg_50_12_inst : DFF_X1 port map( D => n8707, CK => clk, Q => 
                           registers_50_12_port, QN => n15980);
   registers_reg_51_12_inst : DFF_X1 port map( D => n8706, CK => clk, Q => 
                           registers_51_12_port, QN => n15409);
   registers_reg_52_12_inst : DFF_X1 port map( D => n8705, CK => clk, Q => 
                           net227120, QN => n14948);
   registers_reg_53_12_inst : DFF_X1 port map( D => n8704, CK => clk, Q => 
                           net227119, QN => n15958);
   registers_reg_54_12_inst : DFF_X1 port map( D => n8703, CK => clk, Q => 
                           registers_54_12_port, QN => n14580);
   registers_reg_55_12_inst : DFF_X1 port map( D => n8702, CK => clk, Q => 
                           registers_55_12_port, QN => n12099);
   registers_reg_56_12_inst : DFF_X1 port map( D => n8701, CK => clk, Q => 
                           registers_56_12_port, QN => n16016);
   registers_reg_57_12_inst : DFF_X1 port map( D => n8700, CK => clk, Q => 
                           net227118, QN => n15252);
   registers_reg_58_12_inst : DFF_X1 port map( D => n8699, CK => clk, Q => 
                           net227117, QN => n14919);
   registers_reg_59_12_inst : DFF_X1 port map( D => n8698, CK => clk, Q => 
                           registers_59_12_port, QN => n15441);
   registers_reg_60_12_inst : DFF_X1 port map( D => n8697, CK => clk, Q => 
                           registers_60_12_port, QN => n14652);
   registers_reg_61_12_inst : DFF_X1 port map( D => n8696, CK => clk, Q => 
                           net227116, QN => n15643);
   registers_reg_62_12_inst : DFF_X1 port map( D => n8695, CK => clk, Q => 
                           registers_62_12_port, QN => n15132);
   registers_reg_63_12_inst : DFF_X1 port map( D => n8694, CK => clk, Q => 
                           registers_63_12_port, QN => n14515);
   to_mem_reg_12_inst : DFF_X1 port map( D => n8693, CK => clk, Q => net271379,
                           QN => n7713);
   registers_reg_64_12_inst : DFF_X1 port map( D => n8692, CK => clk, Q => 
                           net227115, QN => n16154);
   registers_reg_65_12_inst : DFF_X1 port map( D => n8691, CK => clk, Q => 
                           net227114, QN => n16103);
   registers_reg_66_12_inst : DFF_X1 port map( D => n8690, CK => clk, Q => 
                           net227113, QN => n16069);
   registers_reg_67_12_inst : DFF_X1 port map( D => n8689, CK => clk, Q => 
                           net271378, QN => n14235);
   registers_reg_68_12_inst : DFF_X1 port map( D => n8688, CK => clk, Q => 
                           registers_68_12_port, QN => n16191);
   registers_reg_69_12_inst : DFF_X1 port map( D => n8687, CK => clk, Q => 
                           net227112, QN => n16165);
   registers_reg_70_12_inst : DFF_X1 port map( D => n8686, CK => clk, Q => 
                           net227111, QN => n16068);
   registers_reg_0_11_inst : DFF_X1 port map( D => n8685, CK => clk, Q => 
                           registers_0_11_port, QN => n15862);
   registers_reg_1_11_inst : DFF_X1 port map( D => n8684, CK => clk, Q => 
                           registers_1_11_port, QN => n15600);
   registers_reg_2_11_inst : DFF_X1 port map( D => n8683, CK => clk, Q => 
                           registers_2_11_port, QN => n14791);
   registers_reg_3_11_inst : DFF_X1 port map( D => n8682, CK => clk, Q => 
                           net227110, QN => n15769);
   registers_reg_4_11_inst : DFF_X1 port map( D => n8681, CK => clk, Q => 
                           registers_4_11_port, QN => n15532);
   registers_reg_5_11_inst : DFF_X1 port map( D => n8680, CK => clk, Q => 
                           registers_5_11_port, QN => n14732);
   registers_reg_6_11_inst : DFF_X1 port map( D => n8679, CK => clk, Q => 
                           net271377, QN => n12602);
   registers_reg_7_11_inst : DFF_X1 port map( D => n8678, CK => clk, Q => 
                           registers_7_11_port, QN => n15337);
   registers_reg_8_11_inst : DFF_X1 port map( D => n8677, CK => clk, Q => 
                           net227109, QN => n15220);
   registers_reg_9_11_inst : DFF_X1 port map( D => n8676, CK => clk, Q => 
                           registers_9_11_port, QN => n14339);
   registers_reg_10_11_inst : DFF_X1 port map( D => n8675, CK => clk, Q => 
                           registers_10_11_port, QN => n14733);
   registers_reg_11_11_inst : DFF_X1 port map( D => n8674, CK => clk, Q => 
                           registers_11_11_port, QN => n14445);
   registers_reg_12_11_inst : DFF_X1 port map( D => n8673, CK => clk, Q => 
                           registers_12_11_port, QN => n15679);
   registers_reg_13_11_inst : DFF_X1 port map( D => n8672, CK => clk, Q => 
                           net227108, QN => n15091);
   registers_reg_14_11_inst : DFF_X1 port map( D => n8671, CK => clk, Q => 
                           net271376, QN => n11891);
   registers_reg_15_11_inst : DFF_X1 port map( D => n8670, CK => clk, Q => 
                           registers_15_11_port, QN => n15302);
   registers_reg_16_11_inst : DFF_X1 port map( D => n8669, CK => clk, Q => 
                           registers_16_11_port, QN => n15709);
   registers_reg_17_11_inst : DFF_X1 port map( D => n8668, CK => clk, Q => 
                           registers_17_11_port, QN => n14615);
   registers_reg_18_11_inst : DFF_X1 port map( D => n8667, CK => clk, Q => 
                           registers_18_11_port, QN => n14382);
   registers_reg_19_11_inst : DFF_X1 port map( D => n8666, CK => clk, Q => 
                           registers_19_11_port, QN => n15821);
   registers_reg_20_11_inst : DFF_X1 port map( D => n8665, CK => clk, Q => 
                           net271375, QN => n14841);
   registers_reg_21_11_inst : DFF_X1 port map( D => n8664, CK => clk, Q => 
                           net271374, QN => n12215);
   registers_reg_22_11_inst : DFF_X1 port map( D => n8663, CK => clk, Q => 
                           registers_22_11_port, QN => n15382);
   registers_reg_23_11_inst : DFF_X1 port map( D => n8662, CK => clk, Q => 
                           registers_23_11_port, QN => n15892);
   registers_reg_24_11_inst : DFF_X1 port map( D => n8661, CK => clk, Q => 
                           net227107, QN => n15190);
   registers_reg_25_11_inst : DFF_X1 port map( D => n8660, CK => clk, Q => 
                           registers_25_11_port, QN => n14309);
   registers_reg_26_11_inst : DFF_X1 port map( D => n8659, CK => clk, Q => 
                           net271373, QN => n12600);
   registers_reg_27_11_inst : DFF_X1 port map( D => n8658, CK => clk, Q => 
                           net271372, QN => n12027);
   registers_reg_28_11_inst : DFF_X1 port map( D => n8657, CK => clk, Q => 
                           net227106, QN => n15013);
   registers_reg_29_11_inst : DFF_X1 port map( D => n8656, CK => clk, Q => 
                           registers_29_11_port, QN => n15820);
   registers_reg_30_11_inst : DFF_X1 port map( D => n8655, CK => clk, Q => 
                           registers_30_11_port, QN => n14687);
   registers_reg_31_11_inst : DFF_X1 port map( D => n8654, CK => clk, Q => 
                           net227105, QN => n15745);
   registers_reg_32_11_inst : DFF_X1 port map( D => n8653, CK => clk, Q => 
                           net271371, QN => n12320);
   registers_reg_33_11_inst : DFF_X1 port map( D => n8652, CK => clk, Q => 
                           net271370, QN => n11852);
   registers_reg_34_11_inst : DFF_X1 port map( D => n8651, CK => clk, Q => 
                           registers_34_11_port, QN => n15505);
   registers_reg_35_11_inst : DFF_X1 port map( D => n8650, CK => clk, Q => 
                           net227104, QN => n15599);
   registers_reg_36_11_inst : DFF_X1 port map( D => n8649, CK => clk, Q => 
                           registers_36_11_port, QN => n15162);
   registers_reg_37_11_inst : DFF_X1 port map( D => n8648, CK => clk, Q => 
                           registers_37_11_port, QN => n14381);
   registers_reg_38_11_inst : DFF_X1 port map( D => n8647, CK => clk, Q => 
                           registers_38_11_port, QN => n15046);
   registers_reg_39_11_inst : DFF_X1 port map( D => n8646, CK => clk, Q => 
                           net271369, QN => n12181);
   registers_reg_40_11_inst : DFF_X1 port map( D => n8645, CK => clk, Q => 
                           registers_40_11_port, QN => n15092);
   registers_reg_41_11_inst : DFF_X1 port map( D => n8644, CK => clk, Q => 
                           registers_41_11_port, QN => n14446);
   registers_reg_42_11_inst : DFF_X1 port map( D => n8643, CK => clk, Q => 
                           registers_42_11_port, QN => n15930);
   registers_reg_43_11_inst : DFF_X1 port map( D => n8642, CK => clk, Q => 
                           registers_43_11_port, QN => n14897);
   registers_reg_44_11_inst : DFF_X1 port map( D => n8641, CK => clk, Q => 
                           registers_44_11_port, QN => n15475);
   registers_reg_45_11_inst : DFF_X1 port map( D => n8640, CK => clk, Q => 
                           registers_45_11_port, QN => n14792);
   registers_reg_46_11_inst : DFF_X1 port map( D => n8639, CK => clk, Q => 
                           net227103, QN => n12003);
   registers_reg_47_11_inst : DFF_X1 port map( D => n8638, CK => clk, Q => 
                           registers_47_11_port, QN => n14556);
   registers_reg_48_11_inst : DFF_X1 port map( D => n8637, CK => clk, Q => 
                           registers_48_11_port, QN => n15561);
   registers_reg_49_11_inst : DFF_X1 port map( D => n8636, CK => clk, Q => 
                           registers_49_11_port, QN => n14493);
   registers_reg_50_11_inst : DFF_X1 port map( D => n8635, CK => clk, Q => 
                           registers_50_11_port, QN => n15979);
   registers_reg_51_11_inst : DFF_X1 port map( D => n8634, CK => clk, Q => 
                           registers_51_11_port, QN => n15408);
   registers_reg_52_11_inst : DFF_X1 port map( D => n8633, CK => clk, Q => 
                           net227102, QN => n14947);
   registers_reg_53_11_inst : DFF_X1 port map( D => n8632, CK => clk, Q => 
                           net227101, QN => n15957);
   registers_reg_54_11_inst : DFF_X1 port map( D => n8631, CK => clk, Q => 
                           registers_54_11_port, QN => n14579);
   registers_reg_55_11_inst : DFF_X1 port map( D => n8630, CK => clk, Q => 
                           registers_55_11_port, QN => n12098);
   registers_reg_56_11_inst : DFF_X1 port map( D => n8629, CK => clk, Q => 
                           registers_56_11_port, QN => n16015);
   registers_reg_57_11_inst : DFF_X1 port map( D => n8628, CK => clk, Q => 
                           net227100, QN => n15251);
   registers_reg_58_11_inst : DFF_X1 port map( D => n8627, CK => clk, Q => 
                           net227099, QN => n14918);
   registers_reg_59_11_inst : DFF_X1 port map( D => n8626, CK => clk, Q => 
                           registers_59_11_port, QN => n15440);
   registers_reg_60_11_inst : DFF_X1 port map( D => n8625, CK => clk, Q => 
                           registers_60_11_port, QN => n14651);
   registers_reg_61_11_inst : DFF_X1 port map( D => n8624, CK => clk, Q => 
                           net227098, QN => n15642);
   registers_reg_62_11_inst : DFF_X1 port map( D => n8623, CK => clk, Q => 
                           registers_62_11_port, QN => n15131);
   registers_reg_63_11_inst : DFF_X1 port map( D => n8622, CK => clk, Q => 
                           registers_63_11_port, QN => n14514);
   to_mem_reg_11_inst : DFF_X1 port map( D => n8621, CK => clk, Q => net271368,
                           QN => n7714);
   registers_reg_64_11_inst : DFF_X1 port map( D => n8620, CK => clk, Q => 
                           net227097, QN => n16153);
   registers_reg_65_11_inst : DFF_X1 port map( D => n8619, CK => clk, Q => 
                           net227096, QN => n16102);
   registers_reg_66_11_inst : DFF_X1 port map( D => n8618, CK => clk, Q => 
                           net227095, QN => n16067);
   registers_reg_67_11_inst : DFF_X1 port map( D => n8617, CK => clk, Q => 
                           net271367, QN => n14230);
   registers_reg_68_11_inst : DFF_X1 port map( D => n8616, CK => clk, Q => 
                           registers_68_11_port, QN => n16190);
   registers_reg_69_11_inst : DFF_X1 port map( D => n8615, CK => clk, Q => 
                           net227094, QN => n16164);
   registers_reg_70_11_inst : DFF_X1 port map( D => n8614, CK => clk, Q => 
                           net227093, QN => n16066);
   registers_reg_0_10_inst : DFF_X1 port map( D => n8613, CK => clk, Q => 
                           registers_0_10_port, QN => n15861);
   registers_reg_1_10_inst : DFF_X1 port map( D => n8612, CK => clk, Q => 
                           registers_1_10_port, QN => n15598);
   registers_reg_2_10_inst : DFF_X1 port map( D => n8611, CK => clk, Q => 
                           registers_2_10_port, QN => n14789);
   registers_reg_3_10_inst : DFF_X1 port map( D => n8610, CK => clk, Q => 
                           net227092, QN => n15768);
   registers_reg_4_10_inst : DFF_X1 port map( D => n8609, CK => clk, Q => 
                           registers_4_10_port, QN => n15531);
   registers_reg_5_10_inst : DFF_X1 port map( D => n8608, CK => clk, Q => 
                           registers_5_10_port, QN => n14730);
   registers_reg_6_10_inst : DFF_X1 port map( D => n8607, CK => clk, Q => 
                           net271366, QN => n12551);
   registers_reg_7_10_inst : DFF_X1 port map( D => n8606, CK => clk, Q => 
                           registers_7_10_port, QN => n15336);
   registers_reg_8_10_inst : DFF_X1 port map( D => n8605, CK => clk, Q => 
                           net227091, QN => n15219);
   registers_reg_9_10_inst : DFF_X1 port map( D => n8604, CK => clk, Q => 
                           registers_9_10_port, QN => n14338);
   registers_reg_10_10_inst : DFF_X1 port map( D => n8603, CK => clk, Q => 
                           registers_10_10_port, QN => n14731);
   registers_reg_11_10_inst : DFF_X1 port map( D => n8602, CK => clk, Q => 
                           registers_11_10_port, QN => n14443);
   registers_reg_12_10_inst : DFF_X1 port map( D => n8601, CK => clk, Q => 
                           registers_12_10_port, QN => n15678);
   registers_reg_13_10_inst : DFF_X1 port map( D => n8600, CK => clk, Q => 
                           net227090, QN => n15089);
   registers_reg_14_10_inst : DFF_X1 port map( D => n8599, CK => clk, Q => 
                           net271365, QN => n11890);
   registers_reg_15_10_inst : DFF_X1 port map( D => n8598, CK => clk, Q => 
                           registers_15_10_port, QN => n15301);
   registers_reg_16_10_inst : DFF_X1 port map( D => n8597, CK => clk, Q => 
                           registers_16_10_port, QN => n15708);
   registers_reg_17_10_inst : DFF_X1 port map( D => n8596, CK => clk, Q => 
                           registers_17_10_port, QN => n14614);
   registers_reg_18_10_inst : DFF_X1 port map( D => n8595, CK => clk, Q => 
                           registers_18_10_port, QN => n14380);
   registers_reg_19_10_inst : DFF_X1 port map( D => n8594, CK => clk, Q => 
                           registers_19_10_port, QN => n15819);
   registers_reg_20_10_inst : DFF_X1 port map( D => n8593, CK => clk, Q => 
                           net271364, QN => n14840);
   registers_reg_21_10_inst : DFF_X1 port map( D => n8592, CK => clk, Q => 
                           net271363, QN => n12214);
   registers_reg_22_10_inst : DFF_X1 port map( D => n8591, CK => clk, Q => 
                           registers_22_10_port, QN => n15381);
   registers_reg_23_10_inst : DFF_X1 port map( D => n8590, CK => clk, Q => 
                           registers_23_10_port, QN => n15891);
   registers_reg_24_10_inst : DFF_X1 port map( D => n8589, CK => clk, Q => 
                           net227089, QN => n15189);
   registers_reg_25_10_inst : DFF_X1 port map( D => n8588, CK => clk, Q => 
                           registers_25_10_port, QN => n14308);
   registers_reg_26_10_inst : DFF_X1 port map( D => n8587, CK => clk, Q => 
                           net271362, QN => n12411);
   registers_reg_27_10_inst : DFF_X1 port map( D => n8586, CK => clk, Q => 
                           net271361, QN => n12026);
   registers_reg_28_10_inst : DFF_X1 port map( D => n8585, CK => clk, Q => 
                           net227088, QN => n15012);
   registers_reg_29_10_inst : DFF_X1 port map( D => n8584, CK => clk, Q => 
                           registers_29_10_port, QN => n15818);
   registers_reg_30_10_inst : DFF_X1 port map( D => n8583, CK => clk, Q => 
                           registers_30_10_port, QN => n14686);
   registers_reg_31_10_inst : DFF_X1 port map( D => n8582, CK => clk, Q => 
                           net227087, QN => n15744);
   registers_reg_32_10_inst : DFF_X1 port map( D => n8581, CK => clk, Q => 
                           net271360, QN => n12319);
   registers_reg_33_10_inst : DFF_X1 port map( D => n8580, CK => clk, Q => 
                           net271359, QN => n11851);
   registers_reg_34_10_inst : DFF_X1 port map( D => n8579, CK => clk, Q => 
                           registers_34_10_port, QN => n15504);
   registers_reg_35_10_inst : DFF_X1 port map( D => n8578, CK => clk, Q => 
                           net227086, QN => n15597);
   registers_reg_36_10_inst : DFF_X1 port map( D => n8577, CK => clk, Q => 
                           registers_36_10_port, QN => n15161);
   registers_reg_37_10_inst : DFF_X1 port map( D => n8576, CK => clk, Q => 
                           registers_37_10_port, QN => n14379);
   registers_reg_38_10_inst : DFF_X1 port map( D => n8575, CK => clk, Q => 
                           registers_38_10_port, QN => n15045);
   registers_reg_39_10_inst : DFF_X1 port map( D => n8574, CK => clk, Q => 
                           net271358, QN => n12180);
   registers_reg_40_10_inst : DFF_X1 port map( D => n8573, CK => clk, Q => 
                           registers_40_10_port, QN => n15090);
   registers_reg_41_10_inst : DFF_X1 port map( D => n8572, CK => clk, Q => 
                           registers_41_10_port, QN => n14444);
   registers_reg_42_10_inst : DFF_X1 port map( D => n8571, CK => clk, Q => 
                           registers_42_10_port, QN => n15929);
   registers_reg_43_10_inst : DFF_X1 port map( D => n8570, CK => clk, Q => 
                           registers_43_10_port, QN => n14896);
   registers_reg_44_10_inst : DFF_X1 port map( D => n8569, CK => clk, Q => 
                           registers_44_10_port, QN => n15474);
   registers_reg_45_10_inst : DFF_X1 port map( D => n8568, CK => clk, Q => 
                           registers_45_10_port, QN => n14790);
   registers_reg_46_10_inst : DFF_X1 port map( D => n8567, CK => clk, Q => 
                           net227085, QN => n12002);
   registers_reg_47_10_inst : DFF_X1 port map( D => n8566, CK => clk, Q => 
                           registers_47_10_port, QN => n14555);
   registers_reg_48_10_inst : DFF_X1 port map( D => n8565, CK => clk, Q => 
                           registers_48_10_port, QN => n15560);
   registers_reg_49_10_inst : DFF_X1 port map( D => n8564, CK => clk, Q => 
                           registers_49_10_port, QN => n14492);
   registers_reg_50_10_inst : DFF_X1 port map( D => n8563, CK => clk, Q => 
                           registers_50_10_port, QN => n15978);
   registers_reg_51_10_inst : DFF_X1 port map( D => n8562, CK => clk, Q => 
                           registers_51_10_port, QN => n15407);
   registers_reg_52_10_inst : DFF_X1 port map( D => n8561, CK => clk, Q => 
                           net227084, QN => n14946);
   registers_reg_53_10_inst : DFF_X1 port map( D => n8560, CK => clk, Q => 
                           net227083, QN => n15956);
   registers_reg_54_10_inst : DFF_X1 port map( D => n8559, CK => clk, Q => 
                           registers_54_10_port, QN => n14578);
   registers_reg_55_10_inst : DFF_X1 port map( D => n8558, CK => clk, Q => 
                           registers_55_10_port, QN => n12060);
   registers_reg_56_10_inst : DFF_X1 port map( D => n8557, CK => clk, Q => 
                           registers_56_10_port, QN => n16014);
   registers_reg_57_10_inst : DFF_X1 port map( D => n8556, CK => clk, Q => 
                           net227082, QN => n15250);
   registers_reg_58_10_inst : DFF_X1 port map( D => n8555, CK => clk, Q => 
                           net227081, QN => n14917);
   registers_reg_59_10_inst : DFF_X1 port map( D => n8554, CK => clk, Q => 
                           registers_59_10_port, QN => n15439);
   registers_reg_60_10_inst : DFF_X1 port map( D => n8553, CK => clk, Q => 
                           registers_60_10_port, QN => n14650);
   registers_reg_61_10_inst : DFF_X1 port map( D => n8552, CK => clk, Q => 
                           net227080, QN => n15641);
   registers_reg_62_10_inst : DFF_X1 port map( D => n8551, CK => clk, Q => 
                           registers_62_10_port, QN => n15130);
   registers_reg_63_10_inst : DFF_X1 port map( D => n8550, CK => clk, Q => 
                           registers_63_10_port, QN => n14513);
   to_mem_reg_10_inst : DFF_X1 port map( D => n8549, CK => clk, Q => net271357,
                           QN => n7715);
   registers_reg_64_10_inst : DFF_X1 port map( D => n8548, CK => clk, Q => 
                           net227079, QN => n16152);
   registers_reg_65_10_inst : DFF_X1 port map( D => n8547, CK => clk, Q => 
                           net227078, QN => n16101);
   registers_reg_66_10_inst : DFF_X1 port map( D => n8546, CK => clk, Q => 
                           net227077, QN => n16065);
   registers_reg_67_10_inst : DFF_X1 port map( D => n8545, CK => clk, Q => 
                           net271356, QN => n14227);
   registers_reg_68_10_inst : DFF_X1 port map( D => n8544, CK => clk, Q => 
                           registers_68_10_port, QN => n16189);
   registers_reg_69_10_inst : DFF_X1 port map( D => n8543, CK => clk, Q => 
                           net227076, QN => n16163);
   registers_reg_70_10_inst : DFF_X1 port map( D => n8542, CK => clk, Q => 
                           net227075, QN => n16064);
   registers_reg_0_9_inst : DFF_X1 port map( D => n8541, CK => clk, Q => 
                           registers_0_9_port, QN => n15860);
   registers_reg_1_9_inst : DFF_X1 port map( D => n8540, CK => clk, Q => 
                           registers_1_9_port, QN => n15596);
   registers_reg_2_9_inst : DFF_X1 port map( D => n8539, CK => clk, Q => 
                           registers_2_9_port, QN => n14787);
   registers_reg_3_9_inst : DFF_X1 port map( D => n8538, CK => clk, Q => 
                           net227074, QN => n15767);
   registers_reg_4_9_inst : DFF_X1 port map( D => n8537, CK => clk, Q => 
                           registers_4_9_port, QN => n15530);
   registers_reg_5_9_inst : DFF_X1 port map( D => n8536, CK => clk, Q => 
                           registers_5_9_port, QN => n14728);
   registers_reg_6_9_inst : DFF_X1 port map( D => n8535, CK => clk, Q => 
                           net271355, QN => n12410);
   registers_reg_7_9_inst : DFF_X1 port map( D => n8534, CK => clk, Q => 
                           registers_7_9_port, QN => n15335);
   registers_reg_8_9_inst : DFF_X1 port map( D => n8533, CK => clk, Q => 
                           net227073, QN => n15218);
   registers_reg_9_9_inst : DFF_X1 port map( D => n8532, CK => clk, Q => 
                           registers_9_9_port, QN => n14337);
   registers_reg_10_9_inst : DFF_X1 port map( D => n8531, CK => clk, Q => 
                           registers_10_9_port, QN => n14729);
   registers_reg_11_9_inst : DFF_X1 port map( D => n8530, CK => clk, Q => 
                           registers_11_9_port, QN => n14441);
   registers_reg_12_9_inst : DFF_X1 port map( D => n8529, CK => clk, Q => 
                           registers_12_9_port, QN => n15677);
   registers_reg_13_9_inst : DFF_X1 port map( D => n8528, CK => clk, Q => 
                           net227072, QN => n15087);
   registers_reg_14_9_inst : DFF_X1 port map( D => n8527, CK => clk, Q => 
                           net271354, QN => n11889);
   registers_reg_15_9_inst : DFF_X1 port map( D => n8526, CK => clk, Q => 
                           registers_15_9_port, QN => n15300);
   registers_reg_16_9_inst : DFF_X1 port map( D => n8525, CK => clk, Q => 
                           registers_16_9_port, QN => n15707);
   registers_reg_17_9_inst : DFF_X1 port map( D => n8524, CK => clk, Q => 
                           registers_17_9_port, QN => n14613);
   registers_reg_18_9_inst : DFF_X1 port map( D => n8523, CK => clk, Q => 
                           registers_18_9_port, QN => n14378);
   registers_reg_19_9_inst : DFF_X1 port map( D => n8522, CK => clk, Q => 
                           registers_19_9_port, QN => n15817);
   registers_reg_20_9_inst : DFF_X1 port map( D => n8521, CK => clk, Q => 
                           net271353, QN => n14839);
   registers_reg_21_9_inst : DFF_X1 port map( D => n8520, CK => clk, Q => 
                           net271352, QN => n12213);
   registers_reg_22_9_inst : DFF_X1 port map( D => n8519, CK => clk, Q => 
                           registers_22_9_port, QN => n15380);
   registers_reg_23_9_inst : DFF_X1 port map( D => n8518, CK => clk, Q => 
                           registers_23_9_port, QN => n15890);
   registers_reg_24_9_inst : DFF_X1 port map( D => n8517, CK => clk, Q => 
                           net227071, QN => n15188);
   registers_reg_25_9_inst : DFF_X1 port map( D => n8516, CK => clk, Q => 
                           registers_25_9_port, QN => n14307);
   registers_reg_26_9_inst : DFF_X1 port map( D => n8515, CK => clk, Q => 
                           net271351, QN => n12409);
   registers_reg_27_9_inst : DFF_X1 port map( D => n8514, CK => clk, Q => 
                           net271350, QN => n12025);
   registers_reg_28_9_inst : DFF_X1 port map( D => n8513, CK => clk, Q => 
                           net227070, QN => n15011);
   registers_reg_29_9_inst : DFF_X1 port map( D => n8512, CK => clk, Q => 
                           registers_29_9_port, QN => n15816);
   registers_reg_30_9_inst : DFF_X1 port map( D => n8511, CK => clk, Q => 
                           registers_30_9_port, QN => n14685);
   registers_reg_31_9_inst : DFF_X1 port map( D => n8510, CK => clk, Q => 
                           net227069, QN => n15743);
   registers_reg_32_9_inst : DFF_X1 port map( D => n8509, CK => clk, Q => 
                           net271349, QN => n12318);
   registers_reg_33_9_inst : DFF_X1 port map( D => n8508, CK => clk, Q => 
                           net271348, QN => n11850);
   registers_reg_34_9_inst : DFF_X1 port map( D => n8507, CK => clk, Q => 
                           registers_34_9_port, QN => n15503);
   registers_reg_35_9_inst : DFF_X1 port map( D => n8506, CK => clk, Q => 
                           net227068, QN => n15595);
   registers_reg_36_9_inst : DFF_X1 port map( D => n8505, CK => clk, Q => 
                           registers_36_9_port, QN => n15160);
   registers_reg_37_9_inst : DFF_X1 port map( D => n8504, CK => clk, Q => 
                           registers_37_9_port, QN => n14377);
   registers_reg_38_9_inst : DFF_X1 port map( D => n8503, CK => clk, Q => 
                           registers_38_9_port, QN => n15044);
   registers_reg_39_9_inst : DFF_X1 port map( D => n8502, CK => clk, Q => 
                           net271347, QN => n12179);
   registers_reg_40_9_inst : DFF_X1 port map( D => n8501, CK => clk, Q => 
                           registers_40_9_port, QN => n15088);
   registers_reg_41_9_inst : DFF_X1 port map( D => n8500, CK => clk, Q => 
                           registers_41_9_port, QN => n14442);
   registers_reg_42_9_inst : DFF_X1 port map( D => n8499, CK => clk, Q => 
                           registers_42_9_port, QN => n15928);
   registers_reg_43_9_inst : DFF_X1 port map( D => n8498, CK => clk, Q => 
                           registers_43_9_port, QN => n14895);
   registers_reg_44_9_inst : DFF_X1 port map( D => n8497, CK => clk, Q => 
                           registers_44_9_port, QN => n15473);
   registers_reg_45_9_inst : DFF_X1 port map( D => n8496, CK => clk, Q => 
                           registers_45_9_port, QN => n14788);
   registers_reg_46_9_inst : DFF_X1 port map( D => n8495, CK => clk, Q => 
                           net227067, QN => n12001);
   registers_reg_47_9_inst : DFF_X1 port map( D => n8494, CK => clk, Q => 
                           registers_47_9_port, QN => n14554);
   registers_reg_48_9_inst : DFF_X1 port map( D => n8493, CK => clk, Q => 
                           registers_48_9_port, QN => n15559);
   registers_reg_49_9_inst : DFF_X1 port map( D => n8492, CK => clk, Q => 
                           registers_49_9_port, QN => n14491);
   registers_reg_50_9_inst : DFF_X1 port map( D => n8491, CK => clk, Q => 
                           registers_50_9_port, QN => n15977);
   registers_reg_51_9_inst : DFF_X1 port map( D => n8490, CK => clk, Q => 
                           registers_51_9_port, QN => n15406);
   registers_reg_52_9_inst : DFF_X1 port map( D => n8489, CK => clk, Q => 
                           net227066, QN => n14945);
   registers_reg_53_9_inst : DFF_X1 port map( D => n8488, CK => clk, Q => 
                           net227065, QN => n15919);
   registers_reg_54_9_inst : DFF_X1 port map( D => n8487, CK => clk, Q => 
                           registers_54_9_port, QN => n14577);
   registers_reg_55_9_inst : DFF_X1 port map( D => n8486, CK => clk, Q => 
                           registers_55_9_port, QN => n12059);
   registers_reg_56_9_inst : DFF_X1 port map( D => n8485, CK => clk, Q => 
                           registers_56_9_port, QN => n16003);
   registers_reg_57_9_inst : DFF_X1 port map( D => n8484, CK => clk, Q => 
                           net227064, QN => n15249);
   registers_reg_58_9_inst : DFF_X1 port map( D => n8483, CK => clk, Q => 
                           net227063, QN => n14916);
   registers_reg_59_9_inst : DFF_X1 port map( D => n8482, CK => clk, Q => 
                           registers_59_9_port, QN => n15438);
   registers_reg_60_9_inst : DFF_X1 port map( D => n8481, CK => clk, Q => 
                           registers_60_9_port, QN => n14649);
   registers_reg_61_9_inst : DFF_X1 port map( D => n8480, CK => clk, Q => 
                           net227062, QN => n15640);
   registers_reg_62_9_inst : DFF_X1 port map( D => n8479, CK => clk, Q => 
                           registers_62_9_port, QN => n15129);
   registers_reg_63_9_inst : DFF_X1 port map( D => n8478, CK => clk, Q => 
                           registers_63_9_port, QN => n14512);
   to_mem_reg_9_inst : DFF_X1 port map( D => n8477, CK => clk, Q => net271346, 
                           QN => n7716);
   registers_reg_64_9_inst : DFF_X1 port map( D => n8476, CK => clk, Q => 
                           net227061, QN => n16151);
   registers_reg_65_9_inst : DFF_X1 port map( D => n8475, CK => clk, Q => 
                           net227060, QN => n16100);
   registers_reg_66_9_inst : DFF_X1 port map( D => n8474, CK => clk, Q => 
                           net227059, QN => n16063);
   registers_reg_67_9_inst : DFF_X1 port map( D => n8473, CK => clk, Q => 
                           net271345, QN => n14225);
   registers_reg_68_9_inst : DFF_X1 port map( D => n8472, CK => clk, Q => 
                           registers_68_9_port, QN => n16188);
   registers_reg_69_9_inst : DFF_X1 port map( D => n8471, CK => clk, Q => 
                           net227058, QN => n16162);
   registers_reg_70_9_inst : DFF_X1 port map( D => n8470, CK => clk, Q => 
                           net227057, QN => n16062);
   registers_reg_0_8_inst : DFF_X1 port map( D => n8469, CK => clk, Q => 
                           registers_0_8_port, QN => n15859);
   registers_reg_1_8_inst : DFF_X1 port map( D => n8468, CK => clk, Q => 
                           registers_1_8_port, QN => n15594);
   registers_reg_2_8_inst : DFF_X1 port map( D => n8467, CK => clk, Q => 
                           registers_2_8_port, QN => n14785);
   registers_reg_3_8_inst : DFF_X1 port map( D => n8466, CK => clk, Q => 
                           net227056, QN => n15766);
   registers_reg_4_8_inst : DFF_X1 port map( D => n8465, CK => clk, Q => 
                           registers_4_8_port, QN => n15529);
   registers_reg_5_8_inst : DFF_X1 port map( D => n8464, CK => clk, Q => 
                           registers_5_8_port, QN => n14726);
   registers_reg_6_8_inst : DFF_X1 port map( D => n8463, CK => clk, Q => 
                           net271344, QN => n12408);
   registers_reg_7_8_inst : DFF_X1 port map( D => n8462, CK => clk, Q => 
                           registers_7_8_port, QN => n15334);
   registers_reg_8_8_inst : DFF_X1 port map( D => n8461, CK => clk, Q => 
                           net227055, QN => n15217);
   registers_reg_9_8_inst : DFF_X1 port map( D => n8460, CK => clk, Q => 
                           registers_9_8_port, QN => n14336);
   registers_reg_10_8_inst : DFF_X1 port map( D => n8459, CK => clk, Q => 
                           registers_10_8_port, QN => n14727);
   registers_reg_11_8_inst : DFF_X1 port map( D => n8458, CK => clk, Q => 
                           registers_11_8_port, QN => n14439);
   registers_reg_12_8_inst : DFF_X1 port map( D => n8457, CK => clk, Q => 
                           registers_12_8_port, QN => n15676);
   registers_reg_13_8_inst : DFF_X1 port map( D => n8456, CK => clk, Q => 
                           net227054, QN => n15085);
   registers_reg_14_8_inst : DFF_X1 port map( D => n8455, CK => clk, Q => 
                           net271343, QN => n11888);
   registers_reg_15_8_inst : DFF_X1 port map( D => n8454, CK => clk, Q => 
                           registers_15_8_port, QN => n15299);
   registers_reg_16_8_inst : DFF_X1 port map( D => n8453, CK => clk, Q => 
                           registers_16_8_port, QN => n15706);
   registers_reg_17_8_inst : DFF_X1 port map( D => n8452, CK => clk, Q => 
                           registers_17_8_port, QN => n14612);
   registers_reg_18_8_inst : DFF_X1 port map( D => n8451, CK => clk, Q => 
                           registers_18_8_port, QN => n14376);
   registers_reg_19_8_inst : DFF_X1 port map( D => n8450, CK => clk, Q => 
                           registers_19_8_port, QN => n15815);
   registers_reg_20_8_inst : DFF_X1 port map( D => n8449, CK => clk, Q => 
                           net271342, QN => n14838);
   registers_reg_21_8_inst : DFF_X1 port map( D => n8448, CK => clk, Q => 
                           net271341, QN => n12212);
   registers_reg_22_8_inst : DFF_X1 port map( D => n8447, CK => clk, Q => 
                           registers_22_8_port, QN => n15379);
   registers_reg_23_8_inst : DFF_X1 port map( D => n8446, CK => clk, Q => 
                           registers_23_8_port, QN => n15888);
   registers_reg_24_8_inst : DFF_X1 port map( D => n8445, CK => clk, Q => 
                           net227053, QN => n15187);
   registers_reg_25_8_inst : DFF_X1 port map( D => n8444, CK => clk, Q => 
                           registers_25_8_port, QN => n14306);
   registers_reg_26_8_inst : DFF_X1 port map( D => n8443, CK => clk, Q => 
                           net271340, QN => n12407);
   registers_reg_27_8_inst : DFF_X1 port map( D => n8442, CK => clk, Q => 
                           net271339, QN => n12024);
   registers_reg_28_8_inst : DFF_X1 port map( D => n8441, CK => clk, Q => 
                           net227052, QN => n15010);
   registers_reg_29_8_inst : DFF_X1 port map( D => n8440, CK => clk, Q => 
                           registers_29_8_port, QN => n15812);
   registers_reg_30_8_inst : DFF_X1 port map( D => n8439, CK => clk, Q => 
                           registers_30_8_port, QN => n14684);
   registers_reg_31_8_inst : DFF_X1 port map( D => n8438, CK => clk, Q => 
                           net227051, QN => n15742);
   registers_reg_32_8_inst : DFF_X1 port map( D => n8437, CK => clk, Q => 
                           net271338, QN => n12317);
   registers_reg_33_8_inst : DFF_X1 port map( D => n8436, CK => clk, Q => 
                           net271337, QN => n11849);
   registers_reg_34_8_inst : DFF_X1 port map( D => n8435, CK => clk, Q => 
                           registers_34_8_port, QN => n15502);
   registers_reg_35_8_inst : DFF_X1 port map( D => n8434, CK => clk, Q => 
                           net227050, QN => n15593);
   registers_reg_36_8_inst : DFF_X1 port map( D => n8433, CK => clk, Q => 
                           registers_36_8_port, QN => n15159);
   registers_reg_37_8_inst : DFF_X1 port map( D => n8432, CK => clk, Q => 
                           registers_37_8_port, QN => n14375);
   registers_reg_38_8_inst : DFF_X1 port map( D => n8431, CK => clk, Q => 
                           registers_38_8_port, QN => n15043);
   registers_reg_39_8_inst : DFF_X1 port map( D => n8430, CK => clk, Q => 
                           net271336, QN => n12178);
   registers_reg_40_8_inst : DFF_X1 port map( D => n8429, CK => clk, Q => 
                           registers_40_8_port, QN => n15086);
   registers_reg_41_8_inst : DFF_X1 port map( D => n8428, CK => clk, Q => 
                           registers_41_8_port, QN => n14440);
   registers_reg_42_8_inst : DFF_X1 port map( D => n8427, CK => clk, Q => 
                           registers_42_8_port, QN => n15927);
   registers_reg_43_8_inst : DFF_X1 port map( D => n8426, CK => clk, Q => 
                           registers_43_8_port, QN => n14894);
   registers_reg_44_8_inst : DFF_X1 port map( D => n8425, CK => clk, Q => 
                           registers_44_8_port, QN => n15472);
   registers_reg_45_8_inst : DFF_X1 port map( D => n8424, CK => clk, Q => 
                           registers_45_8_port, QN => n14786);
   registers_reg_46_8_inst : DFF_X1 port map( D => n8423, CK => clk, Q => 
                           net227049, QN => n12000);
   registers_reg_47_8_inst : DFF_X1 port map( D => n8422, CK => clk, Q => 
                           registers_47_8_port, QN => n14553);
   registers_reg_48_8_inst : DFF_X1 port map( D => n8421, CK => clk, Q => 
                           registers_48_8_port, QN => n15558);
   registers_reg_49_8_inst : DFF_X1 port map( D => n8420, CK => clk, Q => 
                           registers_49_8_port, QN => n14490);
   registers_reg_50_8_inst : DFF_X1 port map( D => n8419, CK => clk, Q => 
                           registers_50_8_port, QN => n15976);
   registers_reg_51_8_inst : DFF_X1 port map( D => n8418, CK => clk, Q => 
                           registers_51_8_port, QN => n15405);
   registers_reg_52_8_inst : DFF_X1 port map( D => n8417, CK => clk, Q => 
                           net227048, QN => n14944);
   registers_reg_53_8_inst : DFF_X1 port map( D => n8416, CK => clk, Q => 
                           net227047, QN => n15918);
   registers_reg_54_8_inst : DFF_X1 port map( D => n8415, CK => clk, Q => 
                           registers_54_8_port, QN => n14576);
   registers_reg_55_8_inst : DFF_X1 port map( D => n8414, CK => clk, Q => 
                           registers_55_8_port, QN => n12058);
   registers_reg_56_8_inst : DFF_X1 port map( D => n8413, CK => clk, Q => 
                           registers_56_8_port, QN => n16013);
   registers_reg_57_8_inst : DFF_X1 port map( D => n8412, CK => clk, Q => 
                           net227046, QN => n15248);
   registers_reg_58_8_inst : DFF_X1 port map( D => n8411, CK => clk, Q => 
                           net227045, QN => n14915);
   registers_reg_59_8_inst : DFF_X1 port map( D => n8410, CK => clk, Q => 
                           registers_59_8_port, QN => n15437);
   registers_reg_60_8_inst : DFF_X1 port map( D => n8409, CK => clk, Q => 
                           registers_60_8_port, QN => n14648);
   registers_reg_61_8_inst : DFF_X1 port map( D => n8408, CK => clk, Q => 
                           net227044, QN => n15639);
   registers_reg_62_8_inst : DFF_X1 port map( D => n8407, CK => clk, Q => 
                           registers_62_8_port, QN => n15128);
   registers_reg_63_8_inst : DFF_X1 port map( D => n8406, CK => clk, Q => 
                           registers_63_8_port, QN => n14511);
   to_mem_reg_8_inst : DFF_X1 port map( D => n8405, CK => clk, Q => net271335, 
                           QN => n7717);
   registers_reg_64_8_inst : DFF_X1 port map( D => n8404, CK => clk, Q => 
                           net227043, QN => n16150);
   registers_reg_65_8_inst : DFF_X1 port map( D => n8403, CK => clk, Q => 
                           net227042, QN => n16099);
   registers_reg_66_8_inst : DFF_X1 port map( D => n8402, CK => clk, Q => 
                           net227041, QN => n16061);
   registers_reg_67_8_inst : DFF_X1 port map( D => n8401, CK => clk, Q => 
                           net271334, QN => n14219);
   registers_reg_68_8_inst : DFF_X1 port map( D => n8400, CK => clk, Q => 
                           registers_68_8_port, QN => n16187);
   registers_reg_69_8_inst : DFF_X1 port map( D => n8399, CK => clk, Q => 
                           net227040, QN => n16161);
   registers_reg_70_8_inst : DFF_X1 port map( D => n8398, CK => clk, Q => 
                           net227039, QN => n16039);
   registers_reg_0_7_inst : DFF_X1 port map( D => n8397, CK => clk, Q => 
                           registers_0_7_port, QN => n15858);
   registers_reg_1_7_inst : DFF_X1 port map( D => n8396, CK => clk, Q => 
                           registers_1_7_port, QN => n15592);
   registers_reg_2_7_inst : DFF_X1 port map( D => n8395, CK => clk, Q => 
                           registers_2_7_port, QN => n14783);
   registers_reg_3_7_inst : DFF_X1 port map( D => n8394, CK => clk, Q => 
                           net227038, QN => n15765);
   registers_reg_4_7_inst : DFF_X1 port map( D => n8393, CK => clk, Q => 
                           registers_4_7_port, QN => n15528);
   registers_reg_5_7_inst : DFF_X1 port map( D => n8392, CK => clk, Q => 
                           registers_5_7_port, QN => n14724);
   registers_reg_6_7_inst : DFF_X1 port map( D => n8391, CK => clk, Q => 
                           net271333, QN => n12369);
   registers_reg_7_7_inst : DFF_X1 port map( D => n8390, CK => clk, Q => 
                           registers_7_7_port, QN => n15333);
   registers_reg_8_7_inst : DFF_X1 port map( D => n8389, CK => clk, Q => 
                           net227037, QN => n15216);
   registers_reg_9_7_inst : DFF_X1 port map( D => n8388, CK => clk, Q => 
                           registers_9_7_port, QN => n14335);
   registers_reg_10_7_inst : DFF_X1 port map( D => n8387, CK => clk, Q => 
                           registers_10_7_port, QN => n14725);
   registers_reg_11_7_inst : DFF_X1 port map( D => n8386, CK => clk, Q => 
                           registers_11_7_port, QN => n14437);
   registers_reg_12_7_inst : DFF_X1 port map( D => n8385, CK => clk, Q => 
                           registers_12_7_port, QN => n15675);
   registers_reg_13_7_inst : DFF_X1 port map( D => n8384, CK => clk, Q => 
                           net227036, QN => n15083);
   registers_reg_14_7_inst : DFF_X1 port map( D => n8383, CK => clk, Q => 
                           net271332, QN => n11887);
   registers_reg_15_7_inst : DFF_X1 port map( D => n8382, CK => clk, Q => 
                           registers_15_7_port, QN => n15298);
   registers_reg_16_7_inst : DFF_X1 port map( D => n8381, CK => clk, Q => 
                           registers_16_7_port, QN => n15705);
   registers_reg_17_7_inst : DFF_X1 port map( D => n8380, CK => clk, Q => 
                           registers_17_7_port, QN => n14611);
   registers_reg_18_7_inst : DFF_X1 port map( D => n8379, CK => clk, Q => 
                           registers_18_7_port, QN => n14374);
   registers_reg_19_7_inst : DFF_X1 port map( D => n8378, CK => clk, Q => 
                           registers_19_7_port, QN => n15811);
   registers_reg_20_7_inst : DFF_X1 port map( D => n8377, CK => clk, Q => 
                           net271331, QN => n14837);
   registers_reg_21_7_inst : DFF_X1 port map( D => n8376, CK => clk, Q => 
                           net271330, QN => n12211);
   registers_reg_22_7_inst : DFF_X1 port map( D => n8375, CK => clk, Q => 
                           registers_22_7_port, QN => n15378);
   registers_reg_23_7_inst : DFF_X1 port map( D => n8374, CK => clk, Q => 
                           registers_23_7_port, QN => n15887);
   registers_reg_24_7_inst : DFF_X1 port map( D => n8373, CK => clk, Q => 
                           net227035, QN => n15186);
   registers_reg_25_7_inst : DFF_X1 port map( D => n8372, CK => clk, Q => 
                           registers_25_7_port, QN => n14305);
   registers_reg_26_7_inst : DFF_X1 port map( D => n8371, CK => clk, Q => 
                           net271329, QN => n12368);
   registers_reg_27_7_inst : DFF_X1 port map( D => n8370, CK => clk, Q => 
                           net271328, QN => n12023);
   registers_reg_28_7_inst : DFF_X1 port map( D => n8369, CK => clk, Q => 
                           net227034, QN => n15009);
   registers_reg_29_7_inst : DFF_X1 port map( D => n8368, CK => clk, Q => 
                           registers_29_7_port, QN => n15810);
   registers_reg_30_7_inst : DFF_X1 port map( D => n8367, CK => clk, Q => 
                           registers_30_7_port, QN => n14683);
   registers_reg_31_7_inst : DFF_X1 port map( D => n8366, CK => clk, Q => 
                           net227033, QN => n15741);
   registers_reg_32_7_inst : DFF_X1 port map( D => n8365, CK => clk, Q => 
                           net271327, QN => n12316);
   registers_reg_33_7_inst : DFF_X1 port map( D => n8364, CK => clk, Q => 
                           net271326, QN => n11847);
   registers_reg_34_7_inst : DFF_X1 port map( D => n8363, CK => clk, Q => 
                           registers_34_7_port, QN => n15501);
   registers_reg_35_7_inst : DFF_X1 port map( D => n8362, CK => clk, Q => 
                           net227032, QN => n15591);
   registers_reg_36_7_inst : DFF_X1 port map( D => n8361, CK => clk, Q => 
                           registers_36_7_port, QN => n15158);
   registers_reg_37_7_inst : DFF_X1 port map( D => n8360, CK => clk, Q => 
                           registers_37_7_port, QN => n14373);
   registers_reg_38_7_inst : DFF_X1 port map( D => n8359, CK => clk, Q => 
                           registers_38_7_port, QN => n15042);
   registers_reg_39_7_inst : DFF_X1 port map( D => n8358, CK => clk, Q => 
                           net271325, QN => n12177);
   registers_reg_40_7_inst : DFF_X1 port map( D => n8357, CK => clk, Q => 
                           registers_40_7_port, QN => n15084);
   registers_reg_41_7_inst : DFF_X1 port map( D => n8356, CK => clk, Q => 
                           registers_41_7_port, QN => n14438);
   registers_reg_42_7_inst : DFF_X1 port map( D => n8355, CK => clk, Q => 
                           registers_42_7_port, QN => n15925);
   registers_reg_43_7_inst : DFF_X1 port map( D => n8354, CK => clk, Q => 
                           registers_43_7_port, QN => n14893);
   registers_reg_44_7_inst : DFF_X1 port map( D => n8353, CK => clk, Q => 
                           registers_44_7_port, QN => n15471);
   registers_reg_45_7_inst : DFF_X1 port map( D => n8352, CK => clk, Q => 
                           registers_45_7_port, QN => n14784);
   registers_reg_46_7_inst : DFF_X1 port map( D => n8351, CK => clk, Q => 
                           net227031, QN => n11999);
   registers_reg_47_7_inst : DFF_X1 port map( D => n8350, CK => clk, Q => 
                           registers_47_7_port, QN => n14552);
   registers_reg_48_7_inst : DFF_X1 port map( D => n8349, CK => clk, Q => 
                           registers_48_7_port, QN => n15557);
   registers_reg_49_7_inst : DFF_X1 port map( D => n8348, CK => clk, Q => 
                           registers_49_7_port, QN => n14489);
   registers_reg_50_7_inst : DFF_X1 port map( D => n8347, CK => clk, Q => 
                           registers_50_7_port, QN => n15974);
   registers_reg_51_7_inst : DFF_X1 port map( D => n8346, CK => clk, Q => 
                           registers_51_7_port, QN => n15404);
   registers_reg_52_7_inst : DFF_X1 port map( D => n8345, CK => clk, Q => 
                           net227030, QN => n14943);
   registers_reg_53_7_inst : DFF_X1 port map( D => n8344, CK => clk, Q => 
                           net227029, QN => n15917);
   registers_reg_54_7_inst : DFF_X1 port map( D => n8343, CK => clk, Q => 
                           registers_54_7_port, QN => n14575);
   registers_reg_55_7_inst : DFF_X1 port map( D => n8342, CK => clk, Q => 
                           registers_55_7_port, QN => n12057);
   registers_reg_56_7_inst : DFF_X1 port map( D => n8341, CK => clk, Q => 
                           registers_56_7_port, QN => n16002);
   registers_reg_57_7_inst : DFF_X1 port map( D => n8340, CK => clk, Q => 
                           net227028, QN => n15247);
   registers_reg_58_7_inst : DFF_X1 port map( D => n8339, CK => clk, Q => 
                           net227027, QN => n14914);
   registers_reg_59_7_inst : DFF_X1 port map( D => n8338, CK => clk, Q => 
                           registers_59_7_port, QN => n15436);
   registers_reg_60_7_inst : DFF_X1 port map( D => n8337, CK => clk, Q => 
                           registers_60_7_port, QN => n14647);
   registers_reg_61_7_inst : DFF_X1 port map( D => n8336, CK => clk, Q => 
                           net227026, QN => n15638);
   registers_reg_62_7_inst : DFF_X1 port map( D => n8335, CK => clk, Q => 
                           registers_62_7_port, QN => n15127);
   registers_reg_63_7_inst : DFF_X1 port map( D => n8334, CK => clk, Q => 
                           registers_63_7_port, QN => n14510);
   to_mem_reg_7_inst : DFF_X1 port map( D => n8333, CK => clk, Q => net271324, 
                           QN => n7718);
   registers_reg_64_7_inst : DFF_X1 port map( D => n8332, CK => clk, Q => 
                           net227025, QN => n16149);
   registers_reg_65_7_inst : DFF_X1 port map( D => n8331, CK => clk, Q => 
                           net227024, QN => n16098);
   registers_reg_66_7_inst : DFF_X1 port map( D => n8330, CK => clk, Q => 
                           net227023, QN => n16060);
   registers_reg_67_7_inst : DFF_X1 port map( D => n8329, CK => clk, Q => 
                           net271323, QN => n14216);
   registers_reg_68_7_inst : DFF_X1 port map( D => n8328, CK => clk, Q => 
                           registers_68_7_port, QN => n16186);
   registers_reg_69_7_inst : DFF_X1 port map( D => n8327, CK => clk, Q => 
                           net227022, QN => n16128);
   registers_reg_70_7_inst : DFF_X1 port map( D => n8326, CK => clk, Q => 
                           net227021, QN => n16038);
   registers_reg_0_6_inst : DFF_X1 port map( D => n8325, CK => clk, Q => 
                           registers_0_6_port, QN => n15802);
   registers_reg_1_6_inst : DFF_X1 port map( D => n8324, CK => clk, Q => 
                           registers_1_6_port, QN => n15579);
   registers_reg_2_6_inst : DFF_X1 port map( D => n8323, CK => clk, Q => 
                           registers_2_6_port, QN => n14781);
   registers_reg_3_6_inst : DFF_X1 port map( D => n8322, CK => clk, Q => 
                           net227020, QN => n15764);
   registers_reg_4_6_inst : DFF_X1 port map( D => n8321, CK => clk, Q => 
                           registers_4_6_port, QN => n15527);
   registers_reg_5_6_inst : DFF_X1 port map( D => n8320, CK => clk, Q => 
                           registers_5_6_port, QN => n14722);
   registers_reg_6_6_inst : DFF_X1 port map( D => n8319, CK => clk, Q => 
                           net271322, QN => n12367);
   registers_reg_7_6_inst : DFF_X1 port map( D => n8318, CK => clk, Q => 
                           registers_7_6_port, QN => n15332);
   registers_reg_8_6_inst : DFF_X1 port map( D => n8317, CK => clk, Q => 
                           net227019, QN => n15215);
   registers_reg_9_6_inst : DFF_X1 port map( D => n8316, CK => clk, Q => 
                           registers_9_6_port, QN => n14334);
   registers_reg_10_6_inst : DFF_X1 port map( D => n8315, CK => clk, Q => 
                           registers_10_6_port, QN => n14723);
   registers_reg_11_6_inst : DFF_X1 port map( D => n8314, CK => clk, Q => 
                           registers_11_6_port, QN => n14435);
   registers_reg_12_6_inst : DFF_X1 port map( D => n8313, CK => clk, Q => 
                           registers_12_6_port, QN => n15674);
   registers_reg_13_6_inst : DFF_X1 port map( D => n8312, CK => clk, Q => 
                           net227018, QN => n15081);
   registers_reg_14_6_inst : DFF_X1 port map( D => n8311, CK => clk, Q => 
                           net271321, QN => n11886);
   registers_reg_15_6_inst : DFF_X1 port map( D => n8310, CK => clk, Q => 
                           registers_15_6_port, QN => n15297);
   registers_reg_16_6_inst : DFF_X1 port map( D => n8309, CK => clk, Q => 
                           registers_16_6_port, QN => n15704);
   registers_reg_17_6_inst : DFF_X1 port map( D => n8308, CK => clk, Q => 
                           registers_17_6_port, QN => n14610);
   registers_reg_18_6_inst : DFF_X1 port map( D => n8307, CK => clk, Q => 
                           registers_18_6_port, QN => n14372);
   registers_reg_19_6_inst : DFF_X1 port map( D => n8306, CK => clk, Q => 
                           registers_19_6_port, QN => n15809);
   registers_reg_20_6_inst : DFF_X1 port map( D => n8305, CK => clk, Q => 
                           net271320, QN => n14836);
   registers_reg_21_6_inst : DFF_X1 port map( D => n8304, CK => clk, Q => 
                           net271319, QN => n12210);
   registers_reg_22_6_inst : DFF_X1 port map( D => n8303, CK => clk, Q => 
                           registers_22_6_port, QN => n15376);
   registers_reg_23_6_inst : DFF_X1 port map( D => n8302, CK => clk, Q => 
                           registers_23_6_port, QN => n15886);
   registers_reg_24_6_inst : DFF_X1 port map( D => n8301, CK => clk, Q => 
                           net227017, QN => n15185);
   registers_reg_25_6_inst : DFF_X1 port map( D => n8300, CK => clk, Q => 
                           registers_25_6_port, QN => n14304);
   registers_reg_26_6_inst : DFF_X1 port map( D => n8299, CK => clk, Q => 
                           net271318, QN => n12366);
   registers_reg_27_6_inst : DFF_X1 port map( D => n8298, CK => clk, Q => 
                           net271317, QN => n12022);
   registers_reg_28_6_inst : DFF_X1 port map( D => n8297, CK => clk, Q => 
                           net227016, QN => n15008);
   registers_reg_29_6_inst : DFF_X1 port map( D => n8296, CK => clk, Q => 
                           registers_29_6_port, QN => n15808);
   registers_reg_30_6_inst : DFF_X1 port map( D => n8295, CK => clk, Q => 
                           registers_30_6_port, QN => n14682);
   registers_reg_31_6_inst : DFF_X1 port map( D => n8294, CK => clk, Q => 
                           net227015, QN => n15740);
   registers_reg_32_6_inst : DFF_X1 port map( D => n8293, CK => clk, Q => 
                           net271316, QN => n12315);
   registers_reg_33_6_inst : DFF_X1 port map( D => n8292, CK => clk, Q => 
                           net271315, QN => n11846);
   registers_reg_34_6_inst : DFF_X1 port map( D => n8291, CK => clk, Q => 
                           registers_34_6_port, QN => n15500);
   registers_reg_35_6_inst : DFF_X1 port map( D => n8290, CK => clk, Q => 
                           net227014, QN => n15589);
   registers_reg_36_6_inst : DFF_X1 port map( D => n8289, CK => clk, Q => 
                           registers_36_6_port, QN => n15157);
   registers_reg_37_6_inst : DFF_X1 port map( D => n8288, CK => clk, Q => 
                           registers_37_6_port, QN => n14369);
   registers_reg_38_6_inst : DFF_X1 port map( D => n8287, CK => clk, Q => 
                           registers_38_6_port, QN => n15040);
   registers_reg_39_6_inst : DFF_X1 port map( D => n8286, CK => clk, Q => 
                           net271314, QN => n12176);
   registers_reg_40_6_inst : DFF_X1 port map( D => n8285, CK => clk, Q => 
                           registers_40_6_port, QN => n15082);
   registers_reg_41_6_inst : DFF_X1 port map( D => n8284, CK => clk, Q => 
                           registers_41_6_port, QN => n14436);
   registers_reg_42_6_inst : DFF_X1 port map( D => n8283, CK => clk, Q => 
                           registers_42_6_port, QN => n15924);
   registers_reg_43_6_inst : DFF_X1 port map( D => n8282, CK => clk, Q => 
                           registers_43_6_port, QN => n14892);
   registers_reg_44_6_inst : DFF_X1 port map( D => n8281, CK => clk, Q => 
                           registers_44_6_port, QN => n15470);
   registers_reg_45_6_inst : DFF_X1 port map( D => n8280, CK => clk, Q => 
                           registers_45_6_port, QN => n14782);
   registers_reg_46_6_inst : DFF_X1 port map( D => n8279, CK => clk, Q => 
                           net227013, QN => n11998);
   registers_reg_47_6_inst : DFF_X1 port map( D => n8278, CK => clk, Q => 
                           registers_47_6_port, QN => n14551);
   registers_reg_48_6_inst : DFF_X1 port map( D => n8277, CK => clk, Q => 
                           registers_48_6_port, QN => n15556);
   registers_reg_49_6_inst : DFF_X1 port map( D => n8276, CK => clk, Q => 
                           registers_49_6_port, QN => n14488);
   registers_reg_50_6_inst : DFF_X1 port map( D => n8275, CK => clk, Q => 
                           registers_50_6_port, QN => n15973);
   registers_reg_51_6_inst : DFF_X1 port map( D => n8274, CK => clk, Q => 
                           registers_51_6_port, QN => n15403);
   registers_reg_52_6_inst : DFF_X1 port map( D => n8273, CK => clk, Q => 
                           net227012, QN => n14942);
   registers_reg_53_6_inst : DFF_X1 port map( D => n8272, CK => clk, Q => 
                           net227011, QN => n15916);
   registers_reg_54_6_inst : DFF_X1 port map( D => n8271, CK => clk, Q => 
                           registers_54_6_port, QN => n14574);
   registers_reg_55_6_inst : DFF_X1 port map( D => n8270, CK => clk, Q => 
                           registers_55_6_port, QN => n12056);
   registers_reg_56_6_inst : DFF_X1 port map( D => n8269, CK => clk, Q => 
                           registers_56_6_port, QN => n16001);
   registers_reg_57_6_inst : DFF_X1 port map( D => n8268, CK => clk, Q => 
                           net227010, QN => n15246);
   registers_reg_58_6_inst : DFF_X1 port map( D => n8267, CK => clk, Q => 
                           net227009, QN => n14913);
   registers_reg_59_6_inst : DFF_X1 port map( D => n8266, CK => clk, Q => 
                           registers_59_6_port, QN => n15435);
   registers_reg_60_6_inst : DFF_X1 port map( D => n8265, CK => clk, Q => 
                           registers_60_6_port, QN => n14646);
   registers_reg_61_6_inst : DFF_X1 port map( D => n8264, CK => clk, Q => 
                           net227008, QN => n15637);
   registers_reg_62_6_inst : DFF_X1 port map( D => n8263, CK => clk, Q => 
                           registers_62_6_port, QN => n15126);
   registers_reg_63_6_inst : DFF_X1 port map( D => n8262, CK => clk, Q => 
                           registers_63_6_port, QN => n14509);
   to_mem_reg_6_inst : DFF_X1 port map( D => n8261, CK => clk, Q => net271313, 
                           QN => n7719);
   registers_reg_64_6_inst : DFF_X1 port map( D => n8260, CK => clk, Q => 
                           net227007, QN => net271312);
   registers_reg_65_6_inst : DFF_X1 port map( D => n8259, CK => clk, Q => 
                           net227006, QN => net271311);
   registers_reg_66_6_inst : DFF_X1 port map( D => n8258, CK => clk, Q => 
                           net227005, QN => net271310);
   registers_reg_67_6_inst : DFF_X1 port map( D => n8257, CK => clk, Q => 
                           net271309, QN => n14053);
   registers_reg_68_6_inst : DFF_X1 port map( D => n8256, CK => clk, Q => 
                           registers_68_6_port, QN => net271308);
   registers_reg_69_6_inst : DFF_X1 port map( D => n8255, CK => clk, Q => 
                           net227004, QN => net271307);
   registers_reg_70_6_inst : DFF_X1 port map( D => n8254, CK => clk, Q => 
                           net227003, QN => net271306);
   registers_reg_40_5_inst : DFF_X1 port map( D => n8253, CK => clk, Q => 
                           registers_40_5_port, QN => n14996);
   registers_reg_41_5_inst : DFF_X1 port map( D => n8252, CK => clk, Q => 
                           registers_41_5_port, QN => n14293);
   registers_reg_42_5_inst : DFF_X1 port map( D => n8251, CK => clk, Q => 
                           registers_42_5_port, QN => net271305);
   registers_reg_43_5_inst : DFF_X1 port map( D => n8250, CK => clk, Q => 
                           registers_43_5_port, QN => n14862);
   registers_reg_44_5_inst : DFF_X1 port map( D => n8249, CK => clk, Q => 
                           registers_44_5_port, QN => n15357);
   registers_reg_45_5_inst : DFF_X1 port map( D => n8248, CK => clk, Q => 
                           registers_45_5_port, QN => n14642);
   registers_reg_46_5_inst : DFF_X1 port map( D => n8247, CK => clk, Q => 
                           net227002, QN => n11906);
   registers_reg_47_5_inst : DFF_X1 port map( D => n8246, CK => clk, Q => 
                           registers_47_5_port, QN => n14537);
   registers_reg_48_5_inst : DFF_X1 port map( D => n8245, CK => clk, Q => 
                           registers_48_5_port, QN => n15360);
   registers_reg_49_5_inst : DFF_X1 port map( D => n8244, CK => clk, Q => 
                           registers_49_5_port, QN => n14295);
   registers_reg_50_5_inst : DFF_X1 port map( D => n8243, CK => clk, Q => 
                           registers_50_5_port, QN => net271304);
   registers_reg_51_5_inst : DFF_X1 port map( D => n8242, CK => clk, Q => 
                           registers_51_5_port, QN => n15352);
   registers_reg_52_5_inst : DFF_X1 port map( D => n8241, CK => clk, Q => 
                           net227001, QN => n14867);
   registers_reg_53_5_inst : DFF_X1 port map( D => n8240, CK => clk, Q => 
                           net227000, QN => net271303);
   registers_reg_54_5_inst : DFF_X1 port map( D => n8239, CK => clk, Q => 
                           registers_54_5_port, QN => n14539);
   registers_reg_55_5_inst : DFF_X1 port map( D => n8238, CK => clk, Q => 
                           registers_55_5_port, QN => n12051);
   registers_reg_56_5_inst : DFF_X1 port map( D => n8237, CK => clk, Q => 
                           registers_56_5_port, QN => net271302);
   registers_reg_57_5_inst : DFF_X1 port map( D => n8236, CK => clk, Q => 
                           net226999, QN => n15242);
   registers_reg_58_5_inst : DFF_X1 port map( D => n8235, CK => clk, Q => 
                           net226998, QN => n14865);
   registers_reg_59_5_inst : DFF_X1 port map( D => n8234, CK => clk, Q => 
                           registers_59_5_port, QN => n15355);
   registers_reg_60_5_inst : DFF_X1 port map( D => n8233, CK => clk, Q => 
                           registers_60_5_port, QN => n14637);
   registers_reg_61_5_inst : DFF_X1 port map( D => n8232, CK => clk, Q => 
                           net226997, QN => n15364);
   registers_reg_62_5_inst : DFF_X1 port map( D => n8231, CK => clk, Q => 
                           registers_62_5_port, QN => n14999);
   registers_reg_63_5_inst : DFF_X1 port map( D => n8230, CK => clk, Q => 
                           registers_63_5_port, QN => n14298);
   registers_reg_0_5_inst : DFF_X1 port map( D => n8229, CK => clk, Q => 
                           registers_0_5_port, QN => n15800);
   registers_reg_1_5_inst : DFF_X1 port map( D => n8228, CK => clk, Q => 
                           registers_1_5_port, QN => n15584);
   registers_reg_2_5_inst : DFF_X1 port map( D => n8227, CK => clk, Q => 
                           registers_2_5_port, QN => n14780);
   registers_reg_3_5_inst : DFF_X1 port map( D => n8226, CK => clk, Q => 
                           net226996, QN => n15763);
   registers_reg_4_5_inst : DFF_X1 port map( D => n8225, CK => clk, Q => 
                           registers_4_5_port, QN => n15526);
   registers_reg_5_5_inst : DFF_X1 port map( D => n8224, CK => clk, Q => 
                           registers_5_5_port, QN => n14720);
   registers_reg_6_5_inst : DFF_X1 port map( D => n8223, CK => clk, Q => 
                           net271301, QN => n12365);
   registers_reg_7_5_inst : DFF_X1 port map( D => n8222, CK => clk, Q => 
                           registers_7_5_port, QN => n15331);
   registers_reg_8_5_inst : DFF_X1 port map( D => n8221, CK => clk, Q => 
                           net226995, QN => n15214);
   registers_reg_9_5_inst : DFF_X1 port map( D => n8220, CK => clk, Q => 
                           registers_9_5_port, QN => n14333);
   registers_reg_10_5_inst : DFF_X1 port map( D => n8219, CK => clk, Q => 
                           registers_10_5_port, QN => n14721);
   registers_reg_11_5_inst : DFF_X1 port map( D => n8218, CK => clk, Q => 
                           registers_11_5_port, QN => n14434);
   registers_reg_12_5_inst : DFF_X1 port map( D => n8217, CK => clk, Q => 
                           registers_12_5_port, QN => n15673);
   registers_reg_13_5_inst : DFF_X1 port map( D => n8216, CK => clk, Q => 
                           net226994, QN => n15080);
   registers_reg_14_5_inst : DFF_X1 port map( D => n8215, CK => clk, Q => 
                           net271300, QN => n11885);
   registers_reg_15_5_inst : DFF_X1 port map( D => n8214, CK => clk, Q => 
                           registers_15_5_port, QN => n15296);
   registers_reg_16_5_inst : DFF_X1 port map( D => n8213, CK => clk, Q => 
                           registers_16_5_port, QN => n15703);
   registers_reg_17_5_inst : DFF_X1 port map( D => n8212, CK => clk, Q => 
                           registers_17_5_port, QN => n14609);
   registers_reg_18_5_inst : DFF_X1 port map( D => n8211, CK => clk, Q => 
                           registers_18_5_port, QN => n14368);
   registers_reg_19_5_inst : DFF_X1 port map( D => n8210, CK => clk, Q => 
                           registers_19_5_port, QN => n15807);
   registers_reg_20_5_inst : DFF_X1 port map( D => n8209, CK => clk, Q => 
                           net271299, QN => n14835);
   registers_reg_21_5_inst : DFF_X1 port map( D => n8208, CK => clk, Q => 
                           net271298, QN => n12209);
   registers_reg_22_5_inst : DFF_X1 port map( D => n8207, CK => clk, Q => 
                           registers_22_5_port, QN => n15375);
   registers_reg_23_5_inst : DFF_X1 port map( D => n8206, CK => clk, Q => 
                           registers_23_5_port, QN => n15885);
   registers_reg_24_5_inst : DFF_X1 port map( D => n8205, CK => clk, Q => 
                           net226993, QN => n15184);
   registers_reg_25_5_inst : DFF_X1 port map( D => n8204, CK => clk, Q => 
                           registers_25_5_port, QN => n14303);
   registers_reg_26_5_inst : DFF_X1 port map( D => n8203, CK => clk, Q => 
                           net271297, QN => n12364);
   registers_reg_27_5_inst : DFF_X1 port map( D => n8202, CK => clk, Q => 
                           net271296, QN => n12021);
   registers_reg_28_5_inst : DFF_X1 port map( D => n8201, CK => clk, Q => 
                           net226992, QN => n15007);
   registers_reg_29_5_inst : DFF_X1 port map( D => n8200, CK => clk, Q => 
                           registers_29_5_port, QN => n15806);
   registers_reg_30_5_inst : DFF_X1 port map( D => n8199, CK => clk, Q => 
                           registers_30_5_port, QN => n14681);
   registers_reg_31_5_inst : DFF_X1 port map( D => n8198, CK => clk, Q => 
                           net226991, QN => n15739);
   registers_reg_32_5_inst : DFF_X1 port map( D => n8197, CK => clk, Q => 
                           net271295, QN => n12308);
   registers_reg_33_5_inst : DFF_X1 port map( D => n8196, CK => clk, Q => 
                           net271294, QN => n11584);
   registers_reg_34_5_inst : DFF_X1 port map( D => n8195, CK => clk, Q => 
                           registers_34_5_port, QN => n15358);
   registers_reg_35_5_inst : DFF_X1 port map( D => n8194, CK => clk, Q => 
                           net226990, QN => n15363);
   registers_reg_36_5_inst : DFF_X1 port map( D => n8193, CK => clk, Q => 
                           registers_36_5_port, QN => n15000);
   registers_reg_37_5_inst : DFF_X1 port map( D => n8192, CK => clk, Q => 
                           registers_37_5_port, QN => n14290);
   registers_reg_38_5_inst : DFF_X1 port map( D => n8191, CK => clk, Q => 
                           registers_38_5_port, QN => n14993);
   registers_reg_39_5_inst : DFF_X1 port map( D => n8190, CK => clk, Q => 
                           net271293, QN => n12162);
   to_mem_reg_5_inst : DFF_X1 port map( D => n8189, CK => clk, Q => net271292, 
                           QN => n7720);
   registers_reg_64_5_inst : DFF_X1 port map( D => n8188, CK => clk, Q => 
                           net226989, QN => n16125);
   registers_reg_65_5_inst : DFF_X1 port map( D => n8187, CK => clk, Q => 
                           net226988, QN => n16087);
   registers_reg_66_5_inst : DFF_X1 port map( D => n8186, CK => clk, Q => 
                           net226987, QN => n16041);
   registers_reg_67_5_inst : DFF_X1 port map( D => n8185, CK => clk, Q => 
                           net271291, QN => n14212);
   registers_reg_68_5_inst : DFF_X1 port map( D => n8184, CK => clk, Q => 
                           registers_68_5_port, QN => n16175);
   registers_reg_69_5_inst : DFF_X1 port map( D => n8183, CK => clk, Q => 
                           net226986, QN => n16127);
   registers_reg_70_5_inst : DFF_X1 port map( D => n8182, CK => clk, Q => 
                           net226985, QN => n16037);
   registers_reg_24_4_inst : DFF_X1 port map( D => n8181, CK => clk, Q => 
                           net226984, QN => n15002);
   registers_reg_25_4_inst : DFF_X1 port map( D => n8180, CK => clk, Q => 
                           registers_25_4_port, QN => n14283);
   registers_reg_26_4_inst : DFF_X1 port map( D => n8179, CK => clk, Q => 
                           net271290, QN => n12341);
   registers_reg_27_4_inst : DFF_X1 port map( D => n8178, CK => clk, Q => 
                           net271289, QN => n12017);
   registers_reg_28_4_inst : DFF_X1 port map( D => n8177, CK => clk, Q => 
                           net226983, QN => n14990);
   registers_reg_29_4_inst : DFF_X1 port map( D => n8176, CK => clk, Q => 
                           registers_29_4_port, QN => net271288);
   registers_reg_30_4_inst : DFF_X1 port map( D => n8175, CK => clk, Q => 
                           registers_30_4_port, QN => n14639);
   registers_reg_31_4_inst : DFF_X1 port map( D => n8174, CK => clk, Q => 
                           net226982, QN => n15368);
   registers_reg_48_4_inst : DFF_X1 port map( D => n8173, CK => clk, Q => 
                           registers_48_4_port, QN => n15359);
   registers_reg_49_4_inst : DFF_X1 port map( D => n8172, CK => clk, Q => 
                           registers_49_4_port, QN => n14294);
   registers_reg_50_4_inst : DFF_X1 port map( D => n8171, CK => clk, Q => 
                           registers_50_4_port, QN => net271287);
   registers_reg_51_4_inst : DFF_X1 port map( D => n8170, CK => clk, Q => 
                           registers_51_4_port, QN => n15351);
   registers_reg_52_4_inst : DFF_X1 port map( D => n8169, CK => clk, Q => 
                           net226981, QN => n14866);
   registers_reg_53_4_inst : DFF_X1 port map( D => n8168, CK => clk, Q => 
                           net226980, QN => net271286);
   registers_reg_54_4_inst : DFF_X1 port map( D => n8167, CK => clk, Q => 
                           registers_54_4_port, QN => n14538);
   registers_reg_55_4_inst : DFF_X1 port map( D => n8166, CK => clk, Q => 
                           registers_55_4_port, QN => n12050);
   registers_reg_56_4_inst : DFF_X1 port map( D => n8165, CK => clk, Q => 
                           registers_56_4_port, QN => net271285);
   registers_reg_57_4_inst : DFF_X1 port map( D => n8164, CK => clk, Q => 
                           net226979, QN => n15241);
   registers_reg_58_4_inst : DFF_X1 port map( D => n8163, CK => clk, Q => 
                           net226978, QN => n14864);
   registers_reg_59_4_inst : DFF_X1 port map( D => n8162, CK => clk, Q => 
                           registers_59_4_port, QN => n15354);
   registers_reg_60_4_inst : DFF_X1 port map( D => n8161, CK => clk, Q => 
                           registers_60_4_port, QN => n14636);
   registers_reg_61_4_inst : DFF_X1 port map( D => n8160, CK => clk, Q => 
                           net226977, QN => n15362);
   registers_reg_62_4_inst : DFF_X1 port map( D => n8159, CK => clk, Q => 
                           registers_62_4_port, QN => n14998);
   registers_reg_63_4_inst : DFF_X1 port map( D => n8158, CK => clk, Q => 
                           registers_63_4_port, QN => n14297);
   registers_reg_0_4_inst : DFF_X1 port map( D => n8157, CK => clk, Q => 
                           registers_0_4_port, QN => n15799);
   registers_reg_1_4_inst : DFF_X1 port map( D => n8156, CK => clk, Q => 
                           registers_1_4_port, QN => n15583);
   registers_reg_2_4_inst : DFF_X1 port map( D => n8155, CK => clk, Q => 
                           registers_2_4_port, QN => n14778);
   registers_reg_3_4_inst : DFF_X1 port map( D => n8154, CK => clk, Q => 
                           net226976, QN => n15762);
   registers_reg_4_4_inst : DFF_X1 port map( D => n8153, CK => clk, Q => 
                           registers_4_4_port, QN => n15525);
   registers_reg_5_4_inst : DFF_X1 port map( D => n8152, CK => clk, Q => 
                           registers_5_4_port, QN => n14718);
   registers_reg_6_4_inst : DFF_X1 port map( D => n8151, CK => clk, Q => 
                           net271284, QN => n12363);
   registers_reg_7_4_inst : DFF_X1 port map( D => n8150, CK => clk, Q => 
                           registers_7_4_port, QN => n15330);
   registers_reg_8_4_inst : DFF_X1 port map( D => n8149, CK => clk, Q => 
                           net226975, QN => n15213);
   registers_reg_9_4_inst : DFF_X1 port map( D => n8148, CK => clk, Q => 
                           registers_9_4_port, QN => n14332);
   registers_reg_10_4_inst : DFF_X1 port map( D => n8147, CK => clk, Q => 
                           registers_10_4_port, QN => n14719);
   registers_reg_11_4_inst : DFF_X1 port map( D => n8146, CK => clk, Q => 
                           registers_11_4_port, QN => n14432);
   registers_reg_12_4_inst : DFF_X1 port map( D => n8145, CK => clk, Q => 
                           registers_12_4_port, QN => n15672);
   registers_reg_13_4_inst : DFF_X1 port map( D => n8144, CK => clk, Q => 
                           net226974, QN => n15078);
   registers_reg_14_4_inst : DFF_X1 port map( D => n8143, CK => clk, Q => 
                           net271283, QN => n11884);
   registers_reg_15_4_inst : DFF_X1 port map( D => n8142, CK => clk, Q => 
                           registers_15_4_port, QN => n15295);
   registers_reg_16_4_inst : DFF_X1 port map( D => n8141, CK => clk, Q => 
                           registers_16_4_port, QN => n15366);
   registers_reg_17_4_inst : DFF_X1 port map( D => n8140, CK => clk, Q => 
                           registers_17_4_port, QN => n14569);
   registers_reg_18_4_inst : DFF_X1 port map( D => n8139, CK => clk, Q => 
                           registers_18_4_port, QN => n14289);
   registers_reg_19_4_inst : DFF_X1 port map( D => n8138, CK => clk, Q => 
                           registers_19_4_port, QN => net271282);
   registers_reg_20_4_inst : DFF_X1 port map( D => n8137, CK => clk, Q => 
                           net271281, QN => n14823);
   registers_reg_21_4_inst : DFF_X1 port map( D => n8136, CK => clk, Q => 
                           net271280, QN => n12195);
   registers_reg_22_4_inst : DFF_X1 port map( D => n8135, CK => clk, Q => 
                           registers_22_4_port, QN => n15350);
   registers_reg_23_4_inst : DFF_X1 port map( D => n8134, CK => clk, Q => 
                           registers_23_4_port, QN => net271279);
   registers_reg_32_4_inst : DFF_X1 port map( D => n8133, CK => clk, Q => 
                           net271278, QN => n12313);
   registers_reg_33_4_inst : DFF_X1 port map( D => n8132, CK => clk, Q => 
                           net271277, QN => n11844);
   registers_reg_34_4_inst : DFF_X1 port map( D => n8131, CK => clk, Q => 
                           registers_34_4_port, QN => n15499);
   registers_reg_35_4_inst : DFF_X1 port map( D => n8130, CK => clk, Q => 
                           net226973, QN => n15588);
   registers_reg_36_4_inst : DFF_X1 port map( D => n8129, CK => clk, Q => 
                           registers_36_4_port, QN => n15155);
   registers_reg_37_4_inst : DFF_X1 port map( D => n8128, CK => clk, Q => 
                           registers_37_4_port, QN => n14367);
   registers_reg_38_4_inst : DFF_X1 port map( D => n8127, CK => clk, Q => 
                           registers_38_4_port, QN => n15039);
   registers_reg_39_4_inst : DFF_X1 port map( D => n8126, CK => clk, Q => 
                           net271276, QN => n12175);
   registers_reg_40_4_inst : DFF_X1 port map( D => n8125, CK => clk, Q => 
                           registers_40_4_port, QN => n15079);
   registers_reg_41_4_inst : DFF_X1 port map( D => n8124, CK => clk, Q => 
                           registers_41_4_port, QN => n14433);
   registers_reg_42_4_inst : DFF_X1 port map( D => n8123, CK => clk, Q => 
                           registers_42_4_port, QN => n15923);
   registers_reg_43_4_inst : DFF_X1 port map( D => n8122, CK => clk, Q => 
                           registers_43_4_port, QN => n14891);
   registers_reg_44_4_inst : DFF_X1 port map( D => n8121, CK => clk, Q => 
                           registers_44_4_port, QN => n15469);
   registers_reg_45_4_inst : DFF_X1 port map( D => n8120, CK => clk, Q => 
                           registers_45_4_port, QN => n14779);
   registers_reg_46_4_inst : DFF_X1 port map( D => n8119, CK => clk, Q => 
                           net226972, QN => n11997);
   registers_reg_47_4_inst : DFF_X1 port map( D => n8118, CK => clk, Q => 
                           registers_47_4_port, QN => n14550);
   to_mem_reg_4_inst : DFF_X1 port map( D => n8117, CK => clk, Q => net271275, 
                           QN => n7721);
   registers_reg_64_4_inst : DFF_X1 port map( D => n8116, CK => clk, Q => 
                           net226971, QN => n16124);
   registers_reg_65_4_inst : DFF_X1 port map( D => n8115, CK => clk, Q => 
                           net226970, QN => n16086);
   registers_reg_66_4_inst : DFF_X1 port map( D => n8114, CK => clk, Q => 
                           net226969, QN => n16040);
   registers_reg_67_4_inst : DFF_X1 port map( D => n8113, CK => clk, Q => 
                           net271274, QN => n14071);
   registers_reg_68_4_inst : DFF_X1 port map( D => n8112, CK => clk, Q => 
                           registers_68_4_port, QN => n16174);
   registers_reg_69_4_inst : DFF_X1 port map( D => n8111, CK => clk, Q => 
                           net226968, QN => n16126);
   registers_reg_70_4_inst : DFF_X1 port map( D => n8110, CK => clk, Q => 
                           net226967, QN => n16036);
   registers_reg_71_31_inst : DFF_X1 port map( D => n8109, CK => clk, Q => 
                           net226966, QN => n14051);
   out1_reg_31_inst : DFF_X1 port map( D => n8108, CK => clk, Q => out1(31), QN
                           => net226965);
   registers_reg_71_30_inst : DFF_X1 port map( D => n8107, CK => clk, Q => 
                           net226964, QN => n14860);
   out1_reg_30_inst : DFF_X1 port map( D => n8106, CK => clk, Q => out1(30), QN
                           => net226963);
   registers_reg_71_29_inst : DFF_X1 port map( D => n8105, CK => clk, Q => 
                           net226962, QN => n14988);
   out1_reg_29_inst : DFF_X1 port map( D => n8104, CK => clk, Q => out1(29), QN
                           => net226961);
   registers_reg_71_28_inst : DFF_X1 port map( D => n8103, CK => clk, Q => 
                           net226960, QN => n14987);
   out1_reg_28_inst : DFF_X1 port map( D => n8102, CK => clk, Q => out1(28), QN
                           => net226959);
   registers_reg_71_27_inst : DFF_X1 port map( D => n8101, CK => clk, Q => 
                           net226958, QN => n14986);
   out1_reg_27_inst : DFF_X1 port map( D => n8100, CK => clk, Q => out1(27), QN
                           => net226957);
   registers_reg_71_26_inst : DFF_X1 port map( D => n8099, CK => clk, Q => 
                           net226956, QN => n14985);
   out1_reg_26_inst : DFF_X1 port map( D => n8098, CK => clk, Q => out1(26), QN
                           => net226955);
   registers_reg_71_25_inst : DFF_X1 port map( D => n8097, CK => clk, Q => 
                           net226954, QN => n14984);
   out1_reg_25_inst : DFF_X1 port map( D => n8096, CK => clk, Q => out1(25), QN
                           => net226953);
   registers_reg_71_24_inst : DFF_X1 port map( D => n8095, CK => clk, Q => 
                           net226952, QN => n14983);
   out1_reg_24_inst : DFF_X1 port map( D => n8094, CK => clk, Q => out1(24), QN
                           => net226951);
   registers_reg_71_23_inst : DFF_X1 port map( D => n8093, CK => clk, Q => 
                           net226950, QN => n14979);
   out1_reg_23_inst : DFF_X1 port map( D => n8092, CK => clk, Q => out1(23), QN
                           => net226949);
   registers_reg_71_22_inst : DFF_X1 port map( D => n8091, CK => clk, Q => 
                           net226948, QN => n14982);
   out1_reg_22_inst : DFF_X1 port map( D => n8090, CK => clk, Q => out1(22), QN
                           => net226947);
   registers_reg_71_21_inst : DFF_X1 port map( D => n8089, CK => clk, Q => 
                           net226946, QN => n14981);
   out1_reg_21_inst : DFF_X1 port map( D => n8088, CK => clk, Q => out1(21), QN
                           => net226945);
   registers_reg_71_20_inst : DFF_X1 port map( D => n8087, CK => clk, Q => 
                           net226944, QN => n14978);
   out1_reg_20_inst : DFF_X1 port map( D => n8086, CK => clk, Q => out1(20), QN
                           => net226943);
   registers_reg_71_19_inst : DFF_X1 port map( D => n8085, CK => clk, Q => 
                           net226942, QN => n14977);
   out1_reg_19_inst : DFF_X1 port map( D => n8084, CK => clk, Q => out1(19), QN
                           => net226941);
   registers_reg_71_18_inst : DFF_X1 port map( D => n8083, CK => clk, Q => 
                           net226940, QN => n14976);
   out1_reg_18_inst : DFF_X1 port map( D => n8082, CK => clk, Q => out1(18), QN
                           => net226939);
   registers_reg_71_17_inst : DFF_X1 port map( D => n8081, CK => clk, Q => 
                           net226938, QN => n14975);
   out1_reg_17_inst : DFF_X1 port map( D => n8080, CK => clk, Q => out1(17), QN
                           => net226937);
   registers_reg_71_16_inst : DFF_X1 port map( D => n8079, CK => clk, Q => 
                           net226936, QN => n14974);
   out1_reg_16_inst : DFF_X1 port map( D => n8078, CK => clk, Q => out1(16), QN
                           => net226935);
   registers_reg_71_15_inst : DFF_X1 port map( D => n8077, CK => clk, Q => 
                           net226934, QN => n14973);
   out1_reg_15_inst : DFF_X1 port map( D => n8076, CK => clk, Q => out1(15), QN
                           => net226933);
   registers_reg_71_14_inst : DFF_X1 port map( D => n8075, CK => clk, Q => 
                           net226932, QN => n14972);
   out1_reg_14_inst : DFF_X1 port map( D => n8074, CK => clk, Q => out1(14), QN
                           => net226931);
   registers_reg_71_13_inst : DFF_X1 port map( D => n8073, CK => clk, Q => 
                           net226930, QN => n14971);
   out1_reg_13_inst : DFF_X1 port map( D => n8072, CK => clk, Q => out1(13), QN
                           => net226929);
   registers_reg_71_12_inst : DFF_X1 port map( D => n8071, CK => clk, Q => 
                           net226928, QN => n14970);
   out1_reg_12_inst : DFF_X1 port map( D => n8070, CK => clk, Q => out1(12), QN
                           => net226927);
   registers_reg_71_11_inst : DFF_X1 port map( D => n8069, CK => clk, Q => 
                           net226926, QN => n14969);
   out1_reg_11_inst : DFF_X1 port map( D => n8068, CK => clk, Q => out1(11), QN
                           => net226925);
   registers_reg_71_10_inst : DFF_X1 port map( D => n8067, CK => clk, Q => 
                           net226924, QN => n14968);
   out1_reg_10_inst : DFF_X1 port map( D => n8066, CK => clk, Q => out1(10), QN
                           => net226923);
   registers_reg_71_9_inst : DFF_X1 port map( D => n8065, CK => clk, Q => 
                           net226922, QN => n14967);
   out1_reg_9_inst : DFF_X1 port map( D => n8064, CK => clk, Q => out1(9), QN 
                           => net226921);
   registers_reg_71_8_inst : DFF_X1 port map( D => n8063, CK => clk, Q => 
                           net226920, QN => n14966);
   out1_reg_8_inst : DFF_X1 port map( D => n8062, CK => clk, Q => out1(8), QN 
                           => net226919);
   registers_reg_71_7_inst : DFF_X1 port map( D => n8061, CK => clk, Q => 
                           net226918, QN => n14965);
   out1_reg_7_inst : DFF_X1 port map( D => n8060, CK => clk, Q => out1(7), QN 
                           => net226917);
   registers_reg_71_6_inst : DFF_X1 port map( D => n8059, CK => clk, Q => 
                           net226916, QN => n14868);
   out1_reg_6_inst : DFF_X1 port map( D => n8058, CK => clk, Q => out1(6), QN 
                           => net226915);
   registers_reg_71_5_inst : DFF_X1 port map( D => n8057, CK => clk, Q => 
                           net226914, QN => n14964);
   out1_reg_5_inst : DFF_X1 port map( D => n8056, CK => clk, Q => out1(5), QN 
                           => net226913);
   registers_reg_71_4_inst : DFF_X1 port map( D => n8055, CK => clk, Q => 
                           net226912, QN => n14963);
   out1_reg_4_inst : DFF_X1 port map( D => n8054, CK => clk, Q => out1(4), QN 
                           => net226911);
   registers_reg_24_3_inst : DFF_X1 port map( D => n8053, CK => clk, Q => 
                           net226910, QN => n15001);
   registers_reg_25_3_inst : DFF_X1 port map( D => n8052, CK => clk, Q => 
                           registers_25_3_port, QN => n14282);
   registers_reg_26_3_inst : DFF_X1 port map( D => n8051, CK => clk, Q => 
                           net271273, QN => n12340);
   registers_reg_27_3_inst : DFF_X1 port map( D => n8050, CK => clk, Q => 
                           net271272, QN => n12016);
   registers_reg_28_3_inst : DFF_X1 port map( D => n8049, CK => clk, Q => 
                           net226909, QN => n14989);
   registers_reg_29_3_inst : DFF_X1 port map( D => n8048, CK => clk, Q => 
                           registers_29_3_port, QN => net271271);
   registers_reg_30_3_inst : DFF_X1 port map( D => n8047, CK => clk, Q => 
                           registers_30_3_port, QN => n14638);
   registers_reg_31_3_inst : DFF_X1 port map( D => n8046, CK => clk, Q => 
                           net226908, QN => n15367);
   registers_reg_40_3_inst : DFF_X1 port map( D => n8045, CK => clk, Q => 
                           registers_40_3_port, QN => n14995);
   registers_reg_41_3_inst : DFF_X1 port map( D => n8044, CK => clk, Q => 
                           registers_41_3_port, QN => n14292);
   registers_reg_42_3_inst : DFF_X1 port map( D => n8043, CK => clk, Q => 
                           registers_42_3_port, QN => net271270);
   registers_reg_43_3_inst : DFF_X1 port map( D => n8042, CK => clk, Q => 
                           registers_43_3_port, QN => n14861);
   registers_reg_44_3_inst : DFF_X1 port map( D => n8041, CK => clk, Q => 
                           registers_44_3_port, QN => n15356);
   registers_reg_45_3_inst : DFF_X1 port map( D => n8040, CK => clk, Q => 
                           registers_45_3_port, QN => n14641);
   registers_reg_46_3_inst : DFF_X1 port map( D => n8039, CK => clk, Q => 
                           net226907, QN => n11905);
   registers_reg_47_3_inst : DFF_X1 port map( D => n8038, CK => clk, Q => 
                           registers_47_3_port, QN => n14536);
   registers_reg_56_3_inst : DFF_X1 port map( D => n8037, CK => clk, Q => 
                           registers_56_3_port, QN => net271269);
   registers_reg_57_3_inst : DFF_X1 port map( D => n8036, CK => clk, Q => 
                           net226906, QN => n15240);
   registers_reg_58_3_inst : DFF_X1 port map( D => n8035, CK => clk, Q => 
                           net226905, QN => n14863);
   registers_reg_59_3_inst : DFF_X1 port map( D => n8034, CK => clk, Q => 
                           registers_59_3_port, QN => n15353);
   registers_reg_60_3_inst : DFF_X1 port map( D => n8033, CK => clk, Q => 
                           registers_60_3_port, QN => n14635);
   registers_reg_61_3_inst : DFF_X1 port map( D => n8032, CK => clk, Q => 
                           net226904, QN => n15361);
   registers_reg_62_3_inst : DFF_X1 port map( D => n8031, CK => clk, Q => 
                           registers_62_3_port, QN => n14997);
   registers_reg_63_3_inst : DFF_X1 port map( D => n8030, CK => clk, Q => 
                           registers_63_3_port, QN => n14296);
   registers_reg_0_3_inst : DFF_X1 port map( D => n8029, CK => clk, Q => 
                           registers_0_3_port, QN => n15798);
   registers_reg_1_3_inst : DFF_X1 port map( D => n8028, CK => clk, Q => 
                           registers_1_3_port, QN => n15582);
   registers_reg_2_3_inst : DFF_X1 port map( D => n8027, CK => clk, Q => 
                           registers_2_3_port, QN => n14777);
   registers_reg_3_3_inst : DFF_X1 port map( D => n8026, CK => clk, Q => 
                           net226903, QN => n15761);
   registers_reg_4_3_inst : DFF_X1 port map( D => n8025, CK => clk, Q => 
                           registers_4_3_port, QN => n15524);
   registers_reg_5_3_inst : DFF_X1 port map( D => n8024, CK => clk, Q => 
                           registers_5_3_port, QN => n14717);
   registers_reg_6_3_inst : DFF_X1 port map( D => n8023, CK => clk, Q => 
                           net271268, QN => n12362);
   registers_reg_7_3_inst : DFF_X1 port map( D => n8022, CK => clk, Q => 
                           registers_7_3_port, QN => n15329);
   registers_reg_8_3_inst : DFF_X1 port map( D => n8021, CK => clk, Q => 
                           net226902, QN => n15003);
   registers_reg_9_3_inst : DFF_X1 port map( D => n8020, CK => clk, Q => 
                           registers_9_3_port, QN => n14288);
   registers_reg_10_3_inst : DFF_X1 port map( D => n8019, CK => clk, Q => 
                           registers_10_3_port, QN => n14640);
   registers_reg_11_3_inst : DFF_X1 port map( D => n8018, CK => clk, Q => 
                           registers_11_3_port, QN => n14291);
   registers_reg_12_3_inst : DFF_X1 port map( D => n8017, CK => clk, Q => 
                           registers_12_3_port, QN => n15365);
   registers_reg_13_3_inst : DFF_X1 port map( D => n8016, CK => clk, Q => 
                           net226901, QN => n14994);
   registers_reg_14_3_inst : DFF_X1 port map( D => n8015, CK => clk, Q => 
                           net271267, QN => n11627);
   registers_reg_15_3_inst : DFF_X1 port map( D => n8014, CK => clk, Q => 
                           registers_15_3_port, QN => n15284);
   registers_reg_16_3_inst : DFF_X1 port map( D => n8013, CK => clk, Q => 
                           registers_16_3_port, QN => n15702);
   registers_reg_17_3_inst : DFF_X1 port map( D => n8012, CK => clk, Q => 
                           registers_17_3_port, QN => n14608);
   registers_reg_18_3_inst : DFF_X1 port map( D => n8011, CK => clk, Q => 
                           registers_18_3_port, QN => n14366);
   registers_reg_19_3_inst : DFF_X1 port map( D => n8010, CK => clk, Q => 
                           registers_19_3_port, QN => n15805);
   registers_reg_20_3_inst : DFF_X1 port map( D => n8009, CK => clk, Q => 
                           net271266, QN => n14834);
   registers_reg_21_3_inst : DFF_X1 port map( D => n8008, CK => clk, Q => 
                           net271265, QN => n12208);
   registers_reg_22_3_inst : DFF_X1 port map( D => n8007, CK => clk, Q => 
                           registers_22_3_port, QN => n15374);
   registers_reg_23_3_inst : DFF_X1 port map( D => n8006, CK => clk, Q => 
                           registers_23_3_port, QN => n15884);
   registers_reg_32_3_inst : DFF_X1 port map( D => n8005, CK => clk, Q => 
                           net271264, QN => n12312);
   registers_reg_33_3_inst : DFF_X1 port map( D => n8004, CK => clk, Q => 
                           net271263, QN => n11842);
   registers_reg_34_3_inst : DFF_X1 port map( D => n8003, CK => clk, Q => 
                           registers_34_3_port, QN => n15498);
   registers_reg_35_3_inst : DFF_X1 port map( D => n8002, CK => clk, Q => 
                           net226900, QN => n15587);
   registers_reg_36_3_inst : DFF_X1 port map( D => n8001, CK => clk, Q => 
                           registers_36_3_port, QN => n15154);
   registers_reg_37_3_inst : DFF_X1 port map( D => n8000, CK => clk, Q => 
                           registers_37_3_port, QN => n14365);
   registers_reg_38_3_inst : DFF_X1 port map( D => n7999, CK => clk, Q => 
                           registers_38_3_port, QN => n15038);
   registers_reg_39_3_inst : DFF_X1 port map( D => n7998, CK => clk, Q => 
                           net271262, QN => n12174);
   registers_reg_48_3_inst : DFF_X1 port map( D => n7997, CK => clk, Q => 
                           registers_48_3_port, QN => n15555);
   registers_reg_49_3_inst : DFF_X1 port map( D => n7996, CK => clk, Q => 
                           registers_49_3_port, QN => n14487);
   registers_reg_50_3_inst : DFF_X1 port map( D => n7995, CK => clk, Q => 
                           registers_50_3_port, QN => n15972);
   registers_reg_51_3_inst : DFF_X1 port map( D => n7994, CK => clk, Q => 
                           registers_51_3_port, QN => n15402);
   registers_reg_52_3_inst : DFF_X1 port map( D => n7993, CK => clk, Q => 
                           net226899, QN => n14941);
   registers_reg_53_3_inst : DFF_X1 port map( D => n7992, CK => clk, Q => 
                           net226898, QN => n15915);
   registers_reg_54_3_inst : DFF_X1 port map( D => n7991, CK => clk, Q => 
                           registers_54_3_port, QN => n14572);
   registers_reg_55_3_inst : DFF_X1 port map( D => n7990, CK => clk, Q => 
                           registers_55_3_port, QN => n12054);
   to_mem_reg_3_inst : DFF_X1 port map( D => n7989, CK => clk, Q => net271261, 
                           QN => n7722);
   registers_reg_64_3_inst : DFF_X1 port map( D => n7988, CK => clk, Q => 
                           net226897, QN => n16204);
   registers_reg_65_3_inst : DFF_X1 port map( D => n7987, CK => clk, Q => 
                           net226896, QN => n16114);
   registers_reg_66_3_inst : DFF_X1 port map( D => n7986, CK => clk, Q => 
                           net226895, QN => n16122);
   registers_reg_67_3_inst : DFF_X1 port map( D => n7985, CK => clk, Q => 
                           net271260, QN => n14287);
   registers_reg_68_3_inst : DFF_X1 port map( D => n7984, CK => clk, Q => 
                           registers_68_3_port, QN => n16210);
   registers_reg_69_3_inst : DFF_X1 port map( D => n7983, CK => clk, Q => 
                           net226894, QN => n16206);
   registers_reg_70_3_inst : DFF_X1 port map( D => n7982, CK => clk, Q => 
                           net226893, QN => n16119);
   registers_reg_71_3_inst : DFF_X1 port map( D => n7981, CK => clk, Q => 
                           net226892, QN => n14980);
   out1_reg_3_inst : DFF_X1 port map( D => n7980, CK => clk, Q => out1(3), QN 
                           => net226891);
   registers_reg_4_2_inst : DFF_X1 port map( D => n7979, CK => clk, Q => 
                           registers_4_2_port, QN => n15523);
   registers_reg_5_2_inst : DFF_X1 port map( D => n7978, CK => clk, Q => 
                           registers_5_2_port, QN => n14715);
   registers_reg_6_2_inst : DFF_X1 port map( D => n7977, CK => clk, Q => 
                           net271259, QN => n12361);
   registers_reg_7_2_inst : DFF_X1 port map( D => n7976, CK => clk, Q => 
                           registers_7_2_port, QN => n15328);
   registers_reg_12_2_inst : DFF_X1 port map( D => n7975, CK => clk, Q => 
                           registers_12_2_port, QN => n15671);
   registers_reg_13_2_inst : DFF_X1 port map( D => n7974, CK => clk, Q => 
                           net226890, QN => n15076);
   registers_reg_14_2_inst : DFF_X1 port map( D => n7973, CK => clk, Q => 
                           net271258, QN => n11883);
   registers_reg_15_2_inst : DFF_X1 port map( D => n7972, CK => clk, Q => 
                           registers_15_2_port, QN => n15294);
   registers_reg_20_2_inst : DFF_X1 port map( D => n7971, CK => clk, Q => 
                           net271257, QN => n14833);
   registers_reg_21_2_inst : DFF_X1 port map( D => n7970, CK => clk, Q => 
                           net271256, QN => n12207);
   registers_reg_22_2_inst : DFF_X1 port map( D => n7969, CK => clk, Q => 
                           registers_22_2_port, QN => n15372);
   registers_reg_23_2_inst : DFF_X1 port map( D => n7968, CK => clk, Q => 
                           registers_23_2_port, QN => n15883);
   registers_reg_28_2_inst : DFF_X1 port map( D => n7967, CK => clk, Q => 
                           net226889, QN => n15006);
   registers_reg_29_2_inst : DFF_X1 port map( D => n7966, CK => clk, Q => 
                           registers_29_2_port, QN => n15794);
   registers_reg_30_2_inst : DFF_X1 port map( D => n7965, CK => clk, Q => 
                           registers_30_2_port, QN => n14680);
   registers_reg_31_2_inst : DFF_X1 port map( D => n7964, CK => clk, Q => 
                           net226888, QN => n15738);
   registers_reg_36_2_inst : DFF_X1 port map( D => n7963, CK => clk, Q => 
                           registers_36_2_port, QN => n15151);
   registers_reg_37_2_inst : DFF_X1 port map( D => n7962, CK => clk, Q => 
                           registers_37_2_port, QN => n14361);
   registers_reg_38_2_inst : DFF_X1 port map( D => n7961, CK => clk, Q => 
                           registers_38_2_port, QN => n15036);
   registers_reg_39_2_inst : DFF_X1 port map( D => n7960, CK => clk, Q => 
                           net271255, QN => n12173);
   registers_reg_44_2_inst : DFF_X1 port map( D => n7959, CK => clk, Q => 
                           registers_44_2_port, QN => n15468);
   registers_reg_45_2_inst : DFF_X1 port map( D => n7958, CK => clk, Q => 
                           registers_45_2_port, QN => n14776);
   registers_reg_46_2_inst : DFF_X1 port map( D => n7957, CK => clk, Q => 
                           net226887, QN => n11995);
   registers_reg_47_2_inst : DFF_X1 port map( D => n7956, CK => clk, Q => 
                           registers_47_2_port, QN => n14549);
   registers_reg_52_2_inst : DFF_X1 port map( D => n7955, CK => clk, Q => 
                           net226886, QN => n14940);
   registers_reg_53_2_inst : DFF_X1 port map( D => n7954, CK => clk, Q => 
                           net226885, QN => n15913);
   registers_reg_54_2_inst : DFF_X1 port map( D => n7953, CK => clk, Q => 
                           registers_54_2_port, QN => n14571);
   registers_reg_55_2_inst : DFF_X1 port map( D => n7952, CK => clk, Q => 
                           registers_55_2_port, QN => n12053);
   registers_reg_60_2_inst : DFF_X1 port map( D => n7951, CK => clk, Q => 
                           registers_60_2_port, QN => n14643);
   registers_reg_61_2_inst : DFF_X1 port map( D => n7950, CK => clk, Q => 
                           net226884, QN => n15578);
   registers_reg_62_2_inst : DFF_X1 port map( D => n7949, CK => clk, Q => 
                           registers_62_2_port, QN => n15125);
   registers_reg_63_2_inst : DFF_X1 port map( D => n7948, CK => clk, Q => 
                           registers_63_2_port, QN => n14508);
   registers_reg_0_2_inst : DFF_X1 port map( D => n7947, CK => clk, Q => 
                           registers_0_2_port, QN => n15797);
   registers_reg_1_2_inst : DFF_X1 port map( D => n7946, CK => clk, Q => 
                           registers_1_2_port, QN => n15581);
   registers_reg_2_2_inst : DFF_X1 port map( D => n7945, CK => clk, Q => 
                           registers_2_2_port, QN => n14775);
   registers_reg_3_2_inst : DFF_X1 port map( D => n7944, CK => clk, Q => 
                           net226883, QN => n15760);
   registers_reg_8_2_inst : DFF_X1 port map( D => n7943, CK => clk, Q => 
                           net226882, QN => n15212);
   registers_reg_9_2_inst : DFF_X1 port map( D => n7942, CK => clk, Q => 
                           registers_9_2_port, QN => n14331);
   registers_reg_10_2_inst : DFF_X1 port map( D => n7941, CK => clk, Q => 
                           registers_10_2_port, QN => n14716);
   registers_reg_11_2_inst : DFF_X1 port map( D => n7940, CK => clk, Q => 
                           registers_11_2_port, QN => n14430);
   registers_reg_16_2_inst : DFF_X1 port map( D => n7939, CK => clk, Q => 
                           registers_16_2_port, QN => n15701);
   registers_reg_17_2_inst : DFF_X1 port map( D => n7938, CK => clk, Q => 
                           registers_17_2_port, QN => n14607);
   registers_reg_18_2_inst : DFF_X1 port map( D => n7937, CK => clk, Q => 
                           registers_18_2_port, QN => n14364);
   registers_reg_19_2_inst : DFF_X1 port map( D => n7936, CK => clk, Q => 
                           registers_19_2_port, QN => n15804);
   registers_reg_24_2_inst : DFF_X1 port map( D => n7935, CK => clk, Q => 
                           net226881, QN => n15183);
   registers_reg_25_2_inst : DFF_X1 port map( D => n7934, CK => clk, Q => 
                           registers_25_2_port, QN => n14302);
   registers_reg_26_2_inst : DFF_X1 port map( D => n7933, CK => clk, Q => 
                           net271254, QN => n12360);
   registers_reg_27_2_inst : DFF_X1 port map( D => n7932, CK => clk, Q => 
                           net271253, QN => n12020);
   registers_reg_32_2_inst : DFF_X1 port map( D => n7931, CK => clk, Q => 
                           net271252, QN => n12311);
   registers_reg_33_2_inst : DFF_X1 port map( D => n7930, CK => clk, Q => 
                           net271251, QN => n11799);
   registers_reg_34_2_inst : DFF_X1 port map( D => n7929, CK => clk, Q => 
                           registers_34_2_port, QN => n15497);
   registers_reg_35_2_inst : DFF_X1 port map( D => n7928, CK => clk, Q => 
                           net226880, QN => n15586);
   registers_reg_40_2_inst : DFF_X1 port map( D => n7927, CK => clk, Q => 
                           registers_40_2_port, QN => n15077);
   registers_reg_41_2_inst : DFF_X1 port map( D => n7926, CK => clk, Q => 
                           registers_41_2_port, QN => n14431);
   registers_reg_42_2_inst : DFF_X1 port map( D => n7925, CK => clk, Q => 
                           registers_42_2_port, QN => n15922);
   registers_reg_43_2_inst : DFF_X1 port map( D => n7924, CK => clk, Q => 
                           registers_43_2_port, QN => n14890);
   registers_reg_48_2_inst : DFF_X1 port map( D => n7923, CK => clk, Q => 
                           registers_48_2_port, QN => n15554);
   registers_reg_49_2_inst : DFF_X1 port map( D => n7922, CK => clk, Q => 
                           registers_49_2_port, QN => n14486);
   registers_reg_50_2_inst : DFF_X1 port map( D => n7921, CK => clk, Q => 
                           registers_50_2_port, QN => n15971);
   registers_reg_51_2_inst : DFF_X1 port map( D => n7920, CK => clk, Q => 
                           registers_51_2_port, QN => n15401);
   registers_reg_56_2_inst : DFF_X1 port map( D => n7919, CK => clk, Q => 
                           registers_56_2_port, QN => n16000);
   registers_reg_57_2_inst : DFF_X1 port map( D => n7918, CK => clk, Q => 
                           net226879, QN => n15244);
   registers_reg_58_2_inst : DFF_X1 port map( D => n7917, CK => clk, Q => 
                           net226878, QN => n14912);
   registers_reg_59_2_inst : DFF_X1 port map( D => n7916, CK => clk, Q => 
                           registers_59_2_port, QN => n15434);
   to_mem_reg_2_inst : DFF_X1 port map( D => n7915, CK => clk, Q => net271250, 
                           QN => n7723);
   registers_reg_64_2_inst : DFF_X1 port map( D => n7914, CK => clk, Q => 
                           net226877, QN => n16203);
   registers_reg_65_2_inst : DFF_X1 port map( D => n7913, CK => clk, Q => 
                           net226876, QN => n16113);
   registers_reg_66_2_inst : DFF_X1 port map( D => n7912, CK => clk, Q => 
                           net226875, QN => n16121);
   registers_reg_67_2_inst : DFF_X1 port map( D => n7911, CK => clk, Q => 
                           net271249, QN => n14286);
   registers_reg_68_2_inst : DFF_X1 port map( D => n7910, CK => clk, Q => 
                           registers_68_2_port, QN => n16207);
   registers_reg_69_2_inst : DFF_X1 port map( D => n7909, CK => clk, Q => 
                           net226874, QN => n16200);
   registers_reg_70_2_inst : DFF_X1 port map( D => n7908, CK => clk, Q => 
                           net226873, QN => n16117);
   registers_reg_71_2_inst : DFF_X1 port map( D => n7907, CK => clk, Q => 
                           net226872, QN => n14962);
   out1_reg_2_inst : DFF_X1 port map( D => n7906, CK => clk, Q => out1(2), QN 
                           => net226871);
   registers_reg_2_1_inst : DFF_X1 port map( D => n7905, CK => clk, Q => 
                           registers_2_1_port, QN => n14773);
   registers_reg_3_1_inst : DFF_X1 port map( D => n7904, CK => clk, Q => 
                           net226870, QN => n15759);
   registers_reg_6_1_inst : DFF_X1 port map( D => n7903, CK => clk, Q => 
                           net271248, QN => n12359);
   registers_reg_7_1_inst : DFF_X1 port map( D => n7902, CK => clk, Q => 
                           registers_7_1_port, QN => n15327);
   registers_reg_10_1_inst : DFF_X1 port map( D => n7901, CK => clk, Q => 
                           registers_10_1_port, QN => n14714);
   registers_reg_11_1_inst : DFF_X1 port map( D => n7900, CK => clk, Q => 
                           registers_11_1_port, QN => n14428);
   registers_reg_14_1_inst : DFF_X1 port map( D => n7899, CK => clk, Q => 
                           net271247, QN => n11882);
   registers_reg_15_1_inst : DFF_X1 port map( D => n7898, CK => clk, Q => 
                           registers_15_1_port, QN => n15293);
   registers_reg_18_1_inst : DFF_X1 port map( D => n7897, CK => clk, Q => 
                           registers_18_1_port, QN => n14360);
   registers_reg_19_1_inst : DFF_X1 port map( D => n7896, CK => clk, Q => 
                           registers_19_1_port, QN => n15793);
   registers_reg_22_1_inst : DFF_X1 port map( D => n7895, CK => clk, Q => 
                           registers_22_1_port, QN => n15371);
   registers_reg_23_1_inst : DFF_X1 port map( D => n7894, CK => clk, Q => 
                           registers_23_1_port, QN => n15882);
   registers_reg_26_1_inst : DFF_X1 port map( D => n7893, CK => clk, Q => 
                           net271246, QN => n12358);
   registers_reg_27_1_inst : DFF_X1 port map( D => n7892, CK => clk, Q => 
                           net271245, QN => n12019);
   registers_reg_30_1_inst : DFF_X1 port map( D => n7891, CK => clk, Q => 
                           registers_30_1_port, QN => n14679);
   registers_reg_31_1_inst : DFF_X1 port map( D => n7890, CK => clk, Q => 
                           net226869, QN => n15737);
   registers_reg_34_1_inst : DFF_X1 port map( D => n7889, CK => clk, Q => 
                           registers_34_1_port, QN => n15496);
   registers_reg_35_1_inst : DFF_X1 port map( D => n7888, CK => clk, Q => 
                           net226868, QN => n15577);
   registers_reg_38_1_inst : DFF_X1 port map( D => n7887, CK => clk, Q => 
                           registers_38_1_port, QN => n15035);
   registers_reg_39_1_inst : DFF_X1 port map( D => n7886, CK => clk, Q => 
                           net271244, QN => n12172);
   registers_reg_42_1_inst : DFF_X1 port map( D => n7885, CK => clk, Q => 
                           registers_42_1_port, QN => n15912);
   registers_reg_43_1_inst : DFF_X1 port map( D => n7884, CK => clk, Q => 
                           registers_43_1_port, QN => n14889);
   registers_reg_46_1_inst : DFF_X1 port map( D => n7883, CK => clk, Q => 
                           net226867, QN => n11952);
   registers_reg_47_1_inst : DFF_X1 port map( D => n7882, CK => clk, Q => 
                           registers_47_1_port, QN => n14548);
   registers_reg_50_1_inst : DFF_X1 port map( D => n7881, CK => clk, Q => 
                           registers_50_1_port, QN => n15969);
   registers_reg_51_1_inst : DFF_X1 port map( D => n7880, CK => clk, Q => 
                           registers_51_1_port, QN => n15370);
   registers_reg_54_1_inst : DFF_X1 port map( D => n7879, CK => clk, Q => 
                           registers_54_1_port, QN => n14570);
   registers_reg_55_1_inst : DFF_X1 port map( D => n7878, CK => clk, Q => 
                           registers_55_1_port, QN => n12052);
   registers_reg_58_1_inst : DFF_X1 port map( D => n7877, CK => clk, Q => 
                           net226866, QN => n14911);
   registers_reg_59_1_inst : DFF_X1 port map( D => n7876, CK => clk, Q => 
                           registers_59_1_port, QN => n15433);
   registers_reg_62_1_inst : DFF_X1 port map( D => n7875, CK => clk, Q => 
                           registers_62_1_port, QN => n15124);
   registers_reg_63_1_inst : DFF_X1 port map( D => n7874, CK => clk, Q => 
                           registers_63_1_port, QN => n14507);
   registers_reg_66_1_inst : DFF_X1 port map( D => n7873, CK => clk, Q => 
                           net226865, QN => n16116);
   registers_reg_67_1_inst : DFF_X1 port map( D => n7872, CK => clk, Q => 
                           net271243, QN => n14285);
   registers_reg_0_1_inst : DFF_X1 port map( D => n7871, CK => clk, Q => 
                           registers_0_1_port, QN => n15796);
   registers_reg_1_1_inst : DFF_X1 port map( D => n7870, CK => clk, Q => 
                           registers_1_1_port, QN => n15580);
   registers_reg_4_1_inst : DFF_X1 port map( D => n7869, CK => clk, Q => 
                           registers_4_1_port, QN => n15522);
   registers_reg_5_1_inst : DFF_X1 port map( D => n7868, CK => clk, Q => 
                           registers_5_1_port, QN => n14713);
   registers_reg_8_1_inst : DFF_X1 port map( D => n7867, CK => clk, Q => 
                           net226864, QN => n15211);
   registers_reg_9_1_inst : DFF_X1 port map( D => n7866, CK => clk, Q => 
                           registers_9_1_port, QN => n14330);
   registers_reg_12_1_inst : DFF_X1 port map( D => n7865, CK => clk, Q => 
                           registers_12_1_port, QN => n15670);
   registers_reg_13_1_inst : DFF_X1 port map( D => n7864, CK => clk, Q => 
                           net226863, QN => n15074);
   registers_reg_16_1_inst : DFF_X1 port map( D => n7863, CK => clk, Q => 
                           registers_16_1_port, QN => n15700);
   registers_reg_17_1_inst : DFF_X1 port map( D => n7862, CK => clk, Q => 
                           registers_17_1_port, QN => n14606);
   registers_reg_20_1_inst : DFF_X1 port map( D => n7861, CK => clk, Q => 
                           net271242, QN => n14832);
   registers_reg_21_1_inst : DFF_X1 port map( D => n7860, CK => clk, Q => 
                           net271241, QN => n12206);
   registers_reg_24_1_inst : DFF_X1 port map( D => n7859, CK => clk, Q => 
                           net226862, QN => n15182);
   registers_reg_25_1_inst : DFF_X1 port map( D => n7858, CK => clk, Q => 
                           registers_25_1_port, QN => n14301);
   registers_reg_28_1_inst : DFF_X1 port map( D => n7857, CK => clk, Q => 
                           net226861, QN => n15005);
   registers_reg_29_1_inst : DFF_X1 port map( D => n7856, CK => clk, Q => 
                           registers_29_1_port, QN => n15803);
   registers_reg_32_1_inst : DFF_X1 port map( D => n7855, CK => clk, Q => 
                           net271240, QN => n12310);
   registers_reg_33_1_inst : DFF_X1 port map( D => n7854, CK => clk, Q => 
                           net271239, QN => n11756);
   registers_reg_36_1_inst : DFF_X1 port map( D => n7853, CK => clk, Q => 
                           registers_36_1_port, QN => n15153);
   registers_reg_37_1_inst : DFF_X1 port map( D => n7852, CK => clk, Q => 
                           registers_37_1_port, QN => n14363);
   registers_reg_40_1_inst : DFF_X1 port map( D => n7851, CK => clk, Q => 
                           registers_40_1_port, QN => n15075);
   registers_reg_41_1_inst : DFF_X1 port map( D => n7850, CK => clk, Q => 
                           registers_41_1_port, QN => n14429);
   registers_reg_44_1_inst : DFF_X1 port map( D => n7849, CK => clk, Q => 
                           registers_44_1_port, QN => n15467);
   registers_reg_45_1_inst : DFF_X1 port map( D => n7848, CK => clk, Q => 
                           registers_45_1_port, QN => n14774);
   registers_reg_48_1_inst : DFF_X1 port map( D => n7847, CK => clk, Q => 
                           registers_48_1_port, QN => n15553);
   registers_reg_49_1_inst : DFF_X1 port map( D => n7846, CK => clk, Q => 
                           registers_49_1_port, QN => n14485);
   registers_reg_52_1_inst : DFF_X1 port map( D => n7845, CK => clk, Q => 
                           net226860, QN => n14939);
   registers_reg_53_1_inst : DFF_X1 port map( D => n7844, CK => clk, Q => 
                           net226859, QN => n15914);
   registers_reg_56_1_inst : DFF_X1 port map( D => n7843, CK => clk, Q => 
                           registers_56_1_port, QN => n15999);
   registers_reg_57_1_inst : DFF_X1 port map( D => n7842, CK => clk, Q => 
                           net226858, QN => n15243);
   registers_reg_60_1_inst : DFF_X1 port map( D => n7841, CK => clk, Q => 
                           registers_60_1_port, QN => n14645);
   registers_reg_61_1_inst : DFF_X1 port map( D => n7840, CK => clk, Q => 
                           net226857, QN => n15661);
   to_mem_reg_1_inst : DFF_X1 port map( D => n7839, CK => clk, Q => net271238, 
                           QN => n7724);
   registers_reg_64_1_inst : DFF_X1 port map( D => n7838, CK => clk, Q => 
                           net226856, QN => n16202);
   registers_reg_65_1_inst : DFF_X1 port map( D => n7837, CK => clk, Q => 
                           net226855, QN => n16112);
   registers_reg_68_1_inst : DFF_X1 port map( D => n7836, CK => clk, Q => 
                           registers_68_1_port, QN => n16209);
   registers_reg_69_1_inst : DFF_X1 port map( D => n7835, CK => clk, Q => 
                           net226854, QN => n16205);
   registers_reg_70_1_inst : DFF_X1 port map( D => n7834, CK => clk, Q => 
                           net226853, QN => n16115);
   registers_reg_71_1_inst : DFF_X1 port map( D => n7833, CK => clk, Q => 
                           net226852, QN => n14961);
   out1_reg_1_inst : DFF_X1 port map( D => n7832, CK => clk, Q => out1(1), QN 
                           => net226851);
   registers_reg_1_0_inst : DFF_X1 port map( D => n7831, CK => clk, Q => 
                           registers_1_0_port, QN => n15576);
   registers_reg_3_0_inst : DFF_X1 port map( D => n7830, CK => clk, Q => 
                           net226850, QN => n15758);
   registers_reg_5_0_inst : DFF_X1 port map( D => n7829, CK => clk, Q => 
                           registers_5_0_port, QN => n14711);
   registers_reg_7_0_inst : DFF_X1 port map( D => n7828, CK => clk, Q => 
                           registers_7_0_port, QN => n15326);
   registers_reg_9_0_inst : DFF_X1 port map( D => n7827, CK => clk, Q => 
                           registers_9_0_port, QN => n14329);
   registers_reg_11_0_inst : DFF_X1 port map( D => n7826, CK => clk, Q => 
                           registers_11_0_port, QN => n14426);
   registers_reg_13_0_inst : DFF_X1 port map( D => n7825, CK => clk, Q => 
                           net226849, QN => n15072);
   registers_reg_15_0_inst : DFF_X1 port map( D => n7824, CK => clk, Q => 
                           registers_15_0_port, QN => n15292);
   registers_reg_17_0_inst : DFF_X1 port map( D => n7823, CK => clk, Q => 
                           registers_17_0_port, QN => n14605);
   registers_reg_19_0_inst : DFF_X1 port map( D => n7822, CK => clk, Q => 
                           registers_19_0_port, QN => n15792);
   registers_reg_21_0_inst : DFF_X1 port map( D => n7821, CK => clk, Q => 
                           net271237, QN => n12205);
   registers_reg_23_0_inst : DFF_X1 port map( D => n7820, CK => clk, Q => 
                           registers_23_0_port, QN => n15881);
   registers_reg_25_0_inst : DFF_X1 port map( D => n7819, CK => clk, Q => 
                           registers_25_0_port, QN => n14300);
   registers_reg_27_0_inst : DFF_X1 port map( D => n7818, CK => clk, Q => 
                           net271236, QN => n12018);
   registers_reg_29_0_inst : DFF_X1 port map( D => n7817, CK => clk, Q => 
                           registers_29_0_port, QN => n15791);
   registers_reg_31_0_inst : DFF_X1 port map( D => n7816, CK => clk, Q => 
                           net226848, QN => n15736);
   registers_reg_33_0_inst : DFF_X1 port map( D => n7815, CK => clk, Q => 
                           net271235, QN => n11713);
   registers_reg_35_0_inst : DFF_X1 port map( D => n7814, CK => clk, Q => 
                           net226847, QN => n15575);
   registers_reg_37_0_inst : DFF_X1 port map( D => n7813, CK => clk, Q => 
                           registers_37_0_port, QN => n14359);
   registers_reg_39_0_inst : DFF_X1 port map( D => n7812, CK => clk, Q => 
                           net271234, QN => n12171);
   registers_reg_41_0_inst : DFF_X1 port map( D => n7811, CK => clk, Q => 
                           registers_41_0_port, QN => n14427);
   registers_reg_43_0_inst : DFF_X1 port map( D => n7810, CK => clk, Q => 
                           registers_43_0_port, QN => n14888);
   registers_reg_45_0_inst : DFF_X1 port map( D => n7809, CK => clk, Q => 
                           registers_45_0_port, QN => n14772);
   registers_reg_47_0_inst : DFF_X1 port map( D => n7808, CK => clk, Q => 
                           registers_47_0_port, QN => n14547);
   registers_reg_49_0_inst : DFF_X1 port map( D => n7807, CK => clk, Q => 
                           registers_49_0_port, QN => n14484);
   registers_reg_51_0_inst : DFF_X1 port map( D => n7806, CK => clk, Q => 
                           registers_51_0_port, QN => n15369);
   registers_reg_53_0_inst : DFF_X1 port map( D => n7805, CK => clk, Q => 
                           net226846, QN => n15911);
   registers_reg_55_0_inst : DFF_X1 port map( D => n7804, CK => clk, Q => 
                           registers_55_0_port, QN => n12055);
   registers_reg_57_0_inst : DFF_X1 port map( D => n7803, CK => clk, Q => 
                           net226845, QN => n15245);
   registers_reg_59_0_inst : DFF_X1 port map( D => n7802, CK => clk, Q => 
                           registers_59_0_port, QN => n15432);
   registers_reg_61_0_inst : DFF_X1 port map( D => n7801, CK => clk, Q => 
                           net226844, QN => n15574);
   registers_reg_63_0_inst : DFF_X1 port map( D => n7800, CK => clk, Q => 
                           registers_63_0_port, QN => n14506);
   registers_reg_65_0_inst : DFF_X1 port map( D => n7799, CK => clk, Q => 
                           net226843, QN => n16111);
   registers_reg_67_0_inst : DFF_X1 port map( D => n7798, CK => clk, Q => 
                           net271233, QN => n14284);
   registers_reg_69_0_inst : DFF_X1 port map( D => n7797, CK => clk, Q => 
                           net226842, QN => n16199);
   registers_reg_0_0_inst : DFF_X1 port map( D => n7796, CK => clk, Q => 
                           registers_0_0_port, QN => n15795);
   registers_reg_2_0_inst : DFF_X1 port map( D => n7795, CK => clk, Q => 
                           registers_2_0_port, QN => n14771);
   registers_reg_4_0_inst : DFF_X1 port map( D => n7794, CK => clk, Q => 
                           registers_4_0_port, QN => n15521);
   registers_reg_6_0_inst : DFF_X1 port map( D => n7793, CK => clk, Q => 
                           net271232, QN => n12357);
   registers_reg_8_0_inst : DFF_X1 port map( D => n7792, CK => clk, Q => 
                           net226841, QN => n15210);
   registers_reg_10_0_inst : DFF_X1 port map( D => n7791, CK => clk, Q => 
                           registers_10_0_port, QN => n14712);
   registers_reg_12_0_inst : DFF_X1 port map( D => n7790, CK => clk, Q => 
                           registers_12_0_port, QN => n15669);
   registers_reg_14_0_inst : DFF_X1 port map( D => n7789, CK => clk, Q => 
                           net271231, QN => n11881);
   registers_reg_16_0_inst : DFF_X1 port map( D => n7788, CK => clk, Q => 
                           registers_16_0_port, QN => n15699);
   registers_reg_18_0_inst : DFF_X1 port map( D => n7787, CK => clk, Q => 
                           registers_18_0_port, QN => n14362);
   registers_reg_20_0_inst : DFF_X1 port map( D => n7786, CK => clk, Q => 
                           net271230, QN => n14831);
   registers_reg_22_0_inst : DFF_X1 port map( D => n7785, CK => clk, Q => 
                           registers_22_0_port, QN => n15373);
   registers_reg_24_0_inst : DFF_X1 port map( D => n7784, CK => clk, Q => 
                           net226840, QN => n15181);
   registers_reg_26_0_inst : DFF_X1 port map( D => n7783, CK => clk, Q => 
                           net271229, QN => n12356);
   registers_reg_28_0_inst : DFF_X1 port map( D => n7782, CK => clk, Q => 
                           net226839, QN => n15004);
   registers_reg_30_0_inst : DFF_X1 port map( D => n7781, CK => clk, Q => 
                           registers_30_0_port, QN => n14678);
   registers_reg_32_0_inst : DFF_X1 port map( D => n7780, CK => clk, Q => 
                           net271228, QN => n12309);
   registers_reg_34_0_inst : DFF_X1 port map( D => n7779, CK => clk, Q => 
                           registers_34_0_port, QN => n15495);
   registers_reg_36_0_inst : DFF_X1 port map( D => n7778, CK => clk, Q => 
                           registers_36_0_port, QN => n15152);
   registers_reg_38_0_inst : DFF_X1 port map( D => n7777, CK => clk, Q => 
                           registers_38_0_port, QN => n15037);
   registers_reg_40_0_inst : DFF_X1 port map( D => n7776, CK => clk, Q => 
                           registers_40_0_port, QN => n15073);
   registers_reg_42_0_inst : DFF_X1 port map( D => n7775, CK => clk, Q => 
                           registers_42_0_port, QN => n15921);
   registers_reg_44_0_inst : DFF_X1 port map( D => n7774, CK => clk, Q => 
                           registers_44_0_port, QN => n15466);
   registers_reg_46_0_inst : DFF_X1 port map( D => n7773, CK => clk, Q => 
                           net226838, QN => n11951);
   registers_reg_48_0_inst : DFF_X1 port map( D => n7772, CK => clk, Q => 
                           registers_48_0_port, QN => n15552);
   registers_reg_50_0_inst : DFF_X1 port map( D => n7771, CK => clk, Q => 
                           registers_50_0_port, QN => n15970);
   registers_reg_52_0_inst : DFF_X1 port map( D => n7770, CK => clk, Q => 
                           net226837, QN => n14938);
   registers_reg_54_0_inst : DFF_X1 port map( D => n7769, CK => clk, Q => 
                           registers_54_0_port, QN => n14573);
   registers_reg_56_0_inst : DFF_X1 port map( D => n7768, CK => clk, Q => 
                           registers_56_0_port, QN => n15998);
   registers_reg_58_0_inst : DFF_X1 port map( D => n7767, CK => clk, Q => 
                           net226836, QN => n14910);
   registers_reg_60_0_inst : DFF_X1 port map( D => n7766, CK => clk, Q => 
                           registers_60_0_port, QN => n14669);
   registers_reg_62_0_inst : DFF_X1 port map( D => n7765, CK => clk, Q => 
                           registers_62_0_port, QN => n15123);
   to_mem_reg_0_inst : DFF_X1 port map( D => n7764, CK => clk, Q => net271227, 
                           QN => n7725);
   registers_reg_64_0_inst : DFF_X1 port map( D => n7763, CK => clk, Q => 
                           net226835, QN => n16201);
   registers_reg_66_0_inst : DFF_X1 port map( D => n7762, CK => clk, Q => 
                           net226834, QN => n16120);
   registers_reg_68_0_inst : DFF_X1 port map( D => n7761, CK => clk, Q => 
                           registers_68_0_port, QN => n16208);
   registers_reg_70_0_inst : DFF_X1 port map( D => n7760, CK => clk, Q => 
                           net226833, QN => n16118);
   registers_reg_71_0_inst : DFF_X1 port map( D => n7759, CK => clk, Q => 
                           net226832, QN => n14960);
   out1_reg_0_inst : DFF_X1 port map( D => n7758, CK => clk, Q => out1(0), QN 
                           => net226831);
   out2_reg_31_inst : DFF_X1 port map( D => n7757, CK => clk, Q => out2(31), QN
                           => net226830);
   out2_reg_30_inst : DFF_X1 port map( D => n7756, CK => clk, Q => out2(30), QN
                           => net226829);
   out2_reg_29_inst : DFF_X1 port map( D => n7755, CK => clk, Q => out2(29), QN
                           => net226828);
   out2_reg_28_inst : DFF_X1 port map( D => n7754, CK => clk, Q => out2(28), QN
                           => net226827);
   out2_reg_27_inst : DFF_X1 port map( D => n7753, CK => clk, Q => out2(27), QN
                           => net226826);
   out2_reg_26_inst : DFF_X1 port map( D => n7752, CK => clk, Q => out2(26), QN
                           => net226825);
   out2_reg_25_inst : DFF_X1 port map( D => n7751, CK => clk, Q => out2(25), QN
                           => net226824);
   out2_reg_24_inst : DFF_X1 port map( D => n7750, CK => clk, Q => out2(24), QN
                           => net226823);
   out2_reg_23_inst : DFF_X1 port map( D => n7749, CK => clk, Q => out2(23), QN
                           => net226822);
   out2_reg_22_inst : DFF_X1 port map( D => n7748, CK => clk, Q => out2(22), QN
                           => net226821);
   out2_reg_21_inst : DFF_X1 port map( D => n7747, CK => clk, Q => out2(21), QN
                           => net226820);
   out2_reg_20_inst : DFF_X1 port map( D => n7746, CK => clk, Q => out2(20), QN
                           => net226819);
   out2_reg_19_inst : DFF_X1 port map( D => n7745, CK => clk, Q => out2(19), QN
                           => net226818);
   out2_reg_18_inst : DFF_X1 port map( D => n7744, CK => clk, Q => out2(18), QN
                           => net226817);
   out2_reg_17_inst : DFF_X1 port map( D => n7743, CK => clk, Q => out2(17), QN
                           => net226816);
   out2_reg_16_inst : DFF_X1 port map( D => n7742, CK => clk, Q => out2(16), QN
                           => net226815);
   out2_reg_15_inst : DFF_X1 port map( D => n7741, CK => clk, Q => out2(15), QN
                           => net226814);
   out2_reg_14_inst : DFF_X1 port map( D => n7740, CK => clk, Q => out2(14), QN
                           => net226813);
   out2_reg_13_inst : DFF_X1 port map( D => n7739, CK => clk, Q => out2(13), QN
                           => net226812);
   out2_reg_12_inst : DFF_X1 port map( D => n7738, CK => clk, Q => out2(12), QN
                           => net226811);
   out2_reg_11_inst : DFF_X1 port map( D => n7737, CK => clk, Q => out2(11), QN
                           => net226810);
   out2_reg_10_inst : DFF_X1 port map( D => n7736, CK => clk, Q => out2(10), QN
                           => net226809);
   out2_reg_9_inst : DFF_X1 port map( D => n7735, CK => clk, Q => out2(9), QN 
                           => net226808);
   out2_reg_8_inst : DFF_X1 port map( D => n7734, CK => clk, Q => out2(8), QN 
                           => net226807);
   out2_reg_7_inst : DFF_X1 port map( D => n7733, CK => clk, Q => out2(7), QN 
                           => net226806);
   out2_reg_6_inst : DFF_X1 port map( D => n7732, CK => clk, Q => out2(6), QN 
                           => net226805);
   out2_reg_5_inst : DFF_X1 port map( D => n7731, CK => clk, Q => out2(5), QN 
                           => net226804);
   out2_reg_4_inst : DFF_X1 port map( D => n7730, CK => clk, Q => out2(4), QN 
                           => net226803);
   out2_reg_3_inst : DFF_X1 port map( D => n7729, CK => clk, Q => out2(3), QN 
                           => net226802);
   out2_reg_2_inst : DFF_X1 port map( D => n7728, CK => clk, Q => out2(2), QN 
                           => net226801);
   out2_reg_1_inst : DFF_X1 port map( D => n7727, CK => clk, Q => out2(1), QN 
                           => net226800);
   out2_reg_0_inst : DFF_X1 port map( D => n7726, CK => clk, Q => out2(0), QN 
                           => net226799);
   add_73_U1_1 : FA_X1 port map( A => add_wr(1), B => lastcwp_1_port, CI => 
                           add_73_carry_1_port, CO => add_73_carry_2_port, S =>
                           N273);
   add_73_U1_2 : FA_X1 port map( A => add_wr(2), B => lastcwp_2_port, CI => 
                           add_73_carry_2_port, CO => add_73_carry_3_port, S =>
                           N274);
   add_73_U1_3 : FA_X1 port map( A => add_wr(3), B => lastcwp_3_port, CI => 
                           add_73_carry_3_port, CO => add_73_carry_4_port, S =>
                           N275);
   add_73_U1_4 : FA_X1 port map( A => add_wr(4), B => lastcwp_4_port, CI => 
                           add_73_carry_4_port, CO => add_73_carry_5_port, S =>
                           N276);
   cwp_reg_3_inst : DFF_X1 port map( D => n10175, CK => clk, Q => N9910, QN => 
                           n10187);
   cwp_reg_2_inst : DFF_X1 port map( D => n10177, CK => clk, Q => N9909, QN => 
                           n10188);
   cwp_reg_1_inst : DFF_X1 port map( D => n10179, CK => clk, Q => N9908, QN => 
                           n10189);
   cwp_reg_0_inst : DFF_X1 port map( D => n10180, CK => clk, Q => N9641, QN => 
                           n10190);
   n4 <= '0';
   n76 <= '0';
   n77 <= '0';
   U8886 : NOR4_X2 port map( A1 => n14173, A2 => N9924, A3 => N9926, A4 => call
                           , ZN => n14105);
   U8949 : NOR4_X2 port map( A1 => N9922, A2 => N9924, A3 => N9926, A4 => call,
                           ZN => n14095);
   U9269 : NAND3_X1 port map( A1 => n10513, A2 => n10514, A3 => n10515, ZN => 
                           n8108);
   U9270 : NAND3_X1 port map( A1 => n10665, A2 => n10666, A3 => n10667, ZN => 
                           n8106);
   U9271 : NAND3_X1 port map( A1 => n10724, A2 => n10725, A3 => n10726, ZN => 
                           n8104);
   U9272 : NAND3_X1 port map( A1 => n10767, A2 => n10768, A3 => n10769, ZN => 
                           n8102);
   U9273 : NAND3_X1 port map( A1 => n10810, A2 => n10811, A3 => n10812, ZN => 
                           n8100);
   U9274 : NAND3_X1 port map( A1 => n10853, A2 => n10854, A3 => n10855, ZN => 
                           n8098);
   U9275 : NAND3_X1 port map( A1 => n10896, A2 => n10897, A3 => n10898, ZN => 
                           n8096);
   U9276 : NAND3_X1 port map( A1 => n10939, A2 => n10940, A3 => n10941, ZN => 
                           n8094);
   U9277 : NAND3_X1 port map( A1 => n10982, A2 => n10983, A3 => n10984, ZN => 
                           n8092);
   U9278 : NAND3_X1 port map( A1 => n11025, A2 => n11026, A3 => n11027, ZN => 
                           n8090);
   U9279 : NAND3_X1 port map( A1 => n11068, A2 => n11069, A3 => n11070, ZN => 
                           n8088);
   U9280 : NAND3_X1 port map( A1 => n11111, A2 => n11112, A3 => n11113, ZN => 
                           n8086);
   U9281 : NAND3_X1 port map( A1 => n11154, A2 => n11155, A3 => n11156, ZN => 
                           n8084);
   U9282 : NAND3_X1 port map( A1 => n11197, A2 => n11198, A3 => n11199, ZN => 
                           n8082);
   U9283 : NAND3_X1 port map( A1 => n11240, A2 => n11241, A3 => n11242, ZN => 
                           n8080);
   U9284 : NAND3_X1 port map( A1 => n11283, A2 => n11284, A3 => n11285, ZN => 
                           n8078);
   U9285 : NAND3_X1 port map( A1 => n11326, A2 => n11327, A3 => n11328, ZN => 
                           n8076);
   U9286 : NAND3_X1 port map( A1 => n11369, A2 => n11370, A3 => n11371, ZN => 
                           n8074);
   U9287 : NAND3_X1 port map( A1 => n11412, A2 => n11413, A3 => n11414, ZN => 
                           n8072);
   U9288 : NAND3_X1 port map( A1 => n11455, A2 => n11456, A3 => n11457, ZN => 
                           n8070);
   U9289 : NAND3_X1 port map( A1 => n11499, A2 => n11500, A3 => n11501, ZN => 
                           n8068);
   U9290 : NAND3_X1 port map( A1 => n11542, A2 => n11543, A3 => n11544, ZN => 
                           n8066);
   U9291 : NAND3_X1 port map( A1 => n11585, A2 => n11586, A3 => n11587, ZN => 
                           n8064);
   U9292 : NAND3_X1 port map( A1 => n11628, A2 => n11629, A3 => n11630, ZN => 
                           n8062);
   U9293 : NAND3_X1 port map( A1 => n11671, A2 => n11672, A3 => n11673, ZN => 
                           n8060);
   U9294 : NAND3_X1 port map( A1 => n11714, A2 => n11715, A3 => n11716, ZN => 
                           n8058);
   U9295 : NAND3_X1 port map( A1 => n11757, A2 => n11758, A3 => n11759, ZN => 
                           n8056);
   U9296 : NAND3_X1 port map( A1 => n11800, A2 => n11801, A3 => n11802, ZN => 
                           n8054);
   U9297 : NAND3_X1 port map( A1 => n11953, A2 => n11954, A3 => n11955, ZN => 
                           n7980);
   U9298 : NAND3_X1 port map( A1 => n12106, A2 => n12107, A3 => n12108, ZN => 
                           n7906);
   U9299 : NAND3_X1 port map( A1 => n12259, A2 => n12260, A3 => n12261, ZN => 
                           n7832);
   U9300 : NAND3_X1 port map( A1 => n12416, A2 => n12417, A3 => n12418, ZN => 
                           n7758);
   U9301 : XOR2_X1 port map( A => add_wr(3), B => add_rd1(3), Z => n12515);
   U9302 : NAND3_X1 port map( A1 => enable, A2 => n18044, A3 => rd1, ZN => 
                           n10525);
   U9303 : NAND3_X1 port map( A1 => n12516, A2 => n12517, A3 => n12518, ZN => 
                           n7757);
   U9304 : NAND3_X1 port map( A1 => n12635, A2 => n12636, A3 => n12637, ZN => 
                           n7756);
   U9305 : NAND3_X1 port map( A1 => n12679, A2 => n12680, A3 => n12681, ZN => 
                           n7755);
   U9306 : NAND3_X1 port map( A1 => n12721, A2 => n12722, A3 => n12723, ZN => 
                           n7754);
   U9307 : NAND3_X1 port map( A1 => n12763, A2 => n12764, A3 => n12765, ZN => 
                           n7753);
   U9308 : NAND3_X1 port map( A1 => n12805, A2 => n12806, A3 => n12807, ZN => 
                           n7752);
   U9309 : NAND3_X1 port map( A1 => n12847, A2 => n12848, A3 => n12849, ZN => 
                           n7751);
   U9310 : NAND3_X1 port map( A1 => n12889, A2 => n12890, A3 => n12891, ZN => 
                           n7750);
   U9311 : NAND3_X1 port map( A1 => n12931, A2 => n12932, A3 => n12933, ZN => 
                           n7749);
   U9312 : NAND3_X1 port map( A1 => n12973, A2 => n12974, A3 => n12975, ZN => 
                           n7748);
   U9313 : NAND3_X1 port map( A1 => n13015, A2 => n13016, A3 => n13017, ZN => 
                           n7747);
   U9314 : NAND3_X1 port map( A1 => n13057, A2 => n13058, A3 => n13059, ZN => 
                           n7746);
   U9315 : NAND3_X1 port map( A1 => n13099, A2 => n13100, A3 => n13101, ZN => 
                           n7745);
   U9316 : NAND3_X1 port map( A1 => n13141, A2 => n13142, A3 => n13143, ZN => 
                           n7744);
   U9317 : NAND3_X1 port map( A1 => n13183, A2 => n13184, A3 => n13185, ZN => 
                           n7743);
   U9318 : NAND3_X1 port map( A1 => n13225, A2 => n13226, A3 => n13227, ZN => 
                           n7742);
   U9319 : NAND3_X1 port map( A1 => n13267, A2 => n13268, A3 => n13269, ZN => 
                           n7741);
   U9320 : NAND3_X1 port map( A1 => n13309, A2 => n13310, A3 => n13311, ZN => 
                           n7740);
   U9321 : NAND3_X1 port map( A1 => n13351, A2 => n13352, A3 => n13353, ZN => 
                           n7739);
   U9322 : NAND3_X1 port map( A1 => n13393, A2 => n13394, A3 => n13395, ZN => 
                           n7738);
   U9323 : NAND3_X1 port map( A1 => n13435, A2 => n13436, A3 => n13437, ZN => 
                           n7737);
   U9324 : NAND3_X1 port map( A1 => n13477, A2 => n13478, A3 => n13479, ZN => 
                           n7736);
   U9325 : NAND3_X1 port map( A1 => n13519, A2 => n13520, A3 => n13521, ZN => 
                           n7735);
   U9326 : NAND3_X1 port map( A1 => n13561, A2 => n13562, A3 => n13563, ZN => 
                           n7734);
   U9327 : NAND3_X1 port map( A1 => n13603, A2 => n13604, A3 => n13605, ZN => 
                           n7733);
   U9328 : NAND3_X1 port map( A1 => n13645, A2 => n13646, A3 => n13647, ZN => 
                           n7732);
   U9329 : NAND3_X1 port map( A1 => n13687, A2 => n13688, A3 => n13689, ZN => 
                           n7731);
   U9330 : NAND3_X1 port map( A1 => n13729, A2 => n13730, A3 => n13731, ZN => 
                           n7730);
   U9331 : NAND3_X1 port map( A1 => n13771, A2 => n13772, A3 => n13773, ZN => 
                           n7729);
   U9332 : NAND3_X1 port map( A1 => n13813, A2 => n13814, A3 => n13815, ZN => 
                           n7728);
   U9333 : NAND3_X1 port map( A1 => n13855, A2 => n13856, A3 => n13857, ZN => 
                           n7727);
   U9334 : NAND3_X1 port map( A1 => n13897, A2 => n13898, A3 => n13899, ZN => 
                           n7726);
   U9335 : XOR2_X1 port map( A => add_wr(3), B => add_rd2(3), Z => n13995);
   U9336 : NAND3_X1 port map( A1 => enable, A2 => n18044, A3 => rd2, ZN => 
                           n12527);
   U9337 : XOR2_X1 port map( A => n3043, B => n14011, Z => n14010);
   U9338 : NAND3_X1 port map( A1 => call, A2 => n14023, A3 => n14024, ZN => 
                           n13997);
   U9339 : NAND3_X1 port map( A1 => n14025, A2 => n14024, A3 => ret, ZN => 
                           n13998);
   U9340 : XOR2_X1 port map( A => swp_5_port, B => n3043, Z => n14023);
   U9341 : NAND3_X1 port map( A1 => n14129, A2 => r590_carry_5_port, A3 => 
                           n14147, ZN => n14101);
   U9342 : NAND3_X1 port map( A1 => r590_carry_5_port, A2 => n14133, A3 => 
                           n14147, ZN => n14142);
   U9343 : NAND3_X1 port map( A1 => N9926, A2 => N9924, A3 => N9922, ZN => 
                           n14183);
   U9344 : NAND3_X1 port map( A1 => r590_carry_5_port, A2 => n14133, A3 => 
                           n14178, ZN => n14185);
   U9345 : NAND3_X1 port map( A1 => N9924, A2 => n14173, A3 => N9926, ZN => 
                           n14207);
   U9346 : NAND3_X1 port map( A1 => n14178, A2 => r590_carry_5_port, A3 => 
                           n14129, ZN => n14181);
   U9347 : NAND3_X1 port map( A1 => n14193, A2 => call, A3 => n14179, ZN => 
                           n14211);
   U9348 : NAND3_X1 port map( A1 => n14196, A2 => n10189, A3 => n10187, ZN => 
                           n14116);
   U9349 : XOR2_X1 port map( A => n3043, B => n14820, Z => n14178);
   U9353 : XOR2_X1 port map( A => n7587, B => n14229, Z => n14263);
   add_148 : w_reg_file_M8_N8_F4_Nbit32_DW01_add_0 port map( A(5) => n4, A(4) 
                           => add_rd2(4), A(3) => add_rd2(3), A(2) => 
                           add_rd2(2), A(1) => add_rd2(1), A(0) => add_rd2(0), 
                           B(5) => N51637, B(4) => r590_carry_5_port, B(3) => 
                           N9910, B(2) => N9909, B(1) => N9908, B(0) => N9641, 
                           CI => n76, SUM(5) => N46303, SUM(4) => N46302, 
                           SUM(3) => N46301, SUM(2) => N46300, SUM(1) => N46299
                           , SUM(0) => N46298, CO => net226798);
   add_134 : w_reg_file_M8_N8_F4_Nbit32_DW01_add_1 port map( A(5) => n4, A(4) 
                           => add_rd1(4), A(3) => add_rd1(3), A(2) => 
                           add_rd1(2), A(1) => add_rd1(1), A(0) => add_rd1(0), 
                           B(5) => N51637, B(4) => r590_carry_5_port, B(3) => 
                           N9910, B(2) => N9909, B(1) => N9908, B(0) => N9641, 
                           CI => n77, SUM(5) => N45789, SUM(4) => N45788, 
                           SUM(3) => N45787, SUM(2) => N45786, SUM(1) => N45785
                           , SUM(0) => N45784, CO => net226797);
   add_101 : w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0 port map( A(5) => i_5_port, 
                           A(4) => i_4_port, A(3) => i_3_port, A(2) => i_2_port
                           , A(1) => i_1_port, A(0) => i_0_port, SUM(5) => 
                           N9926, SUM(4) => N9925, SUM(3) => N9924, SUM(2) => 
                           N9923, SUM(1) => N9922, SUM(0) => N9921);
   cwp_reg_4_inst : DFF_X1 port map( D => n10182, CK => clk, Q => 
                           r590_carry_5_port, QN => n14820);
   U6 : NOR2_X1 port map( A1 => n13979, A2 => N46298, ZN => n13932);
   U7 : NOR2_X1 port map( A1 => n12498, A2 => N45784, ZN => n12452);
   U8 : TINV_X1 port map( I => n7694, EN => n6613, ZN => to_mem(31));
   U9 : TINV_X1 port map( I => n7695, EN => n6620, ZN => to_mem(30));
   U10 : TINV_X1 port map( I => n7696, EN => n6621, ZN => to_mem(29));
   U11 : TINV_X1 port map( I => n7697, EN => n6624, ZN => to_mem(28));
   U12 : TINV_X1 port map( I => n7698, EN => n6630, ZN => to_mem(27));
   U13 : TINV_X1 port map( I => n7699, EN => n6632, ZN => to_mem(26));
   U14 : TINV_X1 port map( I => n7700, EN => n6634, ZN => to_mem(25));
   U15 : TINV_X1 port map( I => n7701, EN => n6641, ZN => to_mem(24));
   U16 : TINV_X1 port map( I => n7702, EN => n6642, ZN => to_mem(23));
   U17 : TINV_X1 port map( I => n7703, EN => n6646, ZN => to_mem(22));
   U18 : TINV_X1 port map( I => n7704, EN => n6647, ZN => to_mem(21));
   U19 : TINV_X1 port map( I => n7705, EN => n6648, ZN => to_mem(20));
   U20 : TINV_X1 port map( I => n7706, EN => n6649, ZN => to_mem(19));
   U21 : TINV_X1 port map( I => n7707, EN => n6650, ZN => to_mem(18));
   U22 : TINV_X1 port map( I => n7708, EN => n6651, ZN => to_mem(17));
   U23 : TINV_X1 port map( I => n7709, EN => n6652, ZN => to_mem(16));
   U24 : TINV_X1 port map( I => n7710, EN => n6653, ZN => to_mem(15));
   U25 : TINV_X1 port map( I => n7711, EN => n6654, ZN => to_mem(14));
   U26 : TINV_X1 port map( I => n7712, EN => n6655, ZN => to_mem(13));
   U27 : TINV_X1 port map( I => n7713, EN => n6656, ZN => to_mem(12));
   U28 : TINV_X1 port map( I => n7714, EN => n6657, ZN => to_mem(11));
   U29 : TINV_X1 port map( I => n7715, EN => n6658, ZN => to_mem(10));
   U30 : TINV_X1 port map( I => n7716, EN => n6659, ZN => to_mem(9));
   U31 : TINV_X1 port map( I => n7717, EN => n6660, ZN => to_mem(8));
   U32 : TINV_X1 port map( I => n7718, EN => n6671, ZN => to_mem(7));
   U33 : TINV_X1 port map( I => n7719, EN => n6674, ZN => to_mem(6));
   U34 : TINV_X1 port map( I => n7720, EN => n6676, ZN => to_mem(5));
   U35 : TINV_X1 port map( I => n7721, EN => n6683, ZN => to_mem(4));
   U36 : TINV_X1 port map( I => n7722, EN => n6684, ZN => to_mem(3));
   U37 : TINV_X1 port map( I => n7723, EN => n6687, ZN => to_mem(2));
   U38 : TINV_X1 port map( I => n7724, EN => n6693, ZN => to_mem(1));
   U39 : TINV_X1 port map( I => n7725, EN => n6695, ZN => to_mem(0));
   U40 : NOR2_X1 port map( A1 => n13979, A2 => n13978, ZN => n13918);
   U41 : NOR2_X1 port map( A1 => n12498, A2 => n12497, ZN => n12437);
   U42 : NOR2_X1 port map( A1 => N45784, A2 => N45785, ZN => n12451);
   U43 : NOR2_X1 port map( A1 => N46298, A2 => N46299, ZN => n13927);
   U44 : NOR2_X1 port map( A1 => n13978, A2 => N46299, ZN => n13935);
   U45 : NOR2_X1 port map( A1 => n12497, A2 => N45785, ZN => n12454);
   U46 : INV_X1 port map( A => n17984, ZN => n17965);
   U47 : INV_X1 port map( A => n17324, ZN => n17321);
   U48 : INV_X1 port map( A => n17337, ZN => n17334);
   U49 : INV_X1 port map( A => n17350, ZN => n17347);
   U50 : INV_X1 port map( A => n17363, ZN => n17360);
   U51 : INV_X1 port map( A => n17402, ZN => n17399);
   U52 : INV_X1 port map( A => n17428, ZN => n17425);
   U53 : INV_X1 port map( A => n17441, ZN => n17438);
   U54 : INV_X1 port map( A => n17454, ZN => n17450);
   U55 : INV_X1 port map( A => n17467, ZN => n17464);
   U56 : INV_X1 port map( A => n17480, ZN => n17477);
   U57 : INV_X1 port map( A => n17493, ZN => n17490);
   U58 : INV_X1 port map( A => n17506, ZN => n17503);
   U59 : INV_X1 port map( A => n17984, ZN => n17966);
   U60 : INV_X1 port map( A => n17323, ZN => n17320);
   U61 : INV_X1 port map( A => n17427, ZN => n17424);
   U62 : INV_X1 port map( A => n17336, ZN => n17333);
   U63 : INV_X1 port map( A => n17349, ZN => n17346);
   U64 : INV_X1 port map( A => n17440, ZN => n17437);
   U65 : INV_X1 port map( A => n17479, ZN => n17476);
   U66 : INV_X1 port map( A => n17999, ZN => n17989);
   U67 : INV_X1 port map( A => n17362, ZN => n17359);
   U68 : INV_X1 port map( A => n17401, ZN => n17398);
   U69 : INV_X1 port map( A => n17466, ZN => n17463);
   U70 : INV_X1 port map( A => n17492, ZN => n17489);
   U71 : INV_X1 port map( A => n17505, ZN => n17502);
   U72 : INV_X1 port map( A => n17525, ZN => n17522);
   U73 : INV_X1 port map( A => n17999, ZN => n17990);
   U74 : INV_X1 port map( A => n17414, ZN => n17411);
   U75 : INV_X1 port map( A => n17415, ZN => n17412);
   U76 : INV_X1 port map( A => n17524, ZN => n17521);
   U77 : INV_X1 port map( A => n17018, ZN => n17009);
   U78 : INV_X1 port map( A => n17211, ZN => n17202);
   U79 : INV_X1 port map( A => n17855, ZN => n17836);
   U80 : INV_X1 port map( A => n17877, ZN => n17858);
   U81 : INV_X1 port map( A => n17899, ZN => n17880);
   U82 : INV_X1 port map( A => n17921, ZN => n17902);
   U83 : INV_X1 port map( A => n17942, ZN => n17923);
   U84 : INV_X1 port map( A => n17963, ZN => n17944);
   U85 : INV_X1 port map( A => n18007, ZN => n18004);
   U86 : INV_X1 port map( A => n18020, ZN => n18017);
   U87 : INV_X1 port map( A => n16904, ZN => n16901);
   U88 : INV_X1 port map( A => n16938, ZN => n16935);
   U89 : INV_X1 port map( A => n16993, ZN => n16990);
   U90 : INV_X1 port map( A => n17027, ZN => n17024);
   U91 : INV_X1 port map( A => n17040, ZN => n17037);
   U92 : INV_X1 port map( A => n17053, ZN => n17050);
   U93 : INV_X1 port map( A => n17066, ZN => n17063);
   U94 : INV_X1 port map( A => n17079, ZN => n17076);
   U95 : INV_X1 port map( A => n17092, ZN => n17089);
   U96 : INV_X1 port map( A => n17105, ZN => n17102);
   U97 : INV_X1 port map( A => n17131, ZN => n17128);
   U98 : INV_X1 port map( A => n17154, ZN => n17151);
   U99 : INV_X1 port map( A => n17220, ZN => n17217);
   U100 : INV_X1 port map( A => n17233, ZN => n17230);
   U101 : INV_X1 port map( A => n17246, ZN => n17243);
   U102 : INV_X1 port map( A => n17259, ZN => n17256);
   U103 : INV_X1 port map( A => n17272, ZN => n17269);
   U104 : INV_X1 port map( A => n17285, ZN => n17282);
   U105 : INV_X1 port map( A => n17298, ZN => n17295);
   U106 : INV_X1 port map( A => n17376, ZN => n17373);
   U107 : INV_X1 port map( A => n17389, ZN => n17386);
   U108 : INV_X1 port map( A => n17855, ZN => n17837);
   U109 : INV_X1 port map( A => n17877, ZN => n17859);
   U110 : INV_X1 port map( A => n17899, ZN => n17881);
   U111 : INV_X1 port map( A => n17921, ZN => n17903);
   U112 : INV_X1 port map( A => n17942, ZN => n17924);
   U113 : INV_X1 port map( A => n17963, ZN => n17945);
   U114 : INV_X1 port map( A => n17219, ZN => n17216);
   U115 : INV_X1 port map( A => n16937, ZN => n16934);
   U116 : INV_X1 port map( A => n17026, ZN => n17023);
   U117 : INV_X1 port map( A => n17130, ZN => n17127);
   U118 : INV_X1 port map( A => n18006, ZN => n18003);
   U119 : INV_X1 port map( A => n17153, ZN => n17150);
   U120 : INV_X1 port map( A => n16876, ZN => n16866);
   U121 : INV_X1 port map( A => n17271, ZN => n17268);
   U122 : INV_X1 port map( A => n17039, ZN => n17036);
   U123 : INV_X1 port map( A => n17052, ZN => n17049);
   U124 : INV_X1 port map( A => n17078, ZN => n17075);
   U125 : INV_X1 port map( A => n17232, ZN => n17229);
   U126 : INV_X1 port map( A => n17245, ZN => n17242);
   U127 : INV_X1 port map( A => n17375, ZN => n17372);
   U128 : INV_X1 port map( A => n18019, ZN => n18016);
   U129 : INV_X1 port map( A => n16903, ZN => n16900);
   U130 : INV_X1 port map( A => n16992, ZN => n16989);
   U131 : INV_X1 port map( A => n17065, ZN => n17062);
   U132 : INV_X1 port map( A => n17091, ZN => n17088);
   U133 : INV_X1 port map( A => n17104, ZN => n17101);
   U134 : INV_X1 port map( A => n17258, ZN => n17255);
   U135 : INV_X1 port map( A => n17284, ZN => n17281);
   U136 : INV_X1 port map( A => n17297, ZN => n17294);
   U137 : INV_X1 port map( A => n17388, ZN => n17385);
   U138 : INV_X1 port map( A => n17117, ZN => n17114);
   U139 : INV_X1 port map( A => n17310, ZN => n17307);
   U140 : INV_X1 port map( A => n17118, ZN => n17115);
   U141 : INV_X1 port map( A => n17311, ZN => n17308);
   U142 : INV_X1 port map( A => n16929, ZN => n16920);
   U143 : INV_X1 port map( A => n16876, ZN => n16867);
   U144 : INV_X1 port map( A => n16954, ZN => n16945);
   U145 : INV_X1 port map( A => n17180, ZN => n17171);
   U146 : BUF_X1 port map( A => n17518, Z => n17525);
   U147 : BUF_X1 port map( A => n17317, Z => n17323);
   U148 : BUF_X1 port map( A => n17330, Z => n17336);
   U149 : BUF_X1 port map( A => n17343, Z => n17349);
   U150 : BUF_X1 port map( A => n17356, Z => n17362);
   U151 : BUF_X1 port map( A => n17421, Z => n17427);
   U152 : BUF_X1 port map( A => n17434, Z => n17440);
   U153 : BUF_X1 port map( A => n17447, Z => n17453);
   U154 : BUF_X1 port map( A => n17460, Z => n17466);
   U155 : BUF_X1 port map( A => n17473, Z => n17479);
   U156 : BUF_X1 port map( A => n17486, Z => n17492);
   U157 : BUF_X1 port map( A => n17499, Z => n17505);
   U158 : BUF_X1 port map( A => n17395, Z => n17401);
   U159 : BUF_X1 port map( A => n17408, Z => n17414);
   U160 : BUF_X1 port map( A => n17317, Z => n17324);
   U161 : BUF_X1 port map( A => n17330, Z => n17337);
   U162 : BUF_X1 port map( A => n17343, Z => n17350);
   U163 : BUF_X1 port map( A => n17356, Z => n17363);
   U164 : BUF_X1 port map( A => n17421, Z => n17428);
   U165 : BUF_X1 port map( A => n17434, Z => n17441);
   U166 : BUF_X1 port map( A => n17447, Z => n17454);
   U167 : BUF_X1 port map( A => n17460, Z => n17467);
   U168 : BUF_X1 port map( A => n17473, Z => n17480);
   U169 : BUF_X1 port map( A => n17486, Z => n17493);
   U170 : BUF_X1 port map( A => n17499, Z => n17506);
   U171 : BUF_X1 port map( A => n17518, Z => n17524);
   U172 : BUF_X1 port map( A => n17395, Z => n17402);
   U173 : BUF_X1 port map( A => n17408, Z => n17415);
   U174 : BUF_X1 port map( A => n17201, Z => n17200);
   U175 : BUF_X1 port map( A => n17008, Z => n17007);
   U176 : BUF_X1 port map( A => n17318, Z => n17325);
   U177 : BUF_X1 port map( A => n17331, Z => n17338);
   U178 : BUF_X1 port map( A => n17344, Z => n17351);
   U179 : BUF_X1 port map( A => n17357, Z => n17364);
   U180 : BUF_X1 port map( A => n17422, Z => n17429);
   U181 : BUF_X1 port map( A => n17435, Z => n17442);
   U182 : BUF_X1 port map( A => n17448, Z => n17455);
   U183 : BUF_X1 port map( A => n17461, Z => n17468);
   U184 : BUF_X1 port map( A => n17474, Z => n17481);
   U185 : BUF_X1 port map( A => n17487, Z => n17494);
   U186 : BUF_X1 port map( A => n17500, Z => n17507);
   U187 : BUF_X1 port map( A => n17519, Z => n17526);
   U188 : BUF_X1 port map( A => n17396, Z => n17403);
   U189 : BUF_X1 port map( A => n17409, Z => n17416);
   U190 : BUF_X1 port map( A => n17019, Z => n17018);
   U191 : BUF_X1 port map( A => n17212, Z => n17211);
   U192 : BUF_X1 port map( A => n17317, Z => n17322);
   U193 : BUF_X1 port map( A => n17330, Z => n17335);
   U194 : BUF_X1 port map( A => n17343, Z => n17348);
   U195 : BUF_X1 port map( A => n17356, Z => n17361);
   U196 : BUF_X1 port map( A => n17395, Z => n17400);
   U197 : BUF_X1 port map( A => n17408, Z => n17413);
   U198 : BUF_X1 port map( A => n17008, Z => n17000);
   U199 : BUF_X1 port map( A => n17201, Z => n17193);
   U200 : BUF_X1 port map( A => n17421, Z => n17426);
   U201 : BUF_X1 port map( A => n17434, Z => n17439);
   U202 : BUF_X1 port map( A => n17447, Z => n17452);
   U203 : BUF_X1 port map( A => n17460, Z => n17465);
   U204 : BUF_X1 port map( A => n17473, Z => n17478);
   U205 : BUF_X1 port map( A => n17486, Z => n17491);
   U206 : BUF_X1 port map( A => n17499, Z => n17504);
   U207 : BUF_X1 port map( A => n17518, Z => n17523);
   U208 : BUF_X1 port map( A => n17015, Z => n17016);
   U209 : BUF_X1 port map( A => n17208, Z => n17209);
   U210 : BUF_X1 port map( A => n17000, Z => n17006);
   U211 : BUF_X1 port map( A => n17193, Z => n17199);
   U212 : BUF_X1 port map( A => n17019, Z => n17015);
   U213 : BUF_X1 port map( A => n17212, Z => n17208);
   U214 : BUF_X1 port map( A => n17002, Z => n17005);
   U215 : BUF_X1 port map( A => n17195, Z => n17198);
   U216 : BUF_X1 port map( A => n17019, Z => n17013);
   U217 : BUF_X1 port map( A => n17212, Z => n17206);
   U218 : BUF_X1 port map( A => n17001, Z => n17003);
   U219 : BUF_X1 port map( A => n17194, Z => n17196);
   U220 : BUF_X1 port map( A => n17019, Z => n17012);
   U221 : BUF_X1 port map( A => n17212, Z => n17205);
   U222 : BUF_X1 port map( A => n17008, Z => n17002);
   U223 : BUF_X1 port map( A => n17201, Z => n17195);
   U224 : BUF_X1 port map( A => n17019, Z => n17011);
   U225 : BUF_X1 port map( A => n17212, Z => n17204);
   U226 : BUF_X1 port map( A => n17008, Z => n17001);
   U227 : BUF_X1 port map( A => n17201, Z => n17194);
   U228 : BUF_X1 port map( A => n17019, Z => n17010);
   U229 : BUF_X1 port map( A => n17212, Z => n17203);
   U230 : BUF_X1 port map( A => n17002, Z => n17004);
   U231 : BUF_X1 port map( A => n17019, Z => n17014);
   U232 : BUF_X1 port map( A => n17195, Z => n17197);
   U233 : BUF_X1 port map( A => n17212, Z => n17207);
   U234 : BUF_X1 port map( A => n17986, Z => n17991);
   U235 : BUF_X1 port map( A => n17986, Z => n17992);
   U236 : BUF_X1 port map( A => n17422, Z => n17431);
   U237 : BUF_X1 port map( A => n17435, Z => n17444);
   U238 : BUF_X1 port map( A => n17448, Z => n17457);
   U239 : BUF_X1 port map( A => n17461, Z => n17470);
   U240 : BUF_X1 port map( A => n17474, Z => n17483);
   U241 : BUF_X1 port map( A => n17487, Z => n17496);
   U242 : BUF_X1 port map( A => n17500, Z => n17509);
   U243 : BUF_X1 port map( A => n17519, Z => n17528);
   U244 : BUF_X1 port map( A => n17318, Z => n17327);
   U245 : BUF_X1 port map( A => n17331, Z => n17340);
   U246 : BUF_X1 port map( A => n17344, Z => n17353);
   U247 : BUF_X1 port map( A => n17357, Z => n17366);
   U248 : BUF_X1 port map( A => n17318, Z => n17326);
   U249 : BUF_X1 port map( A => n17331, Z => n17339);
   U250 : BUF_X1 port map( A => n17344, Z => n17352);
   U251 : BUF_X1 port map( A => n17357, Z => n17365);
   U252 : BUF_X1 port map( A => n17422, Z => n17430);
   U253 : BUF_X1 port map( A => n17435, Z => n17443);
   U254 : BUF_X1 port map( A => n17448, Z => n17456);
   U255 : BUF_X1 port map( A => n17461, Z => n17469);
   U256 : BUF_X1 port map( A => n17474, Z => n17482);
   U257 : BUF_X1 port map( A => n17487, Z => n17495);
   U258 : BUF_X1 port map( A => n17500, Z => n17508);
   U259 : BUF_X1 port map( A => n17519, Z => n17527);
   U260 : BUF_X1 port map( A => n17988, Z => n17998);
   U261 : BUF_X1 port map( A => n17988, Z => n17997);
   U262 : BUF_X1 port map( A => n17396, Z => n17405);
   U263 : BUF_X1 port map( A => n17409, Z => n17418);
   U264 : BUF_X1 port map( A => n17987, Z => n17996);
   U265 : BUF_X1 port map( A => n17987, Z => n17994);
   U266 : BUF_X1 port map( A => n17987, Z => n17995);
   U267 : BUF_X1 port map( A => n17986, Z => n17993);
   U268 : BUF_X1 port map( A => n17396, Z => n17404);
   U269 : BUF_X1 port map( A => n17409, Z => n17417);
   U270 : BUF_X1 port map( A => n17423, Z => n17432);
   U271 : BUF_X1 port map( A => n17436, Z => n17445);
   U272 : BUF_X1 port map( A => n17449, Z => n17458);
   U273 : BUF_X1 port map( A => n17462, Z => n17471);
   U274 : BUF_X1 port map( A => n17475, Z => n17484);
   U275 : BUF_X1 port map( A => n17488, Z => n17497);
   U276 : BUF_X1 port map( A => n17501, Z => n17510);
   U277 : BUF_X1 port map( A => n17520, Z => n17529);
   U278 : BUF_X1 port map( A => n17319, Z => n17328);
   U279 : BUF_X1 port map( A => n17332, Z => n17341);
   U280 : BUF_X1 port map( A => n17345, Z => n17354);
   U281 : BUF_X1 port map( A => n17358, Z => n17367);
   U282 : BUF_X1 port map( A => n17319, Z => n17329);
   U283 : BUF_X1 port map( A => n17332, Z => n17342);
   U284 : BUF_X1 port map( A => n17345, Z => n17355);
   U285 : BUF_X1 port map( A => n17358, Z => n17368);
   U286 : BUF_X1 port map( A => n17423, Z => n17433);
   U287 : BUF_X1 port map( A => n17436, Z => n17446);
   U288 : BUF_X1 port map( A => n17449, Z => n17459);
   U289 : BUF_X1 port map( A => n17462, Z => n17472);
   U290 : BUF_X1 port map( A => n17475, Z => n17485);
   U291 : BUF_X1 port map( A => n17488, Z => n17498);
   U292 : BUF_X1 port map( A => n17501, Z => n17511);
   U293 : BUF_X1 port map( A => n17520, Z => n17530);
   U294 : BUF_X1 port map( A => n17397, Z => n17406);
   U295 : BUF_X1 port map( A => n17410, Z => n17419);
   U296 : BUF_X1 port map( A => n17397, Z => n17407);
   U297 : BUF_X1 port map( A => n17410, Z => n17420);
   U298 : BUF_X1 port map( A => n17012, Z => n17017);
   U299 : BUF_X1 port map( A => n17205, Z => n17210);
   U300 : BUF_X1 port map( A => n17988, Z => n17999);
   U301 : INV_X1 port map( A => n18052, ZN => n18039);
   U302 : INV_X1 port map( A => n18051, ZN => n18035);
   U303 : INV_X1 port map( A => n18051, ZN => n18036);
   U304 : INV_X1 port map( A => n18052, ZN => n18041);
   U305 : INV_X1 port map( A => n18052, ZN => n18040);
   U306 : INV_X1 port map( A => n18052, ZN => n18038);
   U307 : INV_X1 port map( A => n16695, ZN => n16691);
   U308 : INV_X1 port map( A => n17580, ZN => n17576);
   U309 : INV_X1 port map( A => n17834, ZN => n17824);
   U310 : INV_X1 port map( A => n17558, ZN => n17548);
   U311 : INV_X1 port map( A => n17544, ZN => n17534);
   U312 : INV_X1 port map( A => n17572, ZN => n17562);
   U313 : INV_X1 port map( A => n17599, ZN => n17589);
   U314 : INV_X1 port map( A => n17613, ZN => n17603);
   U315 : INV_X1 port map( A => n17627, ZN => n17617);
   U316 : INV_X1 port map( A => n17627, ZN => n17618);
   U317 : INV_X1 port map( A => n18053, ZN => n18044);
   U318 : BUF_X1 port map( A => n12578, Z => n16322);
   U319 : BUF_X1 port map( A => n12543, Z => n16394);
   U320 : BUF_X1 port map( A => n12619, Z => n16247);
   U321 : BUF_X1 port map( A => n12578, Z => n16323);
   U322 : BUF_X1 port map( A => n12543, Z => n16395);
   U323 : BUF_X1 port map( A => n12619, Z => n16248);
   U324 : BUF_X1 port map( A => n10590, Z => n16574);
   U325 : BUF_X1 port map( A => n10536, Z => n16658);
   U326 : BUF_X1 port map( A => n10642, Z => n16499);
   U327 : BUF_X1 port map( A => n10590, Z => n16575);
   U328 : BUF_X1 port map( A => n10536, Z => n16659);
   U329 : BUF_X1 port map( A => n10642, Z => n16500);
   U330 : INV_X1 port map( A => n18053, ZN => n18043);
   U331 : INV_X1 port map( A => n18053, ZN => n18042);
   U332 : BUF_X1 port map( A => n12553, Z => n16373);
   U333 : BUF_X1 port map( A => n12553, Z => n16374);
   U334 : BUF_X1 port map( A => n10556, Z => n16625);
   U335 : BUF_X1 port map( A => n10556, Z => n16626);
   U336 : INV_X1 port map( A => n17544, ZN => n17535);
   U337 : INV_X1 port map( A => n17558, ZN => n17549);
   U338 : INV_X1 port map( A => n17572, ZN => n17563);
   U339 : INV_X1 port map( A => n17599, ZN => n17590);
   U340 : INV_X1 port map( A => n17613, ZN => n17604);
   U341 : BUF_X1 port map( A => n12566, Z => n16352);
   U342 : BUF_X1 port map( A => n12566, Z => n16353);
   U343 : BUF_X1 port map( A => n10573, Z => n16604);
   U344 : BUF_X1 port map( A => n10573, Z => n16605);
   U345 : BUF_X1 port map( A => n12616, Z => n16256);
   U346 : BUF_X1 port map( A => n12616, Z => n16257);
   U347 : BUF_X1 port map( A => n10637, Z => n16508);
   U348 : BUF_X1 port map( A => n10637, Z => n16509);
   U349 : BUF_X1 port map( A => n12576, Z => n16328);
   U350 : BUF_X1 port map( A => n12541, Z => n16400);
   U351 : BUF_X1 port map( A => n12546, Z => n16388);
   U352 : BUF_X1 port map( A => n12595, Z => n16292);
   U353 : BUF_X1 port map( A => n12576, Z => n16329);
   U354 : BUF_X1 port map( A => n12541, Z => n16401);
   U355 : BUF_X1 port map( A => n12546, Z => n16389);
   U356 : BUF_X1 port map( A => n12595, Z => n16293);
   U357 : BUF_X1 port map( A => n10594, Z => n16568);
   U358 : BUF_X1 port map( A => n10540, Z => n16652);
   U359 : BUF_X1 port map( A => n10547, Z => n16640);
   U360 : BUF_X1 port map( A => n10612, Z => n16544);
   U361 : BUF_X1 port map( A => n10594, Z => n16569);
   U362 : BUF_X1 port map( A => n10540, Z => n16653);
   U363 : BUF_X1 port map( A => n10547, Z => n16641);
   U364 : BUF_X1 port map( A => n10612, Z => n16545);
   U365 : BUF_X1 port map( A => n4248, Z => n17629);
   U366 : BUF_X1 port map( A => n4112, Z => n17809);
   U367 : BUF_X1 port map( A => n4121, Z => n17797);
   U368 : BUF_X1 port map( A => n4128, Z => n17785);
   U369 : BUF_X1 port map( A => n4248, Z => n17628);
   U370 : BUF_X1 port map( A => n4112, Z => n17808);
   U371 : BUF_X1 port map( A => n4121, Z => n17796);
   U372 : BUF_X1 port map( A => n4128, Z => n17784);
   U373 : BUF_X1 port map( A => n12578, Z => n16324);
   U374 : BUF_X1 port map( A => n12543, Z => n16396);
   U375 : BUF_X1 port map( A => n12619, Z => n16249);
   U376 : BUF_X1 port map( A => n10590, Z => n16576);
   U377 : BUF_X1 port map( A => n10536, Z => n16660);
   U378 : BUF_X1 port map( A => n10642, Z => n16501);
   U379 : BUF_X1 port map( A => n12561, Z => n16364);
   U380 : BUF_X1 port map( A => n12537, Z => n16409);
   U381 : BUF_X1 port map( A => n12547, Z => n16385);
   U382 : BUF_X1 port map( A => n12586, Z => n16313);
   U383 : BUF_X1 port map( A => n12628, Z => n16226);
   U384 : BUF_X1 port map( A => n12561, Z => n16365);
   U385 : BUF_X1 port map( A => n12537, Z => n16410);
   U386 : BUF_X1 port map( A => n12547, Z => n16386);
   U387 : BUF_X1 port map( A => n12586, Z => n16314);
   U388 : BUF_X1 port map( A => n12628, Z => n16227);
   U389 : BUF_X1 port map( A => n10566, Z => n16616);
   U390 : BUF_X1 port map( A => n10535, Z => n16661);
   U391 : BUF_X1 port map( A => n10549, Z => n16637);
   U392 : BUF_X1 port map( A => n10600, Z => n16565);
   U393 : BUF_X1 port map( A => n10655, Z => n16478);
   U394 : BUF_X1 port map( A => n10566, Z => n16617);
   U395 : BUF_X1 port map( A => n10535, Z => n16662);
   U396 : BUF_X1 port map( A => n10549, Z => n16638);
   U397 : BUF_X1 port map( A => n10600, Z => n16566);
   U398 : BUF_X1 port map( A => n10655, Z => n16479);
   U399 : BUF_X1 port map( A => n12540, Z => n16403);
   U400 : BUF_X1 port map( A => n12540, Z => n16404);
   U401 : BUF_X1 port map( A => n10538, Z => n16655);
   U402 : BUF_X1 port map( A => n10538, Z => n16656);
   U403 : BUF_X1 port map( A => n4110, Z => n17812);
   U404 : BUF_X1 port map( A => n4110, Z => n17811);
   U405 : BUF_X1 port map( A => n12553, Z => n16375);
   U406 : BUF_X1 port map( A => n10556, Z => n16627);
   U407 : BUF_X1 port map( A => n12566, Z => n16354);
   U408 : BUF_X1 port map( A => n10573, Z => n16606);
   U409 : BUF_X1 port map( A => n12616, Z => n16258);
   U410 : BUF_X1 port map( A => n10637, Z => n16510);
   U411 : BUF_X1 port map( A => n12576, Z => n16330);
   U412 : BUF_X1 port map( A => n12541, Z => n16402);
   U413 : BUF_X1 port map( A => n12546, Z => n16390);
   U414 : BUF_X1 port map( A => n12595, Z => n16294);
   U415 : BUF_X1 port map( A => n10594, Z => n16570);
   U416 : BUF_X1 port map( A => n10540, Z => n16654);
   U417 : BUF_X1 port map( A => n10547, Z => n16642);
   U418 : BUF_X1 port map( A => n10612, Z => n16546);
   U419 : BUF_X1 port map( A => n4248, Z => n17630);
   U420 : BUF_X1 port map( A => n4112, Z => n17810);
   U421 : BUF_X1 port map( A => n4121, Z => n17798);
   U422 : BUF_X1 port map( A => n4128, Z => n17786);
   U423 : BUF_X1 port map( A => n12561, Z => n16366);
   U424 : BUF_X1 port map( A => n12537, Z => n16411);
   U425 : BUF_X1 port map( A => n12547, Z => n16387);
   U426 : BUF_X1 port map( A => n12586, Z => n16315);
   U427 : BUF_X1 port map( A => n12628, Z => n16228);
   U428 : BUF_X1 port map( A => n10566, Z => n16618);
   U429 : BUF_X1 port map( A => n10535, Z => n16663);
   U430 : BUF_X1 port map( A => n10549, Z => n16639);
   U431 : BUF_X1 port map( A => n10600, Z => n16567);
   U432 : BUF_X1 port map( A => n10655, Z => n16480);
   U433 : BUF_X1 port map( A => n12540, Z => n16405);
   U434 : BUF_X1 port map( A => n10538, Z => n16657);
   U435 : BUF_X1 port map( A => n4110, Z => n17813);
   U436 : BUF_X1 port map( A => n18000, Z => n18007);
   U437 : BUF_X1 port map( A => n18013, Z => n18020);
   U438 : BUF_X1 port map( A => n16897, Z => n16903);
   U439 : BUF_X1 port map( A => n16931, Z => n16937);
   U440 : BUF_X1 port map( A => n18000, Z => n18006);
   U441 : BUF_X1 port map( A => n16986, Z => n16992);
   U442 : BUF_X1 port map( A => n17020, Z => n17026);
   U443 : BUF_X1 port map( A => n17033, Z => n17039);
   U444 : BUF_X1 port map( A => n17046, Z => n17052);
   U445 : BUF_X1 port map( A => n17059, Z => n17065);
   U446 : BUF_X1 port map( A => n17072, Z => n17078);
   U447 : BUF_X1 port map( A => n17085, Z => n17091);
   U448 : BUF_X1 port map( A => n17098, Z => n17104);
   U449 : BUF_X1 port map( A => n17111, Z => n17117);
   U450 : BUF_X1 port map( A => n17124, Z => n17130);
   U451 : BUF_X1 port map( A => n17147, Z => n17153);
   U452 : BUF_X1 port map( A => n17213, Z => n17219);
   U453 : BUF_X1 port map( A => n17226, Z => n17232);
   U454 : BUF_X1 port map( A => n17239, Z => n17245);
   U455 : BUF_X1 port map( A => n17252, Z => n17258);
   U456 : BUF_X1 port map( A => n17265, Z => n17271);
   U457 : BUF_X1 port map( A => n17278, Z => n17284);
   U458 : BUF_X1 port map( A => n17291, Z => n17297);
   U459 : BUF_X1 port map( A => n17304, Z => n17310);
   U460 : BUF_X1 port map( A => n17369, Z => n17375);
   U461 : BUF_X1 port map( A => n17382, Z => n17388);
   U462 : BUF_X1 port map( A => n18013, Z => n18019);
   U463 : BUF_X1 port map( A => n16897, Z => n16904);
   U464 : BUF_X1 port map( A => n16931, Z => n16938);
   U465 : BUF_X1 port map( A => n16986, Z => n16993);
   U466 : BUF_X1 port map( A => n17020, Z => n17027);
   U467 : BUF_X1 port map( A => n17033, Z => n17040);
   U468 : BUF_X1 port map( A => n17046, Z => n17053);
   U469 : BUF_X1 port map( A => n17059, Z => n17066);
   U470 : BUF_X1 port map( A => n17072, Z => n17079);
   U471 : BUF_X1 port map( A => n17085, Z => n17092);
   U472 : BUF_X1 port map( A => n17098, Z => n17105);
   U473 : BUF_X1 port map( A => n17111, Z => n17118);
   U474 : BUF_X1 port map( A => n17124, Z => n17131);
   U475 : BUF_X1 port map( A => n17147, Z => n17154);
   U476 : BUF_X1 port map( A => n17213, Z => n17220);
   U477 : BUF_X1 port map( A => n17226, Z => n17233);
   U478 : BUF_X1 port map( A => n17239, Z => n17246);
   U479 : BUF_X1 port map( A => n17252, Z => n17259);
   U480 : BUF_X1 port map( A => n17265, Z => n17272);
   U481 : BUF_X1 port map( A => n17278, Z => n17285);
   U482 : BUF_X1 port map( A => n17291, Z => n17298);
   U483 : BUF_X1 port map( A => n17304, Z => n17311);
   U484 : BUF_X1 port map( A => n17369, Z => n17376);
   U485 : BUF_X1 port map( A => n17382, Z => n17389);
   U486 : BUF_X1 port map( A => n17181, Z => n17179);
   U487 : BUF_X1 port map( A => n17191, Z => n17190);
   U488 : BUF_X1 port map( A => n16886, Z => n16885);
   U489 : BUF_X1 port map( A => n16896, Z => n16895);
   U490 : BUF_X1 port map( A => n16919, Z => n16918);
   U491 : BUF_X1 port map( A => n16955, Z => n16953);
   U492 : BUF_X1 port map( A => n16965, Z => n16964);
   U493 : BUF_X1 port map( A => n16975, Z => n16974);
   U494 : BUF_X1 port map( A => n16985, Z => n16984);
   U495 : BUF_X1 port map( A => n17146, Z => n17145);
   U496 : BUF_X1 port map( A => n17169, Z => n17168);
   U497 : BUF_X1 port map( A => n18001, Z => n18008);
   U498 : BUF_X1 port map( A => n18014, Z => n18021);
   U499 : BUF_X1 port map( A => n16898, Z => n16905);
   U500 : BUF_X1 port map( A => n16932, Z => n16939);
   U501 : BUF_X1 port map( A => n17021, Z => n17028);
   U502 : BUF_X1 port map( A => n17034, Z => n17041);
   U503 : BUF_X1 port map( A => n17047, Z => n17054);
   U504 : BUF_X1 port map( A => n17060, Z => n17067);
   U505 : BUF_X1 port map( A => n17073, Z => n17080);
   U506 : BUF_X1 port map( A => n17086, Z => n17093);
   U507 : BUF_X1 port map( A => n17099, Z => n17106);
   U508 : BUF_X1 port map( A => n17112, Z => n17119);
   U509 : BUF_X1 port map( A => n17125, Z => n17132);
   U510 : BUF_X1 port map( A => n17148, Z => n17155);
   U511 : BUF_X1 port map( A => n17214, Z => n17221);
   U512 : BUF_X1 port map( A => n17227, Z => n17234);
   U513 : BUF_X1 port map( A => n17240, Z => n17247);
   U514 : BUF_X1 port map( A => n17253, Z => n17260);
   U515 : BUF_X1 port map( A => n17266, Z => n17273);
   U516 : BUF_X1 port map( A => n17279, Z => n17286);
   U517 : BUF_X1 port map( A => n17292, Z => n17299);
   U518 : BUF_X1 port map( A => n17305, Z => n17312);
   U519 : BUF_X1 port map( A => n16987, Z => n16994);
   U520 : BUF_X1 port map( A => n17370, Z => n17377);
   U521 : BUF_X1 port map( A => n17383, Z => n17390);
   U522 : BUF_X1 port map( A => n16930, Z => n16929);
   U523 : BUF_X1 port map( A => n16931, Z => n16936);
   U524 : BUF_X1 port map( A => n17124, Z => n17129);
   U525 : BUF_X1 port map( A => n18000, Z => n18005);
   U526 : BUF_X1 port map( A => n18013, Z => n18018);
   U527 : BUF_X1 port map( A => n17020, Z => n17025);
   U528 : BUF_X1 port map( A => n17033, Z => n17038);
   U529 : BUF_X1 port map( A => n17046, Z => n17051);
   U530 : BUF_X1 port map( A => n17059, Z => n17064);
   U531 : BUF_X1 port map( A => n17072, Z => n17077);
   U532 : BUF_X1 port map( A => n17085, Z => n17090);
   U533 : BUF_X1 port map( A => n17098, Z => n17103);
   U534 : BUF_X1 port map( A => n17111, Z => n17116);
   U535 : BUF_X1 port map( A => n17226, Z => n17231);
   U536 : BUF_X1 port map( A => n17239, Z => n17244);
   U537 : BUF_X1 port map( A => n17252, Z => n17257);
   U538 : BUF_X1 port map( A => n17278, Z => n17283);
   U539 : BUF_X1 port map( A => n17291, Z => n17296);
   U540 : BUF_X1 port map( A => n17304, Z => n17309);
   U541 : BUF_X1 port map( A => n17369, Z => n17374);
   U542 : BUF_X1 port map( A => n17382, Z => n17387);
   U543 : BUF_X1 port map( A => n16896, Z => n16888);
   U544 : BUF_X1 port map( A => n16955, Z => n16946);
   U545 : BUF_X1 port map( A => n16965, Z => n16957);
   U546 : BUF_X1 port map( A => n16985, Z => n16977);
   U547 : BUF_X1 port map( A => n17146, Z => n17138);
   U548 : BUF_X1 port map( A => n17181, Z => n17172);
   U549 : BUF_X1 port map( A => n16863, Z => n16868);
   U550 : BUF_X1 port map( A => n16886, Z => n16878);
   U551 : BUF_X1 port map( A => n16919, Z => n16911);
   U552 : BUF_X1 port map( A => n16975, Z => n16967);
   U553 : BUF_X1 port map( A => n17169, Z => n17161);
   U554 : BUF_X1 port map( A => n17191, Z => n17183);
   U555 : BUF_X1 port map( A => n16897, Z => n16902);
   U556 : BUF_X1 port map( A => n17147, Z => n17152);
   U557 : BUF_X1 port map( A => n16986, Z => n16991);
   U558 : BUF_X1 port map( A => n17213, Z => n17218);
   U559 : BUF_X1 port map( A => n17265, Z => n17270);
   U560 : BUF_X1 port map( A => n16926, Z => n16927);
   U561 : BUF_X1 port map( A => n16878, Z => n16884);
   U562 : BUF_X1 port map( A => n16911, Z => n16917);
   U563 : BUF_X1 port map( A => n16967, Z => n16973);
   U564 : BUF_X1 port map( A => n17161, Z => n17167);
   U565 : BUF_X1 port map( A => n17183, Z => n17189);
   U566 : BUF_X1 port map( A => n16888, Z => n16894);
   U567 : BUF_X1 port map( A => n16946, Z => n16952);
   U568 : BUF_X1 port map( A => n16957, Z => n16963);
   U569 : BUF_X1 port map( A => n16977, Z => n16983);
   U570 : BUF_X1 port map( A => n17138, Z => n17144);
   U571 : BUF_X1 port map( A => n17172, Z => n17178);
   U572 : BUF_X1 port map( A => n16930, Z => n16926);
   U573 : BUF_X1 port map( A => n16880, Z => n16883);
   U574 : BUF_X1 port map( A => n16913, Z => n16916);
   U575 : BUF_X1 port map( A => n16969, Z => n16972);
   U576 : BUF_X1 port map( A => n17163, Z => n17166);
   U577 : BUF_X1 port map( A => n17185, Z => n17188);
   U578 : BUF_X1 port map( A => n16890, Z => n16893);
   U579 : BUF_X1 port map( A => n16948, Z => n16951);
   U580 : BUF_X1 port map( A => n16959, Z => n16962);
   U581 : BUF_X1 port map( A => n16979, Z => n16982);
   U582 : BUF_X1 port map( A => n17140, Z => n17143);
   U583 : BUF_X1 port map( A => n17174, Z => n17177);
   U584 : BUF_X1 port map( A => n16930, Z => n16924);
   U585 : BUF_X1 port map( A => n16879, Z => n16881);
   U586 : BUF_X1 port map( A => n16912, Z => n16914);
   U587 : BUF_X1 port map( A => n16968, Z => n16970);
   U588 : BUF_X1 port map( A => n17162, Z => n17164);
   U589 : BUF_X1 port map( A => n17184, Z => n17186);
   U590 : BUF_X1 port map( A => n16889, Z => n16891);
   U591 : BUF_X1 port map( A => n16947, Z => n16949);
   U592 : BUF_X1 port map( A => n16958, Z => n16960);
   U593 : BUF_X1 port map( A => n16978, Z => n16980);
   U594 : BUF_X1 port map( A => n17139, Z => n17141);
   U595 : BUF_X1 port map( A => n17173, Z => n17175);
   U596 : BUF_X1 port map( A => n16930, Z => n16923);
   U597 : BUF_X1 port map( A => n16886, Z => n16880);
   U598 : BUF_X1 port map( A => n16919, Z => n16913);
   U599 : BUF_X1 port map( A => n16975, Z => n16969);
   U600 : BUF_X1 port map( A => n17169, Z => n17163);
   U601 : BUF_X1 port map( A => n17191, Z => n17185);
   U602 : BUF_X1 port map( A => n16896, Z => n16890);
   U603 : BUF_X1 port map( A => n16955, Z => n16948);
   U604 : BUF_X1 port map( A => n16965, Z => n16959);
   U605 : BUF_X1 port map( A => n16985, Z => n16979);
   U606 : BUF_X1 port map( A => n17146, Z => n17140);
   U607 : BUF_X1 port map( A => n17181, Z => n17174);
   U608 : BUF_X1 port map( A => n16930, Z => n16922);
   U609 : BUF_X1 port map( A => n16919, Z => n16912);
   U610 : BUF_X1 port map( A => n17191, Z => n17184);
   U611 : BUF_X1 port map( A => n16896, Z => n16889);
   U612 : BUF_X1 port map( A => n16955, Z => n16947);
   U613 : BUF_X1 port map( A => n16965, Z => n16958);
   U614 : BUF_X1 port map( A => n16985, Z => n16978);
   U615 : BUF_X1 port map( A => n17146, Z => n17139);
   U616 : BUF_X1 port map( A => n17181, Z => n17173);
   U617 : BUF_X1 port map( A => n16886, Z => n16879);
   U618 : BUF_X1 port map( A => n16975, Z => n16968);
   U619 : BUF_X1 port map( A => n17169, Z => n17162);
   U620 : BUF_X1 port map( A => n16930, Z => n16921);
   U621 : BUF_X1 port map( A => n16880, Z => n16882);
   U622 : BUF_X1 port map( A => n16890, Z => n16892);
   U623 : BUF_X1 port map( A => n16913, Z => n16915);
   U624 : BUF_X1 port map( A => n16930, Z => n16925);
   U625 : BUF_X1 port map( A => n16948, Z => n16950);
   U626 : BUF_X1 port map( A => n16959, Z => n16961);
   U627 : BUF_X1 port map( A => n16969, Z => n16971);
   U628 : BUF_X1 port map( A => n16979, Z => n16981);
   U629 : BUF_X1 port map( A => n17140, Z => n17142);
   U630 : BUF_X1 port map( A => n17163, Z => n17165);
   U631 : BUF_X1 port map( A => n17174, Z => n17176);
   U632 : BUF_X1 port map( A => n17185, Z => n17187);
   U633 : BUF_X1 port map( A => n16865, Z => n16874);
   U634 : BUF_X1 port map( A => n17021, Z => n17030);
   U635 : BUF_X1 port map( A => n17034, Z => n17043);
   U636 : BUF_X1 port map( A => n17047, Z => n17056);
   U637 : BUF_X1 port map( A => n17060, Z => n17069);
   U638 : BUF_X1 port map( A => n17073, Z => n17082);
   U639 : BUF_X1 port map( A => n17086, Z => n17095);
   U640 : BUF_X1 port map( A => n17099, Z => n17108);
   U641 : BUF_X1 port map( A => n17112, Z => n17121);
   U642 : BUF_X1 port map( A => n17214, Z => n17223);
   U643 : BUF_X1 port map( A => n17227, Z => n17236);
   U644 : BUF_X1 port map( A => n17240, Z => n17249);
   U645 : BUF_X1 port map( A => n17253, Z => n17262);
   U646 : BUF_X1 port map( A => n17266, Z => n17275);
   U647 : BUF_X1 port map( A => n17279, Z => n17288);
   U648 : BUF_X1 port map( A => n17292, Z => n17301);
   U649 : BUF_X1 port map( A => n17305, Z => n17314);
   U650 : BUF_X1 port map( A => n16864, Z => n16873);
   U651 : BUF_X1 port map( A => n16898, Z => n16907);
   U652 : BUF_X1 port map( A => n16932, Z => n16941);
   U653 : BUF_X1 port map( A => n17125, Z => n17134);
   U654 : BUF_X1 port map( A => n17148, Z => n17157);
   U655 : BUF_X1 port map( A => n18001, Z => n18010);
   U656 : BUF_X1 port map( A => n18014, Z => n18023);
   U657 : BUF_X1 port map( A => n16864, Z => n16871);
   U658 : BUF_X1 port map( A => n18001, Z => n18009);
   U659 : BUF_X1 port map( A => n18014, Z => n18022);
   U660 : BUF_X1 port map( A => n16863, Z => n16870);
   U661 : BUF_X1 port map( A => n16863, Z => n16869);
   U662 : BUF_X1 port map( A => n16864, Z => n16872);
   U663 : BUF_X1 port map( A => n16898, Z => n16906);
   U664 : BUF_X1 port map( A => n16932, Z => n16940);
   U665 : BUF_X1 port map( A => n17021, Z => n17029);
   U666 : BUF_X1 port map( A => n17034, Z => n17042);
   U667 : BUF_X1 port map( A => n17047, Z => n17055);
   U668 : BUF_X1 port map( A => n17060, Z => n17068);
   U669 : BUF_X1 port map( A => n17073, Z => n17081);
   U670 : BUF_X1 port map( A => n17086, Z => n17094);
   U671 : BUF_X1 port map( A => n17099, Z => n17107);
   U672 : BUF_X1 port map( A => n17112, Z => n17120);
   U673 : BUF_X1 port map( A => n17125, Z => n17133);
   U674 : BUF_X1 port map( A => n17148, Z => n17156);
   U675 : BUF_X1 port map( A => n17214, Z => n17222);
   U676 : BUF_X1 port map( A => n17227, Z => n17235);
   U677 : BUF_X1 port map( A => n17240, Z => n17248);
   U678 : BUF_X1 port map( A => n17253, Z => n17261);
   U679 : BUF_X1 port map( A => n17266, Z => n17274);
   U680 : BUF_X1 port map( A => n17279, Z => n17287);
   U681 : BUF_X1 port map( A => n17292, Z => n17300);
   U682 : BUF_X1 port map( A => n17305, Z => n17313);
   U683 : BUF_X1 port map( A => n16865, Z => n16875);
   U684 : BUF_X1 port map( A => n17370, Z => n17379);
   U685 : BUF_X1 port map( A => n17383, Z => n17392);
   U686 : BUF_X1 port map( A => n16987, Z => n16996);
   U687 : BUF_X1 port map( A => n16987, Z => n16995);
   U688 : BUF_X1 port map( A => n17370, Z => n17378);
   U689 : BUF_X1 port map( A => n17383, Z => n17391);
   U690 : BUF_X1 port map( A => n18002, Z => n18012);
   U691 : BUF_X1 port map( A => n18015, Z => n18025);
   U692 : BUF_X1 port map( A => n17022, Z => n17031);
   U693 : BUF_X1 port map( A => n17035, Z => n17044);
   U694 : BUF_X1 port map( A => n17048, Z => n17057);
   U695 : BUF_X1 port map( A => n17061, Z => n17070);
   U696 : BUF_X1 port map( A => n17074, Z => n17083);
   U697 : BUF_X1 port map( A => n17087, Z => n17096);
   U698 : BUF_X1 port map( A => n17100, Z => n17109);
   U699 : BUF_X1 port map( A => n17113, Z => n17122);
   U700 : BUF_X1 port map( A => n17215, Z => n17224);
   U701 : BUF_X1 port map( A => n17228, Z => n17237);
   U702 : BUF_X1 port map( A => n17241, Z => n17250);
   U703 : BUF_X1 port map( A => n17254, Z => n17263);
   U704 : BUF_X1 port map( A => n17267, Z => n17276);
   U705 : BUF_X1 port map( A => n17280, Z => n17289);
   U706 : BUF_X1 port map( A => n17293, Z => n17302);
   U707 : BUF_X1 port map( A => n17306, Z => n17315);
   U708 : BUF_X1 port map( A => n16899, Z => n16908);
   U709 : BUF_X1 port map( A => n16933, Z => n16942);
   U710 : BUF_X1 port map( A => n17126, Z => n17135);
   U711 : BUF_X1 port map( A => n17149, Z => n17158);
   U712 : BUF_X1 port map( A => n18002, Z => n18011);
   U713 : BUF_X1 port map( A => n16899, Z => n16909);
   U714 : BUF_X1 port map( A => n18015, Z => n18024);
   U715 : BUF_X1 port map( A => n16933, Z => n16943);
   U716 : BUF_X1 port map( A => n17022, Z => n17032);
   U717 : BUF_X1 port map( A => n17035, Z => n17045);
   U718 : BUF_X1 port map( A => n17048, Z => n17058);
   U719 : BUF_X1 port map( A => n17061, Z => n17071);
   U720 : BUF_X1 port map( A => n17074, Z => n17084);
   U721 : BUF_X1 port map( A => n17087, Z => n17097);
   U722 : BUF_X1 port map( A => n17100, Z => n17110);
   U723 : BUF_X1 port map( A => n17113, Z => n17123);
   U724 : BUF_X1 port map( A => n17126, Z => n17136);
   U725 : BUF_X1 port map( A => n17149, Z => n17159);
   U726 : BUF_X1 port map( A => n17215, Z => n17225);
   U727 : BUF_X1 port map( A => n17228, Z => n17238);
   U728 : BUF_X1 port map( A => n17241, Z => n17251);
   U729 : BUF_X1 port map( A => n17254, Z => n17264);
   U730 : BUF_X1 port map( A => n17267, Z => n17277);
   U731 : BUF_X1 port map( A => n17280, Z => n17290);
   U732 : BUF_X1 port map( A => n17293, Z => n17303);
   U733 : BUF_X1 port map( A => n17306, Z => n17316);
   U734 : BUF_X1 port map( A => n17371, Z => n17380);
   U735 : BUF_X1 port map( A => n17384, Z => n17393);
   U736 : BUF_X1 port map( A => n16988, Z => n16997);
   U737 : BUF_X1 port map( A => n16988, Z => n16998);
   U738 : BUF_X1 port map( A => n17371, Z => n17381);
   U739 : BUF_X1 port map( A => n17384, Z => n17394);
   U740 : BUF_X1 port map( A => n16923, Z => n16928);
   U741 : BUF_X1 port map( A => n16865, Z => n16876);
   U742 : BUF_X1 port map( A => n16955, Z => n16954);
   U743 : BUF_X1 port map( A => n17181, Z => n17180);
   U744 : BUF_X1 port map( A => n4329, Z => n17317);
   U745 : BUF_X1 port map( A => n4326, Z => n17330);
   U746 : BUF_X1 port map( A => n4323, Z => n17343);
   U747 : BUF_X1 port map( A => n4320, Z => n17356);
   U748 : BUF_X1 port map( A => n4301, Z => n17421);
   U749 : BUF_X1 port map( A => n4298, Z => n17434);
   U750 : BUF_X1 port map( A => n4291, Z => n17447);
   U751 : BUF_X1 port map( A => n4288, Z => n17460);
   U752 : BUF_X1 port map( A => n4285, Z => n17473);
   U753 : BUF_X1 port map( A => n4282, Z => n17486);
   U754 : BUF_X1 port map( A => n4279, Z => n17499);
   U755 : BUF_X1 port map( A => n4275, Z => n17518);
   U756 : BUF_X1 port map( A => n4329, Z => n17318);
   U757 : BUF_X1 port map( A => n4326, Z => n17331);
   U758 : BUF_X1 port map( A => n4323, Z => n17344);
   U759 : BUF_X1 port map( A => n4320, Z => n17357);
   U760 : BUF_X1 port map( A => n4301, Z => n17422);
   U761 : BUF_X1 port map( A => n4298, Z => n17435);
   U762 : BUF_X1 port map( A => n4291, Z => n17448);
   U763 : BUF_X1 port map( A => n4288, Z => n17461);
   U764 : BUF_X1 port map( A => n4285, Z => n17474);
   U765 : BUF_X1 port map( A => n4282, Z => n17487);
   U766 : BUF_X1 port map( A => n4279, Z => n17500);
   U767 : BUF_X1 port map( A => n4275, Z => n17519);
   U768 : BUF_X1 port map( A => n4067, Z => n17988);
   U769 : BUF_X1 port map( A => n4067, Z => n17987);
   U770 : BUF_X1 port map( A => n4067, Z => n17986);
   U771 : BUF_X1 port map( A => n4309, Z => n17395);
   U772 : BUF_X1 port map( A => n4306, Z => n17408);
   U773 : BUF_X1 port map( A => n4309, Z => n17396);
   U774 : BUF_X1 port map( A => n4306, Z => n17409);
   U775 : BUF_X1 port map( A => n4329, Z => n17319);
   U776 : BUF_X1 port map( A => n4326, Z => n17332);
   U777 : BUF_X1 port map( A => n4323, Z => n17345);
   U778 : BUF_X1 port map( A => n4320, Z => n17358);
   U779 : BUF_X1 port map( A => n4301, Z => n17423);
   U780 : BUF_X1 port map( A => n4298, Z => n17436);
   U781 : BUF_X1 port map( A => n4291, Z => n17449);
   U782 : BUF_X1 port map( A => n4288, Z => n17462);
   U783 : BUF_X1 port map( A => n4285, Z => n17475);
   U784 : BUF_X1 port map( A => n4282, Z => n17488);
   U785 : BUF_X1 port map( A => n4279, Z => n17501);
   U786 : BUF_X1 port map( A => n4275, Z => n17520);
   U787 : BUF_X1 port map( A => n4309, Z => n17397);
   U788 : BUF_X1 port map( A => n4306, Z => n17410);
   U789 : INV_X1 port map( A => n16999, ZN => n17008);
   U790 : INV_X1 port map( A => n4420, ZN => n17019);
   U791 : INV_X1 port map( A => n17192, ZN => n17201);
   U792 : INV_X1 port map( A => n4362, ZN => n17212);
   U793 : INV_X1 port map( A => n18051, ZN => n18034);
   U794 : INV_X1 port map( A => n18051, ZN => n18037);
   U795 : INV_X1 port map( A => n17834, ZN => n17823);
   U796 : OAI21_X1 port map( B1 => n14061, B2 => n14063, A => n18039, ZN => 
                           n4070);
   U797 : BUF_X1 port map( A => n4182, Z => n17719);
   U798 : BUF_X1 port map( A => n4226, Z => n17659);
   U799 : BUF_X1 port map( A => n4182, Z => n17718);
   U800 : BUF_X1 port map( A => n4226, Z => n17658);
   U801 : BUF_X1 port map( A => n4117, Z => n17803);
   U802 : BUF_X1 port map( A => n4117, Z => n17802);
   U803 : BUF_X1 port map( A => n4108, Z => n17815);
   U804 : BUF_X1 port map( A => n4108, Z => n17814);
   U805 : BUF_X1 port map( A => n12562, Z => n16361);
   U806 : BUF_X1 port map( A => n12573, Z => n16334);
   U807 : BUF_X1 port map( A => n12568, Z => n16346);
   U808 : BUF_X1 port map( A => n12538, Z => n16406);
   U809 : BUF_X1 port map( A => n12548, Z => n16382);
   U810 : BUF_X1 port map( A => n12604, Z => n16274);
   U811 : BUF_X1 port map( A => n12587, Z => n16310);
   U812 : BUF_X1 port map( A => n12592, Z => n16298);
   U813 : BUF_X1 port map( A => n12597, Z => n16286);
   U814 : BUF_X1 port map( A => n12613, Z => n16262);
   U815 : BUF_X1 port map( A => n12629, Z => n16223);
   U816 : BUF_X1 port map( A => n12562, Z => n16362);
   U817 : BUF_X1 port map( A => n12573, Z => n16335);
   U818 : BUF_X1 port map( A => n12568, Z => n16347);
   U819 : BUF_X1 port map( A => n12538, Z => n16407);
   U820 : BUF_X1 port map( A => n12548, Z => n16383);
   U821 : BUF_X1 port map( A => n12604, Z => n16275);
   U822 : BUF_X1 port map( A => n12587, Z => n16311);
   U823 : BUF_X1 port map( A => n12592, Z => n16299);
   U824 : BUF_X1 port map( A => n12597, Z => n16287);
   U825 : BUF_X1 port map( A => n12613, Z => n16263);
   U826 : BUF_X1 port map( A => n12629, Z => n16224);
   U827 : BUF_X1 port map( A => n10567, Z => n16613);
   U828 : BUF_X1 port map( A => n10583, Z => n16586);
   U829 : BUF_X1 port map( A => n10576, Z => n16598);
   U830 : BUF_X1 port map( A => n10550, Z => n16634);
   U831 : BUF_X1 port map( A => n10543, Z => n16646);
   U832 : BUF_X1 port map( A => n10615, Z => n16538);
   U833 : BUF_X1 port map( A => n10622, Z => n16526);
   U834 : BUF_X1 port map( A => n10601, Z => n16562);
   U835 : BUF_X1 port map( A => n10608, Z => n16550);
   U836 : BUF_X1 port map( A => n10633, Z => n16514);
   U837 : BUF_X1 port map( A => n10656, Z => n16475);
   U838 : BUF_X1 port map( A => n10567, Z => n16614);
   U839 : BUF_X1 port map( A => n10583, Z => n16587);
   U840 : BUF_X1 port map( A => n10576, Z => n16599);
   U841 : BUF_X1 port map( A => n10550, Z => n16635);
   U842 : BUF_X1 port map( A => n10543, Z => n16647);
   U843 : BUF_X1 port map( A => n10615, Z => n16539);
   U844 : BUF_X1 port map( A => n10622, Z => n16527);
   U845 : BUF_X1 port map( A => n10601, Z => n16563);
   U846 : BUF_X1 port map( A => n10608, Z => n16551);
   U847 : BUF_X1 port map( A => n10633, Z => n16515);
   U848 : BUF_X1 port map( A => n10656, Z => n16476);
   U849 : BUF_X1 port map( A => n4162, Z => n17743);
   U850 : BUF_X1 port map( A => n4162, Z => n17742);
   U851 : BUF_X1 port map( A => n12617, Z => n16253);
   U852 : BUF_X1 port map( A => n12617, Z => n16254);
   U853 : BUF_X1 port map( A => n10639, Z => n16505);
   U854 : BUF_X1 port map( A => n10639, Z => n16506);
   U855 : OAI21_X1 port map( B1 => n14074, B2 => n14236, A => n18041, ZN => 
                           n4329);
   U856 : OAI21_X1 port map( B1 => n14073, B2 => n14236, A => n18041, ZN => 
                           n4326);
   U857 : OAI21_X1 port map( B1 => n14072, B2 => n14236, A => n18040, ZN => 
                           n4323);
   U858 : OAI21_X1 port map( B1 => n14070, B2 => n14236, A => n18041, ZN => 
                           n4320);
   U859 : OAI21_X1 port map( B1 => n12414, B2 => n14236, A => n18040, ZN => 
                           n4301);
   U860 : OAI21_X1 port map( B1 => n14058, B2 => n14236, A => n18040, ZN => 
                           n4298);
   U861 : OAI21_X1 port map( B1 => n14228, B2 => n14236, A => n18040, ZN => 
                           n4291);
   U862 : OAI21_X1 port map( B1 => n14226, B2 => n14236, A => n18040, ZN => 
                           n4288);
   U863 : OAI21_X1 port map( B1 => n14222, B2 => n14236, A => n18040, ZN => 
                           n4285);
   U864 : OAI21_X1 port map( B1 => n14221, B2 => n14236, A => n18040, ZN => 
                           n4282);
   U865 : OAI21_X1 port map( B1 => n14218, B2 => n14236, A => n18040, ZN => 
                           n4279);
   U866 : OAI21_X1 port map( B1 => n14215, B2 => n14236, A => n18040, ZN => 
                           n4275);
   U867 : BUF_X1 port map( A => n16454, Z => n16456);
   U868 : BUF_X1 port map( A => n16454, Z => n16457);
   U869 : BUF_X1 port map( A => n16455, Z => n16458);
   U870 : BUF_X1 port map( A => n16707, Z => n16709);
   U871 : BUF_X1 port map( A => n16707, Z => n16710);
   U872 : BUF_X1 port map( A => n16708, Z => n16711);
   U873 : BUF_X1 port map( A => n16716, Z => n16718);
   U874 : BUF_X1 port map( A => n16716, Z => n16719);
   U875 : BUF_X1 port map( A => n16717, Z => n16720);
   U876 : BUF_X1 port map( A => n12565, Z => n16355);
   U877 : BUF_X1 port map( A => n12565, Z => n16356);
   U878 : BUF_X1 port map( A => n10571, Z => n16607);
   U879 : BUF_X1 port map( A => n10571, Z => n16608);
   U880 : BUF_X1 port map( A => n12615, Z => n16259);
   U881 : BUF_X1 port map( A => n12615, Z => n16260);
   U882 : BUF_X1 port map( A => n10635, Z => n16511);
   U883 : BUF_X1 port map( A => n10635, Z => n16512);
   U884 : BUF_X1 port map( A => n12564, Z => n16358);
   U885 : BUF_X1 port map( A => n12564, Z => n16359);
   U886 : BUF_X1 port map( A => n10569, Z => n16610);
   U887 : BUF_X1 port map( A => n10569, Z => n16611);
   U888 : BUF_X1 port map( A => n4182, Z => n17720);
   U889 : BUF_X1 port map( A => n4226, Z => n17660);
   U890 : BUF_X1 port map( A => n4117, Z => n17804);
   U891 : BUF_X1 port map( A => n12622, Z => n16241);
   U892 : BUF_X1 port map( A => n12622, Z => n16242);
   U893 : BUF_X1 port map( A => n10646, Z => n16493);
   U894 : BUF_X1 port map( A => n10646, Z => n16494);
   U895 : BUF_X1 port map( A => n4152, Z => n17758);
   U896 : BUF_X1 port map( A => n4152, Z => n17757);
   U897 : BUF_X1 port map( A => n12581, Z => n16316);
   U898 : BUF_X1 port map( A => n12571, Z => n16340);
   U899 : BUF_X1 port map( A => n12552, Z => n16376);
   U900 : BUF_X1 port map( A => n12556, Z => n16367);
   U901 : BUF_X1 port map( A => n12607, Z => n16268);
   U902 : BUF_X1 port map( A => n12590, Z => n16304);
   U903 : BUF_X1 port map( A => n12601, Z => n16280);
   U904 : BUF_X1 port map( A => n12632, Z => n16217);
   U905 : BUF_X1 port map( A => n12627, Z => n16229);
   U906 : BUF_X1 port map( A => n12581, Z => n16317);
   U907 : BUF_X1 port map( A => n12571, Z => n16341);
   U908 : BUF_X1 port map( A => n12552, Z => n16377);
   U909 : BUF_X1 port map( A => n12556, Z => n16368);
   U910 : BUF_X1 port map( A => n12607, Z => n16269);
   U911 : BUF_X1 port map( A => n12590, Z => n16305);
   U912 : BUF_X1 port map( A => n12601, Z => n16281);
   U913 : BUF_X1 port map( A => n12632, Z => n16218);
   U914 : BUF_X1 port map( A => n12627, Z => n16230);
   U915 : BUF_X1 port map( A => n10587, Z => n16580);
   U916 : BUF_X1 port map( A => n10580, Z => n16592);
   U917 : BUF_X1 port map( A => n10554, Z => n16628);
   U918 : BUF_X1 port map( A => n10560, Z => n16619);
   U919 : BUF_X1 port map( A => n10619, Z => n16532);
   U920 : BUF_X1 port map( A => n10626, Z => n16520);
   U921 : BUF_X1 port map( A => n10605, Z => n16556);
   U922 : BUF_X1 port map( A => n10660, Z => n16469);
   U923 : BUF_X1 port map( A => n10653, Z => n16481);
   U924 : BUF_X1 port map( A => n10587, Z => n16581);
   U925 : BUF_X1 port map( A => n10580, Z => n16593);
   U926 : BUF_X1 port map( A => n10554, Z => n16629);
   U927 : BUF_X1 port map( A => n10560, Z => n16620);
   U928 : BUF_X1 port map( A => n10619, Z => n16533);
   U929 : BUF_X1 port map( A => n10626, Z => n16521);
   U930 : BUF_X1 port map( A => n10605, Z => n16557);
   U931 : BUF_X1 port map( A => n10660, Z => n16470);
   U932 : BUF_X1 port map( A => n10653, Z => n16482);
   U933 : BUF_X1 port map( A => n4192, Z => n17701);
   U934 : BUF_X1 port map( A => n4192, Z => n17700);
   U935 : BUF_X1 port map( A => n4108, Z => n17816);
   U936 : BUF_X1 port map( A => n12562, Z => n16363);
   U937 : BUF_X1 port map( A => n12573, Z => n16336);
   U938 : BUF_X1 port map( A => n12568, Z => n16348);
   U939 : BUF_X1 port map( A => n12538, Z => n16408);
   U940 : BUF_X1 port map( A => n12548, Z => n16384);
   U941 : BUF_X1 port map( A => n12604, Z => n16276);
   U942 : BUF_X1 port map( A => n12587, Z => n16312);
   U943 : BUF_X1 port map( A => n12592, Z => n16300);
   U944 : BUF_X1 port map( A => n12597, Z => n16288);
   U945 : BUF_X1 port map( A => n12613, Z => n16264);
   U946 : BUF_X1 port map( A => n12629, Z => n16225);
   U947 : BUF_X1 port map( A => n10567, Z => n16615);
   U948 : BUF_X1 port map( A => n10583, Z => n16588);
   U949 : BUF_X1 port map( A => n10576, Z => n16600);
   U950 : BUF_X1 port map( A => n10550, Z => n16636);
   U951 : BUF_X1 port map( A => n10543, Z => n16648);
   U952 : BUF_X1 port map( A => n10615, Z => n16540);
   U953 : BUF_X1 port map( A => n10622, Z => n16528);
   U954 : BUF_X1 port map( A => n10601, Z => n16564);
   U955 : BUF_X1 port map( A => n10608, Z => n16552);
   U956 : BUF_X1 port map( A => n10633, Z => n16516);
   U957 : BUF_X1 port map( A => n10656, Z => n16477);
   U958 : BUF_X1 port map( A => n4162, Z => n17744);
   U959 : BUF_X1 port map( A => n12572, Z => n16337);
   U960 : BUF_X1 port map( A => n12577, Z => n16325);
   U961 : BUF_X1 port map( A => n12567, Z => n16349);
   U962 : BUF_X1 port map( A => n12542, Z => n16397);
   U963 : BUF_X1 port map( A => n12603, Z => n16277);
   U964 : BUF_X1 port map( A => n12591, Z => n16301);
   U965 : BUF_X1 port map( A => n12596, Z => n16289);
   U966 : BUF_X1 port map( A => n12612, Z => n16265);
   U967 : BUF_X1 port map( A => n12618, Z => n16250);
   U968 : BUF_X1 port map( A => n12623, Z => n16238);
   U969 : BUF_X1 port map( A => n12572, Z => n16338);
   U970 : BUF_X1 port map( A => n12577, Z => n16326);
   U971 : BUF_X1 port map( A => n12567, Z => n16350);
   U972 : BUF_X1 port map( A => n12542, Z => n16398);
   U973 : BUF_X1 port map( A => n12603, Z => n16278);
   U974 : BUF_X1 port map( A => n12591, Z => n16302);
   U975 : BUF_X1 port map( A => n12596, Z => n16290);
   U976 : BUF_X1 port map( A => n12612, Z => n16266);
   U977 : BUF_X1 port map( A => n12618, Z => n16251);
   U978 : BUF_X1 port map( A => n12623, Z => n16239);
   U979 : BUF_X1 port map( A => n10582, Z => n16589);
   U980 : BUF_X1 port map( A => n10589, Z => n16577);
   U981 : BUF_X1 port map( A => n10575, Z => n16601);
   U982 : BUF_X1 port map( A => n10542, Z => n16649);
   U983 : BUF_X1 port map( A => n10614, Z => n16541);
   U984 : BUF_X1 port map( A => n10621, Z => n16529);
   U985 : BUF_X1 port map( A => n10607, Z => n16553);
   U986 : BUF_X1 port map( A => n10632, Z => n16517);
   U987 : BUF_X1 port map( A => n10641, Z => n16502);
   U988 : BUF_X1 port map( A => n10648, Z => n16490);
   U989 : BUF_X1 port map( A => n10582, Z => n16590);
   U990 : BUF_X1 port map( A => n10589, Z => n16578);
   U991 : BUF_X1 port map( A => n10575, Z => n16602);
   U992 : BUF_X1 port map( A => n10542, Z => n16650);
   U993 : BUF_X1 port map( A => n10614, Z => n16542);
   U994 : BUF_X1 port map( A => n10621, Z => n16530);
   U995 : BUF_X1 port map( A => n10607, Z => n16554);
   U996 : BUF_X1 port map( A => n10632, Z => n16518);
   U997 : BUF_X1 port map( A => n10641, Z => n16503);
   U998 : BUF_X1 port map( A => n10648, Z => n16491);
   U999 : BUF_X1 port map( A => n12575, Z => n16331);
   U1000 : BUF_X1 port map( A => n12550, Z => n16379);
   U1001 : BUF_X1 port map( A => n12606, Z => n16271);
   U1002 : BUF_X1 port map( A => n12621, Z => n16244);
   U1003 : BUF_X1 port map( A => n12575, Z => n16332);
   U1004 : BUF_X1 port map( A => n12550, Z => n16380);
   U1005 : BUF_X1 port map( A => n12606, Z => n16272);
   U1006 : BUF_X1 port map( A => n12621, Z => n16245);
   U1007 : BUF_X1 port map( A => n10592, Z => n16571);
   U1008 : BUF_X1 port map( A => n10624, Z => n16523);
   U1009 : BUF_X1 port map( A => n10644, Z => n16496);
   U1010 : BUF_X1 port map( A => n10592, Z => n16572);
   U1011 : BUF_X1 port map( A => n10624, Z => n16524);
   U1012 : BUF_X1 port map( A => n10644, Z => n16497);
   U1013 : BUF_X1 port map( A => n12580, Z => n16319);
   U1014 : BUF_X1 port map( A => n12545, Z => n16391);
   U1015 : BUF_X1 port map( A => n12555, Z => n16370);
   U1016 : BUF_X1 port map( A => n12589, Z => n16307);
   U1017 : BUF_X1 port map( A => n12631, Z => n16220);
   U1018 : BUF_X1 port map( A => n12580, Z => n16320);
   U1019 : BUF_X1 port map( A => n12545, Z => n16392);
   U1020 : BUF_X1 port map( A => n12555, Z => n16371);
   U1021 : BUF_X1 port map( A => n12589, Z => n16308);
   U1022 : BUF_X1 port map( A => n12631, Z => n16221);
   U1023 : BUF_X1 port map( A => n10585, Z => n16583);
   U1024 : BUF_X1 port map( A => n10552, Z => n16631);
   U1025 : BUF_X1 port map( A => n10558, Z => n16622);
   U1026 : BUF_X1 port map( A => n10617, Z => n16535);
   U1027 : BUF_X1 port map( A => n10603, Z => n16559);
   U1028 : BUF_X1 port map( A => n10658, Z => n16472);
   U1029 : BUF_X1 port map( A => n10585, Z => n16584);
   U1030 : BUF_X1 port map( A => n10552, Z => n16632);
   U1031 : BUF_X1 port map( A => n10558, Z => n16623);
   U1032 : BUF_X1 port map( A => n10617, Z => n16536);
   U1033 : BUF_X1 port map( A => n10603, Z => n16560);
   U1034 : BUF_X1 port map( A => n10658, Z => n16473);
   U1035 : BUF_X1 port map( A => n12570, Z => n16343);
   U1036 : BUF_X1 port map( A => n12594, Z => n16295);
   U1037 : BUF_X1 port map( A => n12599, Z => n16283);
   U1038 : BUF_X1 port map( A => n12626, Z => n16232);
   U1039 : BUF_X1 port map( A => n12570, Z => n16344);
   U1040 : BUF_X1 port map( A => n12594, Z => n16296);
   U1041 : BUF_X1 port map( A => n12599, Z => n16284);
   U1042 : BUF_X1 port map( A => n12626, Z => n16233);
   U1043 : BUF_X1 port map( A => n10578, Z => n16595);
   U1044 : BUF_X1 port map( A => n10545, Z => n16643);
   U1045 : BUF_X1 port map( A => n10610, Z => n16547);
   U1046 : BUF_X1 port map( A => n10651, Z => n16484);
   U1047 : BUF_X1 port map( A => n10578, Z => n16596);
   U1048 : BUF_X1 port map( A => n10545, Z => n16644);
   U1049 : BUF_X1 port map( A => n10610, Z => n16548);
   U1050 : BUF_X1 port map( A => n10651, Z => n16485);
   U1051 : BUF_X1 port map( A => n4164, Z => n17740);
   U1052 : BUF_X1 port map( A => n4164, Z => n17739);
   U1053 : BUF_X1 port map( A => n12617, Z => n16255);
   U1054 : BUF_X1 port map( A => n10639, Z => n16507);
   U1055 : BUF_X1 port map( A => n12565, Z => n16357);
   U1056 : BUF_X1 port map( A => n10571, Z => n16609);
   U1057 : BUF_X1 port map( A => n12615, Z => n16261);
   U1058 : BUF_X1 port map( A => n10635, Z => n16513);
   U1059 : BUF_X1 port map( A => n12564, Z => n16360);
   U1060 : BUF_X1 port map( A => n10569, Z => n16612);
   U1061 : BUF_X1 port map( A => n4152, Z => n17759);
   U1062 : BUF_X1 port map( A => n12622, Z => n16243);
   U1063 : BUF_X1 port map( A => n10646, Z => n16495);
   U1064 : BUF_X1 port map( A => n12607, Z => n16270);
   U1065 : BUF_X1 port map( A => n12581, Z => n16318);
   U1066 : BUF_X1 port map( A => n12571, Z => n16342);
   U1067 : BUF_X1 port map( A => n12552, Z => n16378);
   U1068 : BUF_X1 port map( A => n12556, Z => n16369);
   U1069 : BUF_X1 port map( A => n12590, Z => n16306);
   U1070 : BUF_X1 port map( A => n12601, Z => n16282);
   U1071 : BUF_X1 port map( A => n12632, Z => n16219);
   U1072 : BUF_X1 port map( A => n12627, Z => n16231);
   U1073 : BUF_X1 port map( A => n10587, Z => n16582);
   U1074 : BUF_X1 port map( A => n10626, Z => n16522);
   U1075 : BUF_X1 port map( A => n10580, Z => n16594);
   U1076 : BUF_X1 port map( A => n10554, Z => n16630);
   U1077 : BUF_X1 port map( A => n10560, Z => n16621);
   U1078 : BUF_X1 port map( A => n10619, Z => n16534);
   U1079 : BUF_X1 port map( A => n10605, Z => n16558);
   U1080 : BUF_X1 port map( A => n10660, Z => n16471);
   U1081 : BUF_X1 port map( A => n10653, Z => n16483);
   U1082 : BUF_X1 port map( A => n4192, Z => n17702);
   U1083 : BUF_X1 port map( A => n12575, Z => n16333);
   U1084 : BUF_X1 port map( A => n12550, Z => n16381);
   U1085 : BUF_X1 port map( A => n12606, Z => n16273);
   U1086 : BUF_X1 port map( A => n12621, Z => n16246);
   U1087 : BUF_X1 port map( A => n10592, Z => n16573);
   U1088 : BUF_X1 port map( A => n10624, Z => n16525);
   U1089 : BUF_X1 port map( A => n10644, Z => n16498);
   U1090 : BUF_X1 port map( A => n12572, Z => n16339);
   U1091 : BUF_X1 port map( A => n12577, Z => n16327);
   U1092 : BUF_X1 port map( A => n12567, Z => n16351);
   U1093 : BUF_X1 port map( A => n12542, Z => n16399);
   U1094 : BUF_X1 port map( A => n12603, Z => n16279);
   U1095 : BUF_X1 port map( A => n12591, Z => n16303);
   U1096 : BUF_X1 port map( A => n12596, Z => n16291);
   U1097 : BUF_X1 port map( A => n12612, Z => n16267);
   U1098 : BUF_X1 port map( A => n12618, Z => n16252);
   U1099 : BUF_X1 port map( A => n12623, Z => n16240);
   U1100 : BUF_X1 port map( A => n10582, Z => n16591);
   U1101 : BUF_X1 port map( A => n10589, Z => n16579);
   U1102 : BUF_X1 port map( A => n10575, Z => n16603);
   U1103 : BUF_X1 port map( A => n10542, Z => n16651);
   U1104 : BUF_X1 port map( A => n10614, Z => n16543);
   U1105 : BUF_X1 port map( A => n10621, Z => n16531);
   U1106 : BUF_X1 port map( A => n10607, Z => n16555);
   U1107 : BUF_X1 port map( A => n10632, Z => n16519);
   U1108 : BUF_X1 port map( A => n10641, Z => n16504);
   U1109 : BUF_X1 port map( A => n10648, Z => n16492);
   U1110 : BUF_X1 port map( A => n10585, Z => n16585);
   U1111 : BUF_X1 port map( A => n10552, Z => n16633);
   U1112 : BUF_X1 port map( A => n10558, Z => n16624);
   U1113 : BUF_X1 port map( A => n10617, Z => n16537);
   U1114 : BUF_X1 port map( A => n10603, Z => n16561);
   U1115 : BUF_X1 port map( A => n10658, Z => n16474);
   U1116 : BUF_X1 port map( A => n12580, Z => n16321);
   U1117 : BUF_X1 port map( A => n12545, Z => n16393);
   U1118 : BUF_X1 port map( A => n12555, Z => n16372);
   U1119 : BUF_X1 port map( A => n12589, Z => n16309);
   U1120 : BUF_X1 port map( A => n12631, Z => n16222);
   U1121 : BUF_X1 port map( A => n12570, Z => n16345);
   U1122 : BUF_X1 port map( A => n12594, Z => n16297);
   U1123 : BUF_X1 port map( A => n12599, Z => n16285);
   U1124 : BUF_X1 port map( A => n12626, Z => n16234);
   U1125 : BUF_X1 port map( A => n10578, Z => n16597);
   U1126 : BUF_X1 port map( A => n10545, Z => n16645);
   U1127 : BUF_X1 port map( A => n10610, Z => n16549);
   U1128 : BUF_X1 port map( A => n10651, Z => n16486);
   U1129 : BUF_X1 port map( A => n4164, Z => n17741);
   U1130 : OAI21_X1 port map( B1 => n14061, B2 => n14062, A => n18039, ZN => 
                           n4067);
   U1131 : OAI21_X1 port map( B1 => n14063, B2 => n14237, A => n18041, ZN => 
                           n4309);
   U1132 : OAI21_X1 port map( B1 => n14062, B2 => n14237, A => n18041, ZN => 
                           n4306);
   U1133 : BUF_X1 port map( A => n18054, Z => n18052);
   U1134 : BUF_X1 port map( A => n18054, Z => n18051);
   U1135 : NAND2_X1 port map( A1 => n14258, A2 => n14249, ZN => n14073);
   U1136 : NAND2_X1 port map( A1 => n14258, A2 => n14251, ZN => n14074);
   U1137 : BUF_X1 port map( A => n17822, Z => n17834);
   U1138 : AND2_X1 port map( A1 => n12489, A2 => n12437, ZN => n12440);
   U1139 : BUF_X1 port map( A => n16688, Z => n16695);
   U1140 : BUF_X1 port map( A => n16688, Z => n16694);
   U1141 : BUF_X1 port map( A => n17573, Z => n17580);
   U1142 : BUF_X1 port map( A => n17573, Z => n17579);
   U1143 : BUF_X1 port map( A => n18055, Z => n18050);
   U1144 : BUF_X1 port map( A => n18054, Z => n18053);
   U1145 : NAND2_X1 port map( A1 => n14085, A2 => n14086, ZN => n4112);
   U1146 : NAND2_X1 port map( A1 => n14085, A2 => n14088, ZN => n4121);
   U1147 : NAND2_X1 port map( A1 => n14085, A2 => n14103, ZN => n4128);
   U1148 : BUF_X1 port map( A => n16689, Z => n16696);
   U1149 : BUF_X1 port map( A => n17574, Z => n17581);
   U1150 : NAND2_X1 port map( A1 => n13919, A2 => n13920, ZN => n12540);
   U1151 : NAND2_X1 port map( A1 => n13925, A2 => n13920, ZN => n12546);
   U1152 : NAND2_X1 port map( A1 => n12438, A2 => n12439, ZN => n10538);
   U1153 : NAND2_X1 port map( A1 => n12443, A2 => n12439, ZN => n10547);
   U1154 : NAND2_X1 port map( A1 => n14107, A2 => n14085, ZN => n4248);
   U1155 : NAND2_X1 port map( A1 => n13936, A2 => n13918, ZN => n12566);
   U1156 : NAND2_X1 port map( A1 => n13946, A2 => n13918, ZN => n12576);
   U1157 : NAND2_X1 port map( A1 => n13917, A2 => n13918, ZN => n12541);
   U1158 : NAND2_X1 port map( A1 => n13953, A2 => n13918, ZN => n12595);
   U1159 : NAND2_X1 port map( A1 => n13960, A2 => n13918, ZN => n12616);
   U1160 : NAND2_X1 port map( A1 => n12455, A2 => n12437, ZN => n10573);
   U1161 : NAND2_X1 port map( A1 => n12465, A2 => n12437, ZN => n10594);
   U1162 : NAND2_X1 port map( A1 => n12436, A2 => n12437, ZN => n10540);
   U1163 : NAND2_X1 port map( A1 => n12472, A2 => n12437, ZN => n10612);
   U1164 : NAND2_X1 port map( A1 => n12479, A2 => n12437, ZN => n10637);
   U1165 : NAND2_X1 port map( A1 => n14087, A2 => n14088, ZN => n4110);
   U1166 : INV_X1 port map( A => n14201, ZN => n14088);
   U1167 : AND2_X1 port map( A1 => n13970, A2 => n13918, ZN => n13928);
   U1168 : INV_X1 port map( A => n14097, ZN => n14103);
   U1169 : BUF_X1 port map( A => n16455, Z => n16459);
   U1170 : BUF_X1 port map( A => n16708, Z => n16712);
   U1171 : BUF_X1 port map( A => n16717, Z => n16721);
   U1172 : AND2_X1 port map( A1 => n13926, A2 => n13918, ZN => n12553);
   U1173 : AND2_X1 port map( A1 => n13969, A2 => n13918, ZN => n12619);
   U1174 : AND2_X1 port map( A1 => n13955, A2 => n13918, ZN => n12628);
   U1175 : AND2_X1 port map( A1 => n12450, A2 => n12437, ZN => n10556);
   U1176 : AND2_X1 port map( A1 => n12488, A2 => n12437, ZN => n10642);
   U1177 : AND2_X1 port map( A1 => n12477, A2 => n12437, ZN => n10655);
   U1178 : AND2_X1 port map( A1 => n13920, A2 => n13923, ZN => n12537);
   U1179 : AND2_X1 port map( A1 => n12439, A2 => n12441, ZN => n10535);
   U1180 : BUF_X1 port map( A => n16688, Z => n16693);
   U1181 : BUF_X1 port map( A => n17573, Z => n17578);
   U1182 : AND2_X1 port map( A1 => n13931, A2 => n13920, ZN => n12561);
   U1183 : AND2_X1 port map( A1 => n13929, A2 => n13920, ZN => n12578);
   U1184 : AND2_X1 port map( A1 => n13928, A2 => n13920, ZN => n12543);
   U1185 : AND2_X1 port map( A1 => n13922, A2 => n13920, ZN => n12547);
   U1186 : AND2_X1 port map( A1 => n13933, A2 => n13920, ZN => n12586);
   U1187 : AND2_X1 port map( A1 => n12449, A2 => n12439, ZN => n10566);
   U1188 : AND2_X1 port map( A1 => n12447, A2 => n12439, ZN => n10590);
   U1189 : AND2_X1 port map( A1 => n12440, A2 => n12439, ZN => n10536);
   U1190 : AND2_X1 port map( A1 => n12445, A2 => n12439, ZN => n10549);
   U1191 : AND2_X1 port map( A1 => n12446, A2 => n12439, ZN => n10600);
   U1192 : BUF_X1 port map( A => n17545, Z => n17550);
   U1193 : BUF_X1 port map( A => n17559, Z => n17564);
   U1194 : BUF_X1 port map( A => n17586, Z => n17591);
   U1195 : BUF_X1 port map( A => n17600, Z => n17605);
   U1196 : BUF_X1 port map( A => n17614, Z => n17619);
   U1197 : BUF_X1 port map( A => n17531, Z => n17536);
   U1198 : BUF_X1 port map( A => n17547, Z => n17557);
   U1199 : BUF_X1 port map( A => n17561, Z => n17571);
   U1200 : BUF_X1 port map( A => n17588, Z => n17598);
   U1201 : BUF_X1 port map( A => n17602, Z => n17612);
   U1202 : BUF_X1 port map( A => n17616, Z => n17626);
   U1203 : BUF_X1 port map( A => n16689, Z => n16698);
   U1204 : BUF_X1 port map( A => n16689, Z => n16697);
   U1205 : BUF_X1 port map( A => n17533, Z => n17542);
   U1206 : BUF_X1 port map( A => n17547, Z => n17556);
   U1207 : BUF_X1 port map( A => n17561, Z => n17570);
   U1208 : BUF_X1 port map( A => n17588, Z => n17597);
   U1209 : BUF_X1 port map( A => n17602, Z => n17611);
   U1210 : BUF_X1 port map( A => n17616, Z => n17625);
   U1211 : BUF_X1 port map( A => n17532, Z => n17541);
   U1212 : BUF_X1 port map( A => n17546, Z => n17555);
   U1213 : BUF_X1 port map( A => n17560, Z => n17569);
   U1214 : BUF_X1 port map( A => n17574, Z => n17583);
   U1215 : BUF_X1 port map( A => n17587, Z => n17596);
   U1216 : BUF_X1 port map( A => n17601, Z => n17610);
   U1217 : BUF_X1 port map( A => n17615, Z => n17624);
   U1218 : BUF_X1 port map( A => n17532, Z => n17539);
   U1219 : BUF_X1 port map( A => n17546, Z => n17553);
   U1220 : BUF_X1 port map( A => n17560, Z => n17567);
   U1221 : BUF_X1 port map( A => n17587, Z => n17594);
   U1222 : BUF_X1 port map( A => n17601, Z => n17608);
   U1223 : BUF_X1 port map( A => n17615, Z => n17622);
   U1224 : BUF_X1 port map( A => n17532, Z => n17540);
   U1225 : BUF_X1 port map( A => n17546, Z => n17554);
   U1226 : BUF_X1 port map( A => n17560, Z => n17568);
   U1227 : BUF_X1 port map( A => n17574, Z => n17582);
   U1228 : BUF_X1 port map( A => n17587, Z => n17595);
   U1229 : BUF_X1 port map( A => n17601, Z => n17609);
   U1230 : BUF_X1 port map( A => n17615, Z => n17623);
   U1231 : BUF_X1 port map( A => n17531, Z => n17538);
   U1232 : BUF_X1 port map( A => n17545, Z => n17552);
   U1233 : BUF_X1 port map( A => n17559, Z => n17566);
   U1234 : BUF_X1 port map( A => n17586, Z => n17593);
   U1235 : BUF_X1 port map( A => n17600, Z => n17607);
   U1236 : BUF_X1 port map( A => n17614, Z => n17621);
   U1237 : BUF_X1 port map( A => n17531, Z => n17537);
   U1238 : BUF_X1 port map( A => n17545, Z => n17551);
   U1239 : BUF_X1 port map( A => n17559, Z => n17565);
   U1240 : BUF_X1 port map( A => n17586, Z => n17592);
   U1241 : BUF_X1 port map( A => n17600, Z => n17606);
   U1242 : BUF_X1 port map( A => n17614, Z => n17620);
   U1243 : BUF_X1 port map( A => n17533, Z => n17543);
   U1244 : BUF_X1 port map( A => n16690, Z => n16700);
   U1245 : BUF_X1 port map( A => n17575, Z => n17585);
   U1246 : BUF_X1 port map( A => n16690, Z => n16699);
   U1247 : BUF_X1 port map( A => n17575, Z => n17584);
   U1248 : BUF_X1 port map( A => n4367, Z => n17192);
   U1249 : OAI21_X1 port map( B1 => n14063, B2 => n14244, A => n18042, ZN => 
                           n4367);
   U1250 : BUF_X1 port map( A => n4423, Z => n16999);
   U1251 : OAI21_X1 port map( B1 => n14063, B2 => n14252, A => n18042, ZN => 
                           n4423);
   U1252 : OAI21_X1 port map( B1 => n14062, B2 => n14252, A => n18043, ZN => 
                           n4420);
   U1253 : OAI21_X1 port map( B1 => n14062, B2 => n14244, A => n18042, ZN => 
                           n4362);
   U1254 : BUF_X1 port map( A => n17533, Z => n17544);
   U1255 : BUF_X1 port map( A => n17547, Z => n17558);
   U1256 : BUF_X1 port map( A => n17561, Z => n17572);
   U1257 : BUF_X1 port map( A => n17588, Z => n17599);
   U1258 : BUF_X1 port map( A => n17602, Z => n17613);
   U1259 : INV_X1 port map( A => n14089, ZN => n14086);
   U1260 : INV_X1 port map( A => n14098, ZN => n14158);
   U1261 : BUF_X1 port map( A => n17616, Z => n17627);
   U1262 : BUF_X1 port map( A => n4062, Z => n18000);
   U1263 : BUF_X1 port map( A => n4456, Z => n16897);
   U1264 : BUF_X1 port map( A => n4467, Z => n16865);
   U1265 : BUF_X1 port map( A => n4062, Z => n18001);
   U1266 : BUF_X1 port map( A => n4467, Z => n16864);
   U1267 : BUF_X1 port map( A => n4456, Z => n16898);
   U1268 : BUF_X1 port map( A => n4467, Z => n16863);
   U1269 : BUF_X1 port map( A => n4385, Z => n17124);
   U1270 : BUF_X1 port map( A => n4379, Z => n17147);
   U1271 : BUF_X1 port map( A => n4359, Z => n17213);
   U1272 : BUF_X1 port map( A => n4356, Z => n17226);
   U1273 : BUF_X1 port map( A => n4351, Z => n17239);
   U1274 : BUF_X1 port map( A => n4348, Z => n17252);
   U1275 : BUF_X1 port map( A => n4341, Z => n17265);
   U1276 : BUF_X1 port map( A => n4338, Z => n17278);
   U1277 : BUF_X1 port map( A => n4335, Z => n17291);
   U1278 : BUF_X1 port map( A => n4332, Z => n17304);
   U1279 : BUF_X1 port map( A => n4385, Z => n17125);
   U1280 : BUF_X1 port map( A => n4379, Z => n17148);
   U1281 : BUF_X1 port map( A => n4359, Z => n17214);
   U1282 : BUF_X1 port map( A => n4356, Z => n17227);
   U1283 : BUF_X1 port map( A => n4351, Z => n17240);
   U1284 : BUF_X1 port map( A => n4348, Z => n17253);
   U1285 : BUF_X1 port map( A => n4341, Z => n17266);
   U1286 : BUF_X1 port map( A => n4338, Z => n17279);
   U1287 : BUF_X1 port map( A => n4335, Z => n17292);
   U1288 : BUF_X1 port map( A => n4332, Z => n17305);
   U1289 : BUF_X1 port map( A => n4441, Z => n16931);
   U1290 : BUF_X1 port map( A => n4417, Z => n17020);
   U1291 : BUF_X1 port map( A => n4412, Z => n17033);
   U1292 : BUF_X1 port map( A => n4409, Z => n17046);
   U1293 : BUF_X1 port map( A => n4406, Z => n17059);
   U1294 : BUF_X1 port map( A => n4401, Z => n17072);
   U1295 : BUF_X1 port map( A => n4398, Z => n17085);
   U1296 : BUF_X1 port map( A => n4391, Z => n17098);
   U1297 : BUF_X1 port map( A => n4388, Z => n17111);
   U1298 : BUF_X1 port map( A => n4441, Z => n16932);
   U1299 : BUF_X1 port map( A => n4417, Z => n17021);
   U1300 : BUF_X1 port map( A => n4412, Z => n17034);
   U1301 : BUF_X1 port map( A => n4409, Z => n17047);
   U1302 : BUF_X1 port map( A => n4406, Z => n17060);
   U1303 : BUF_X1 port map( A => n4401, Z => n17073);
   U1304 : BUF_X1 port map( A => n4398, Z => n17086);
   U1305 : BUF_X1 port map( A => n4391, Z => n17099);
   U1306 : BUF_X1 port map( A => n4388, Z => n17112);
   U1307 : BUF_X1 port map( A => n4059, Z => n18013);
   U1308 : BUF_X1 port map( A => n4059, Z => n18014);
   U1309 : BUF_X1 port map( A => n4317, Z => n17369);
   U1310 : BUF_X1 port map( A => n4317, Z => n17370);
   U1311 : BUF_X1 port map( A => n4426, Z => n16986);
   U1312 : BUF_X1 port map( A => n4312, Z => n17382);
   U1313 : BUF_X1 port map( A => n4426, Z => n16987);
   U1314 : BUF_X1 port map( A => n4312, Z => n17383);
   U1315 : BUF_X1 port map( A => n4062, Z => n18002);
   U1316 : BUF_X1 port map( A => n4456, Z => n16899);
   U1317 : BUF_X1 port map( A => n4385, Z => n17126);
   U1318 : BUF_X1 port map( A => n4379, Z => n17149);
   U1319 : BUF_X1 port map( A => n4359, Z => n17215);
   U1320 : BUF_X1 port map( A => n4356, Z => n17228);
   U1321 : BUF_X1 port map( A => n4351, Z => n17241);
   U1322 : BUF_X1 port map( A => n4348, Z => n17254);
   U1323 : BUF_X1 port map( A => n4341, Z => n17267);
   U1324 : BUF_X1 port map( A => n4338, Z => n17280);
   U1325 : BUF_X1 port map( A => n4335, Z => n17293);
   U1326 : BUF_X1 port map( A => n4332, Z => n17306);
   U1327 : BUF_X1 port map( A => n4441, Z => n16933);
   U1328 : BUF_X1 port map( A => n4417, Z => n17022);
   U1329 : BUF_X1 port map( A => n4412, Z => n17035);
   U1330 : BUF_X1 port map( A => n4409, Z => n17048);
   U1331 : BUF_X1 port map( A => n4406, Z => n17061);
   U1332 : BUF_X1 port map( A => n4401, Z => n17074);
   U1333 : BUF_X1 port map( A => n4398, Z => n17087);
   U1334 : BUF_X1 port map( A => n4391, Z => n17100);
   U1335 : BUF_X1 port map( A => n4388, Z => n17113);
   U1336 : BUF_X1 port map( A => n4059, Z => n18015);
   U1337 : BUF_X1 port map( A => n4317, Z => n17371);
   U1338 : BUF_X1 port map( A => n4426, Z => n16988);
   U1339 : BUF_X1 port map( A => n4312, Z => n17384);
   U1340 : INV_X1 port map( A => n16944, ZN => n16955);
   U1341 : INV_X1 port map( A => n16956, ZN => n16965);
   U1342 : INV_X1 port map( A => n16966, ZN => n16975);
   U1343 : INV_X1 port map( A => n17137, ZN => n17146);
   U1344 : INV_X1 port map( A => n17160, ZN => n17169);
   U1345 : INV_X1 port map( A => n16877, ZN => n16886);
   U1346 : INV_X1 port map( A => n16887, ZN => n16896);
   U1347 : INV_X1 port map( A => n16910, ZN => n16919);
   U1348 : INV_X1 port map( A => n4448, ZN => n16930);
   U1349 : INV_X1 port map( A => n16976, ZN => n16985);
   U1350 : INV_X1 port map( A => n17170, ZN => n17181);
   U1351 : INV_X1 port map( A => n17182, ZN => n17191);
   U1352 : BUF_X1 port map( A => n18055, Z => n18048);
   U1353 : BUF_X1 port map( A => n18048, Z => n18047);
   U1354 : BUF_X1 port map( A => n18049, Z => n18046);
   U1355 : BUF_X1 port map( A => n18049, Z => n18045);
   U1356 : BUF_X1 port map( A => n18055, Z => n18049);
   U1357 : BUF_X1 port map( A => n17822, Z => n17832);
   U1358 : BUF_X1 port map( A => n17821, Z => n17831);
   U1359 : BUF_X1 port map( A => n17821, Z => n17830);
   U1360 : BUF_X1 port map( A => n17821, Z => n17829);
   U1361 : BUF_X1 port map( A => n17820, Z => n17828);
   U1362 : BUF_X1 port map( A => n17820, Z => n17827);
   U1363 : BUF_X1 port map( A => n17820, Z => n17826);
   U1364 : BUF_X1 port map( A => n17822, Z => n17833);
   U1365 : NAND3_X1 port map( A1 => n14239, A2 => n14234, A3 => n14240, ZN => 
                           n14236);
   U1366 : OAI22_X1 port map( A1 => n14022, A2 => n14136, B1 => n14096, B2 => 
                           n14134, ZN => n4152);
   U1367 : OAI22_X1 port map( A1 => n14166, A2 => n14124, B1 => n14167, B2 => 
                           n14125, ZN => n4226);
   U1368 : OAI22_X1 port map( A1 => n14120, A2 => n14124, B1 => n14121, B2 => 
                           n14125, ZN => n4182);
   U1369 : OAI21_X1 port map( B1 => n14066, B2 => n14061, A => n18040, ZN => 
                           n4076);
   U1370 : OAI21_X1 port map( B1 => n14064, B2 => n14061, A => n18039, ZN => 
                           n4073);
   U1371 : NOR2_X1 port map( A1 => n14257, A2 => n14259, ZN => n14258);
   U1372 : NOR2_X1 port map( A1 => n14096, A2 => n14097, ZN => n4117);
   U1373 : BUF_X1 port map( A => n12624, Z => n16235);
   U1374 : BUF_X1 port map( A => n12624, Z => n16236);
   U1375 : INV_X1 port map( A => n14099, ZN => n14085);
   U1376 : AND3_X1 port map( A1 => n13980, A2 => n13963, A3 => n13962, ZN => 
                           n13920);
   U1377 : AND3_X1 port map( A1 => n12499, A2 => n12482, A3 => n12481, ZN => 
                           n12439);
   U1378 : INV_X1 port map( A => n14162, ZN => n4192);
   U1379 : OAI22_X1 port map( A1 => n14163, A2 => n14124, B1 => n14164, B2 => 
                           n14125, ZN => n14162);
   U1380 : OAI21_X1 port map( B1 => n14059, B2 => n14228, A => n18041, ZN => 
                           n4467);
   U1381 : OAI21_X1 port map( B1 => n14059, B2 => n12414, A => n18039, ZN => 
                           n4062);
   U1382 : OAI21_X1 port map( B1 => n14059, B2 => n14221, A => n18044, ZN => 
                           n4456);
   U1383 : BUF_X1 port map( A => n10523, Z => n16670);
   U1384 : BUF_X1 port map( A => n10517, Z => n16682);
   U1385 : BUF_X1 port map( A => n10662, Z => n16466);
   U1386 : BUF_X1 port map( A => n10649, Z => n16487);
   U1387 : BUF_X1 port map( A => n4153, Z => n17755);
   U1388 : BUF_X1 port map( A => n4153, Z => n17754);
   U1389 : BUF_X1 port map( A => n4198, Z => n17695);
   U1390 : BUF_X1 port map( A => n4198, Z => n17694);
   U1391 : BUF_X1 port map( A => n4233, Z => n17647);
   U1392 : BUF_X1 port map( A => n4233, Z => n17646);
   U1393 : BUF_X1 port map( A => n4207, Z => n17683);
   U1394 : BUF_X1 port map( A => n4207, Z => n17682);
   U1395 : BUF_X1 port map( A => n4220, Z => n17671);
   U1396 : BUF_X1 port map( A => n4220, Z => n17670);
   U1397 : BUF_X1 port map( A => n4142, Z => n17767);
   U1398 : BUF_X1 port map( A => n4189, Z => n17707);
   U1399 : BUF_X1 port map( A => n4142, Z => n17766);
   U1400 : BUF_X1 port map( A => n4189, Z => n17706);
   U1401 : BUF_X1 port map( A => n4171, Z => n17731);
   U1402 : BUF_X1 port map( A => n4124, Z => n17791);
   U1403 : BUF_X1 port map( A => n4131, Z => n17779);
   U1404 : BUF_X1 port map( A => n4171, Z => n17730);
   U1405 : BUF_X1 port map( A => n4124, Z => n17790);
   U1406 : BUF_X1 port map( A => n4131, Z => n17778);
   U1407 : BUF_X1 port map( A => n10663, Z => n16463);
   U1408 : BUF_X1 port map( A => n10649, Z => n16488);
   U1409 : BUF_X1 port map( A => n10519, Z => n16679);
   U1410 : BUF_X1 port map( A => n10662, Z => n16467);
   U1411 : BUF_X1 port map( A => n10523, Z => n16671);
   U1412 : BUF_X1 port map( A => n10517, Z => n16683);
   U1413 : NOR2_X1 port map( A1 => n14089, A2 => n14090, ZN => n4108);
   U1414 : BUF_X1 port map( A => n10519, Z => n16680);
   U1415 : BUF_X1 port map( A => n4058, Z => n18026);
   U1416 : BUF_X1 port map( A => n4058, Z => n18030);
   U1417 : BUF_X1 port map( A => n4058, Z => n18029);
   U1418 : BUF_X1 port map( A => n4058, Z => n18028);
   U1419 : BUF_X1 port map( A => n4058, Z => n18027);
   U1420 : BUF_X1 port map( A => n10510, Z => n16701);
   U1421 : INV_X1 port map( A => n14034, ZN => n14033);
   U1422 : BUF_X1 port map( A => n4058, Z => n18031);
   U1423 : BUF_X1 port map( A => n12522, Z => n16427);
   U1424 : BUF_X1 port map( A => n12522, Z => n16428);
   U1425 : BUF_X1 port map( A => n10510, Z => n16702);
   U1426 : OAI21_X1 port map( B1 => n14074, B2 => n14241, A => n18042, ZN => 
                           n4385);
   U1427 : OAI21_X1 port map( B1 => n14072, B2 => n14241, A => n18042, ZN => 
                           n4379);
   U1428 : OAI21_X1 port map( B1 => n12414, B2 => n14241, A => n18042, ZN => 
                           n4359);
   U1429 : OAI21_X1 port map( B1 => n14058, B2 => n14241, A => n18041, ZN => 
                           n4356);
   U1430 : OAI21_X1 port map( B1 => n14228, B2 => n14241, A => n18042, ZN => 
                           n4351);
   U1431 : OAI21_X1 port map( B1 => n14226, B2 => n14241, A => n18041, ZN => 
                           n4348);
   U1432 : OAI21_X1 port map( B1 => n14222, B2 => n14241, A => n18039, ZN => 
                           n4341);
   U1433 : OAI21_X1 port map( B1 => n14221, B2 => n14241, A => n18041, ZN => 
                           n4338);
   U1434 : OAI21_X1 port map( B1 => n14218, B2 => n14241, A => n18041, ZN => 
                           n4335);
   U1435 : OAI21_X1 port map( B1 => n14215, B2 => n14241, A => n18041, ZN => 
                           n4332);
   U1436 : BUF_X1 port map( A => n7537, Z => n16731);
   U1437 : BUF_X1 port map( A => n7537, Z => n16732);
   U1438 : BUF_X1 port map( A => n7537, Z => n16733);
   U1439 : BUF_X1 port map( A => n7537, Z => n16734);
   U1440 : BUF_X1 port map( A => n7537, Z => n16735);
   U1441 : BUF_X1 port map( A => n7537, Z => n16736);
   U1442 : BUF_X1 port map( A => n7428, Z => n16737);
   U1443 : BUF_X1 port map( A => n7428, Z => n16738);
   U1444 : BUF_X1 port map( A => n7428, Z => n16739);
   U1445 : BUF_X1 port map( A => n7428, Z => n16740);
   U1446 : BUF_X1 port map( A => n7428, Z => n16741);
   U1447 : BUF_X1 port map( A => n7428, Z => n16742);
   U1448 : BUF_X1 port map( A => n7319, Z => n16743);
   U1449 : BUF_X1 port map( A => n7319, Z => n16744);
   U1450 : BUF_X1 port map( A => n7319, Z => n16745);
   U1451 : BUF_X1 port map( A => n7319, Z => n16746);
   U1452 : BUF_X1 port map( A => n7319, Z => n16747);
   U1453 : BUF_X1 port map( A => n7319, Z => n16748);
   U1454 : BUF_X1 port map( A => n7205, Z => n16749);
   U1455 : BUF_X1 port map( A => n7205, Z => n16750);
   U1456 : BUF_X1 port map( A => n7205, Z => n16751);
   U1457 : BUF_X1 port map( A => n7205, Z => n16752);
   U1458 : BUF_X1 port map( A => n7205, Z => n16753);
   U1459 : BUF_X1 port map( A => n7205, Z => n16754);
   U1460 : BUF_X1 port map( A => n7096, Z => n16755);
   U1461 : BUF_X1 port map( A => n7096, Z => n16756);
   U1462 : BUF_X1 port map( A => n7096, Z => n16757);
   U1463 : BUF_X1 port map( A => n7096, Z => n16758);
   U1464 : BUF_X1 port map( A => n7096, Z => n16759);
   U1465 : BUF_X1 port map( A => n7096, Z => n16760);
   U1466 : BUF_X1 port map( A => n6987, Z => n16761);
   U1467 : BUF_X1 port map( A => n6987, Z => n16762);
   U1468 : BUF_X1 port map( A => n6987, Z => n16763);
   U1469 : BUF_X1 port map( A => n6987, Z => n16764);
   U1470 : BUF_X1 port map( A => n6987, Z => n16765);
   U1471 : BUF_X1 port map( A => n6987, Z => n16766);
   U1472 : BUF_X1 port map( A => n6878, Z => n16767);
   U1473 : BUF_X1 port map( A => n6878, Z => n16768);
   U1474 : BUF_X1 port map( A => n6878, Z => n16769);
   U1475 : BUF_X1 port map( A => n6878, Z => n16770);
   U1476 : BUF_X1 port map( A => n6878, Z => n16771);
   U1477 : BUF_X1 port map( A => n6878, Z => n16772);
   U1478 : BUF_X1 port map( A => n6769, Z => n16773);
   U1479 : BUF_X1 port map( A => n6769, Z => n16774);
   U1480 : BUF_X1 port map( A => n6769, Z => n16775);
   U1481 : BUF_X1 port map( A => n6769, Z => n16776);
   U1482 : BUF_X1 port map( A => n6769, Z => n16777);
   U1483 : BUF_X1 port map( A => n6769, Z => n16778);
   U1484 : BUF_X1 port map( A => n6635, Z => n16779);
   U1485 : BUF_X1 port map( A => n6635, Z => n16780);
   U1486 : BUF_X1 port map( A => n6635, Z => n16781);
   U1487 : BUF_X1 port map( A => n6635, Z => n16782);
   U1488 : BUF_X1 port map( A => n6635, Z => n16783);
   U1489 : BUF_X1 port map( A => n6635, Z => n16784);
   U1490 : BUF_X1 port map( A => n6448, Z => n16785);
   U1491 : BUF_X1 port map( A => n6448, Z => n16786);
   U1492 : BUF_X1 port map( A => n6448, Z => n16787);
   U1493 : BUF_X1 port map( A => n6448, Z => n16788);
   U1494 : BUF_X1 port map( A => n6448, Z => n16789);
   U1495 : BUF_X1 port map( A => n6448, Z => n16790);
   U1496 : BUF_X1 port map( A => n6261, Z => n16791);
   U1497 : BUF_X1 port map( A => n6261, Z => n16792);
   U1498 : BUF_X1 port map( A => n6261, Z => n16793);
   U1499 : BUF_X1 port map( A => n6261, Z => n16794);
   U1500 : BUF_X1 port map( A => n6261, Z => n16795);
   U1501 : BUF_X1 port map( A => n6261, Z => n16796);
   U1502 : BUF_X1 port map( A => n6076, Z => n16797);
   U1503 : BUF_X1 port map( A => n6076, Z => n16798);
   U1504 : BUF_X1 port map( A => n6076, Z => n16799);
   U1505 : BUF_X1 port map( A => n6076, Z => n16800);
   U1506 : BUF_X1 port map( A => n6076, Z => n16801);
   U1507 : BUF_X1 port map( A => n6076, Z => n16802);
   U1508 : BUF_X1 port map( A => n5889, Z => n16803);
   U1509 : BUF_X1 port map( A => n5889, Z => n16804);
   U1510 : BUF_X1 port map( A => n5889, Z => n16805);
   U1511 : BUF_X1 port map( A => n5889, Z => n16806);
   U1512 : BUF_X1 port map( A => n5889, Z => n16807);
   U1513 : BUF_X1 port map( A => n5889, Z => n16808);
   U1514 : BUF_X1 port map( A => n5717, Z => n16809);
   U1515 : BUF_X1 port map( A => n5717, Z => n16810);
   U1516 : BUF_X1 port map( A => n5717, Z => n16811);
   U1517 : BUF_X1 port map( A => n5717, Z => n16812);
   U1518 : BUF_X1 port map( A => n5717, Z => n16813);
   U1519 : BUF_X1 port map( A => n5717, Z => n16814);
   U1520 : BUF_X1 port map( A => n5530, Z => n16815);
   U1521 : BUF_X1 port map( A => n5530, Z => n16816);
   U1522 : BUF_X1 port map( A => n5530, Z => n16817);
   U1523 : BUF_X1 port map( A => n5530, Z => n16818);
   U1524 : BUF_X1 port map( A => n5530, Z => n16819);
   U1525 : BUF_X1 port map( A => n5530, Z => n16820);
   U1526 : BUF_X1 port map( A => n5343, Z => n16821);
   U1527 : BUF_X1 port map( A => n5343, Z => n16822);
   U1528 : BUF_X1 port map( A => n5343, Z => n16823);
   U1529 : BUF_X1 port map( A => n5343, Z => n16824);
   U1530 : BUF_X1 port map( A => n5343, Z => n16825);
   U1531 : BUF_X1 port map( A => n5343, Z => n16826);
   U1532 : BUF_X1 port map( A => n5157, Z => n16827);
   U1533 : BUF_X1 port map( A => n5157, Z => n16828);
   U1534 : BUF_X1 port map( A => n5157, Z => n16829);
   U1535 : BUF_X1 port map( A => n5157, Z => n16830);
   U1536 : BUF_X1 port map( A => n5157, Z => n16831);
   U1537 : BUF_X1 port map( A => n5157, Z => n16832);
   U1538 : BUF_X1 port map( A => n5040, Z => n16833);
   U1539 : BUF_X1 port map( A => n5040, Z => n16834);
   U1540 : BUF_X1 port map( A => n5040, Z => n16835);
   U1541 : BUF_X1 port map( A => n5040, Z => n16836);
   U1542 : BUF_X1 port map( A => n5040, Z => n16837);
   U1543 : BUF_X1 port map( A => n5040, Z => n16838);
   U1544 : BUF_X1 port map( A => n4924, Z => n16839);
   U1545 : BUF_X1 port map( A => n4924, Z => n16840);
   U1546 : BUF_X1 port map( A => n4924, Z => n16841);
   U1547 : BUF_X1 port map( A => n4924, Z => n16842);
   U1548 : BUF_X1 port map( A => n4924, Z => n16843);
   U1549 : BUF_X1 port map( A => n4924, Z => n16844);
   U1550 : BUF_X1 port map( A => n4791, Z => n16845);
   U1551 : BUF_X1 port map( A => n4791, Z => n16846);
   U1552 : BUF_X1 port map( A => n4791, Z => n16847);
   U1553 : BUF_X1 port map( A => n4791, Z => n16848);
   U1554 : BUF_X1 port map( A => n4791, Z => n16849);
   U1555 : BUF_X1 port map( A => n4791, Z => n16850);
   U1556 : BUF_X1 port map( A => n4664, Z => n16851);
   U1557 : BUF_X1 port map( A => n4664, Z => n16852);
   U1558 : BUF_X1 port map( A => n4664, Z => n16853);
   U1559 : BUF_X1 port map( A => n4664, Z => n16854);
   U1560 : BUF_X1 port map( A => n4664, Z => n16855);
   U1561 : BUF_X1 port map( A => n4664, Z => n16856);
   U1562 : BUF_X1 port map( A => n4533, Z => n16857);
   U1563 : BUF_X1 port map( A => n4533, Z => n16858);
   U1564 : BUF_X1 port map( A => n4533, Z => n16859);
   U1565 : BUF_X1 port map( A => n4533, Z => n16860);
   U1566 : BUF_X1 port map( A => n4533, Z => n16861);
   U1567 : BUF_X1 port map( A => n4533, Z => n16862);
   U1568 : BUF_X1 port map( A => n4278, Z => n17512);
   U1569 : BUF_X1 port map( A => n4278, Z => n17513);
   U1570 : BUF_X1 port map( A => n4278, Z => n17514);
   U1571 : BUF_X1 port map( A => n4278, Z => n17515);
   U1572 : BUF_X1 port map( A => n4278, Z => n17516);
   U1573 : BUF_X1 port map( A => n4278, Z => n17517);
   U1574 : BUF_X1 port map( A => n10510, Z => n16706);
   U1575 : BUF_X1 port map( A => n10510, Z => n16705);
   U1576 : BUF_X1 port map( A => n10510, Z => n16704);
   U1577 : BUF_X1 port map( A => n10510, Z => n16703);
   U1578 : BUF_X1 port map( A => n7652, Z => n16725);
   U1579 : BUF_X1 port map( A => n7652, Z => n16726);
   U1580 : BUF_X1 port map( A => n7652, Z => n16727);
   U1581 : BUF_X1 port map( A => n7652, Z => n16728);
   U1582 : BUF_X1 port map( A => n7652, Z => n16729);
   U1583 : BUF_X1 port map( A => n12338, Z => n16436);
   U1584 : BUF_X1 port map( A => n12338, Z => n16437);
   U1585 : BUF_X1 port map( A => n12338, Z => n16438);
   U1586 : BUF_X1 port map( A => n12184, Z => n16442);
   U1587 : BUF_X1 port map( A => n12184, Z => n16443);
   U1588 : BUF_X1 port map( A => n12184, Z => n16444);
   U1589 : BUF_X1 port map( A => n12029, Z => n16448);
   U1590 : BUF_X1 port map( A => n12029, Z => n16449);
   U1591 : BUF_X1 port map( A => n12029, Z => n16450);
   U1592 : OAI21_X1 port map( B1 => n14074, B2 => n14248, A => n18044, ZN => 
                           n4441);
   U1593 : OAI21_X1 port map( B1 => n12414, B2 => n14248, A => n18043, ZN => 
                           n4417);
   U1594 : OAI21_X1 port map( B1 => n14058, B2 => n14248, A => n18043, ZN => 
                           n4412);
   U1595 : OAI21_X1 port map( B1 => n14228, B2 => n14248, A => n18043, ZN => 
                           n4409);
   U1596 : OAI21_X1 port map( B1 => n14226, B2 => n14248, A => n18043, ZN => 
                           n4406);
   U1597 : OAI21_X1 port map( B1 => n14222, B2 => n14248, A => n18043, ZN => 
                           n4401);
   U1598 : OAI21_X1 port map( B1 => n14221, B2 => n14248, A => n18042, ZN => 
                           n4398);
   U1599 : OAI21_X1 port map( B1 => n14218, B2 => n14248, A => n18043, ZN => 
                           n4391);
   U1600 : OAI21_X1 port map( B1 => n14215, B2 => n14248, A => n18042, ZN => 
                           n4388);
   U1601 : BUF_X1 port map( A => n12523, Z => n16424);
   U1602 : BUF_X1 port map( A => n12523, Z => n16425);
   U1603 : BUF_X1 port map( A => n10520, Z => n16677);
   U1604 : BUF_X1 port map( A => n10520, Z => n16676);
   U1605 : BUF_X1 port map( A => n10663, Z => n16464);
   U1606 : OAI21_X1 port map( B1 => n14058, B2 => n14059, A => n18039, ZN => 
                           n4059);
   U1607 : BUF_X1 port map( A => n12524, Z => n16421);
   U1608 : BUF_X1 port map( A => n12519, Z => n16433);
   U1609 : BUF_X1 port map( A => n12524, Z => n16422);
   U1610 : BUF_X1 port map( A => n12519, Z => n16434);
   U1611 : BUF_X1 port map( A => n10522, Z => n16674);
   U1612 : BUF_X1 port map( A => n10516, Z => n16686);
   U1613 : BUF_X1 port map( A => n10522, Z => n16673);
   U1614 : BUF_X1 port map( A => n10516, Z => n16685);
   U1615 : BUF_X1 port map( A => n4153, Z => n17756);
   U1616 : BUF_X1 port map( A => n4198, Z => n17696);
   U1617 : BUF_X1 port map( A => n4233, Z => n17648);
   U1618 : BUF_X1 port map( A => n4207, Z => n17684);
   U1619 : BUF_X1 port map( A => n4220, Z => n17672);
   U1620 : BUF_X1 port map( A => n4142, Z => n17768);
   U1621 : BUF_X1 port map( A => n4189, Z => n17708);
   U1622 : BUF_X1 port map( A => n4168, Z => n17737);
   U1623 : BUF_X1 port map( A => n4237, Z => n17641);
   U1624 : BUF_X1 port map( A => n4168, Z => n17736);
   U1625 : BUF_X1 port map( A => n4237, Z => n17640);
   U1626 : BUF_X1 port map( A => n4230, Z => n17653);
   U1627 : BUF_X1 port map( A => n4230, Z => n17652);
   U1628 : BUF_X1 port map( A => n4159, Z => n17749);
   U1629 : BUF_X1 port map( A => n4211, Z => n17677);
   U1630 : BUF_X1 port map( A => n4159, Z => n17748);
   U1631 : BUF_X1 port map( A => n4211, Z => n17676);
   U1632 : BUF_X1 port map( A => n4135, Z => n17773);
   U1633 : BUF_X1 port map( A => n4135, Z => n17772);
   U1634 : BUF_X1 port map( A => n4175, Z => n17725);
   U1635 : BUF_X1 port map( A => n4186, Z => n17713);
   U1636 : BUF_X1 port map( A => n4175, Z => n17724);
   U1637 : BUF_X1 port map( A => n4186, Z => n17712);
   U1638 : BUF_X1 port map( A => n4150, Z => n17761);
   U1639 : BUF_X1 port map( A => n4150, Z => n17760);
   U1640 : BUF_X1 port map( A => n4161, Z => n17746);
   U1641 : BUF_X1 port map( A => n4195, Z => n17698);
   U1642 : BUF_X1 port map( A => n4161, Z => n17745);
   U1643 : BUF_X1 port map( A => n4195, Z => n17697);
   U1644 : BUF_X1 port map( A => n4232, Z => n17650);
   U1645 : BUF_X1 port map( A => n4232, Z => n17649);
   U1646 : BUF_X1 port map( A => n4206, Z => n17686);
   U1647 : BUF_X1 port map( A => n4206, Z => n17685);
   U1648 : BUF_X1 port map( A => n4188, Z => n17710);
   U1649 : BUF_X1 port map( A => n4219, Z => n17674);
   U1650 : BUF_X1 port map( A => n4188, Z => n17709);
   U1651 : BUF_X1 port map( A => n4219, Z => n17673);
   U1652 : BUF_X1 port map( A => n4141, Z => n17770);
   U1653 : BUF_X1 port map( A => n4181, Z => n17722);
   U1654 : BUF_X1 port map( A => n4225, Z => n17662);
   U1655 : BUF_X1 port map( A => n4239, Z => n17638);
   U1656 : BUF_X1 port map( A => n4114, Z => n17806);
   U1657 : BUF_X1 port map( A => n4141, Z => n17769);
   U1658 : BUF_X1 port map( A => n4181, Z => n17721);
   U1659 : BUF_X1 port map( A => n4225, Z => n17661);
   U1660 : BUF_X1 port map( A => n4239, Z => n17637);
   U1661 : BUF_X1 port map( A => n4114, Z => n17805);
   U1662 : BUF_X1 port map( A => n4200, Z => n17692);
   U1663 : BUF_X1 port map( A => n4209, Z => n17680);
   U1664 : BUF_X1 port map( A => n4200, Z => n17691);
   U1665 : BUF_X1 port map( A => n4209, Z => n17679);
   U1666 : BUF_X1 port map( A => n4157, Z => n17752);
   U1667 : BUF_X1 port map( A => n4235, Z => n17644);
   U1668 : BUF_X1 port map( A => n4228, Z => n17656);
   U1669 : BUF_X1 port map( A => n4157, Z => n17751);
   U1670 : BUF_X1 port map( A => n4235, Z => n17643);
   U1671 : BUF_X1 port map( A => n4228, Z => n17655);
   U1672 : BUF_X1 port map( A => n12633, Z => n16214);
   U1673 : BUF_X1 port map( A => n12633, Z => n16215);
   U1674 : BUF_X1 port map( A => n12525, Z => n16418);
   U1675 : BUF_X1 port map( A => n12520, Z => n16430);
   U1676 : BUF_X1 port map( A => n12525, Z => n16419);
   U1677 : BUF_X1 port map( A => n12520, Z => n16431);
   U1678 : BUF_X1 port map( A => n4124, Z => n17792);
   U1679 : BUF_X1 port map( A => n4131, Z => n17780);
   U1680 : BUF_X1 port map( A => n4171, Z => n17732);
   U1681 : BUF_X1 port map( A => n4184, Z => n17716);
   U1682 : BUF_X1 port map( A => n4119, Z => n17800);
   U1683 : BUF_X1 port map( A => n4126, Z => n17788);
   U1684 : BUF_X1 port map( A => n4133, Z => n17776);
   U1685 : BUF_X1 port map( A => n4184, Z => n17715);
   U1686 : BUF_X1 port map( A => n4119, Z => n17799);
   U1687 : BUF_X1 port map( A => n4126, Z => n17787);
   U1688 : BUF_X1 port map( A => n4133, Z => n17775);
   U1689 : BUF_X1 port map( A => n4173, Z => n17728);
   U1690 : BUF_X1 port map( A => n4242, Z => n17632);
   U1691 : BUF_X1 port map( A => n4173, Z => n17727);
   U1692 : BUF_X1 port map( A => n4242, Z => n17631);
   U1693 : BUF_X1 port map( A => n4170, Z => n17734);
   U1694 : BUF_X1 port map( A => n4107, Z => n17818);
   U1695 : BUF_X1 port map( A => n4123, Z => n17794);
   U1696 : BUF_X1 port map( A => n4130, Z => n17782);
   U1697 : BUF_X1 port map( A => n4170, Z => n17733);
   U1698 : BUF_X1 port map( A => n4107, Z => n17817);
   U1699 : BUF_X1 port map( A => n4123, Z => n17793);
   U1700 : BUF_X1 port map( A => n4130, Z => n17781);
   U1701 : BUF_X1 port map( A => n4148, Z => n17764);
   U1702 : BUF_X1 port map( A => n4191, Z => n17704);
   U1703 : BUF_X1 port map( A => n4222, Z => n17668);
   U1704 : BUF_X1 port map( A => n4148, Z => n17763);
   U1705 : BUF_X1 port map( A => n4191, Z => n17703);
   U1706 : BUF_X1 port map( A => n4222, Z => n17667);
   U1707 : BUF_X1 port map( A => n12522, Z => n16429);
   U1708 : NOR2_X1 port map( A1 => n13975, A2 => n13976, ZN => n13970);
   U1709 : NOR2_X1 port map( A1 => n12494, A2 => n12495, ZN => n12489);
   U1710 : BUF_X1 port map( A => n12523, Z => n16426);
   U1711 : BUF_X1 port map( A => n12634, Z => n16212);
   U1712 : BUF_X1 port map( A => n12634, Z => n16211);
   U1713 : NAND2_X1 port map( A1 => n14260, A2 => n14253, ZN => n14215);
   U1714 : NAND2_X1 port map( A1 => n13932, A2 => n13960, ZN => n12615);
   U1715 : BUF_X1 port map( A => n12524, Z => n16423);
   U1716 : BUF_X1 port map( A => n12519, Z => n16435);
   U1717 : BUF_X1 port map( A => n10520, Z => n16678);
   U1718 : NAND2_X1 port map( A1 => n14260, A2 => n14251, ZN => n14222);
   U1719 : NAND2_X1 port map( A1 => n14260, A2 => n14249, ZN => n14221);
   U1720 : NAND2_X1 port map( A1 => n14253, A2 => n14250, ZN => n14226);
   U1721 : NAND2_X1 port map( A1 => n14260, A2 => n14254, ZN => n14218);
   U1722 : NAND2_X1 port map( A1 => n14254, A2 => n14250, ZN => n14228);
   U1723 : BUF_X1 port map( A => n4161, Z => n17747);
   U1724 : BUF_X1 port map( A => n4195, Z => n17699);
   U1725 : BUF_X1 port map( A => n4232, Z => n17651);
   U1726 : BUF_X1 port map( A => n4168, Z => n17738);
   U1727 : BUF_X1 port map( A => n4237, Z => n17642);
   U1728 : BUF_X1 port map( A => n4230, Z => n17654);
   U1729 : BUF_X1 port map( A => n4206, Z => n17687);
   U1730 : BUF_X1 port map( A => n4188, Z => n17711);
   U1731 : BUF_X1 port map( A => n4219, Z => n17675);
   U1732 : BUF_X1 port map( A => n4159, Z => n17750);
   U1733 : BUF_X1 port map( A => n4211, Z => n17678);
   U1734 : BUF_X1 port map( A => n4141, Z => n17771);
   U1735 : BUF_X1 port map( A => n4181, Z => n17723);
   U1736 : BUF_X1 port map( A => n4225, Z => n17663);
   U1737 : BUF_X1 port map( A => n4239, Z => n17639);
   U1738 : BUF_X1 port map( A => n4114, Z => n17807);
   U1739 : BUF_X1 port map( A => n10522, Z => n16675);
   U1740 : BUF_X1 port map( A => n10516, Z => n16687);
   U1741 : BUF_X1 port map( A => n4135, Z => n17774);
   U1742 : BUF_X1 port map( A => n4200, Z => n17693);
   U1743 : BUF_X1 port map( A => n4209, Z => n17681);
   U1744 : BUF_X1 port map( A => n4175, Z => n17726);
   U1745 : BUF_X1 port map( A => n4186, Z => n17714);
   U1746 : BUF_X1 port map( A => n4157, Z => n17753);
   U1747 : BUF_X1 port map( A => n4235, Z => n17645);
   U1748 : BUF_X1 port map( A => n4228, Z => n17657);
   U1749 : BUF_X1 port map( A => n4150, Z => n17762);
   U1750 : NAND2_X1 port map( A1 => n14251, A2 => n14250, ZN => n12414);
   U1751 : BUF_X1 port map( A => n12624, Z => n16237);
   U1752 : BUF_X1 port map( A => n12633, Z => n16216);
   U1753 : BUF_X1 port map( A => n12525, Z => n16420);
   U1754 : BUF_X1 port map( A => n12520, Z => n16432);
   U1755 : BUF_X1 port map( A => n4184, Z => n17717);
   U1756 : BUF_X1 port map( A => n4119, Z => n17801);
   U1757 : BUF_X1 port map( A => n4126, Z => n17789);
   U1758 : BUF_X1 port map( A => n4133, Z => n17777);
   U1759 : BUF_X1 port map( A => n4173, Z => n17729);
   U1760 : BUF_X1 port map( A => n4242, Z => n17633);
   U1761 : BUF_X1 port map( A => n4123, Z => n17795);
   U1762 : BUF_X1 port map( A => n4130, Z => n17783);
   U1763 : BUF_X1 port map( A => n4170, Z => n17735);
   U1764 : BUF_X1 port map( A => n4107, Z => n17819);
   U1765 : BUF_X1 port map( A => n4148, Z => n17765);
   U1766 : BUF_X1 port map( A => n4191, Z => n17705);
   U1767 : BUF_X1 port map( A => n4222, Z => n17669);
   U1768 : NAND2_X1 port map( A1 => n12452, A2 => n12479, ZN => n10635);
   U1769 : NAND2_X1 port map( A1 => n14249, A2 => n14250, ZN => n14058);
   U1770 : NAND2_X1 port map( A1 => n14138, A2 => n14205, ZN => n14089);
   U1771 : NAND2_X1 port map( A1 => n14137, A2 => n14205, ZN => n14098);
   U1772 : OAI21_X1 port map( B1 => n14066, B2 => n14237, A => n18041, ZN => 
                           n4317);
   U1773 : BUF_X1 port map( A => n12634, Z => n16213);
   U1774 : BUF_X1 port map( A => n4088, Z => n17835);
   U1775 : OAI21_X1 port map( B1 => n14059, B2 => n14074, A => n18040, ZN => 
                           n4088);
   U1776 : BUF_X1 port map( A => n4085, Z => n17857);
   U1777 : OAI21_X1 port map( B1 => n14059, B2 => n14073, A => n18040, ZN => 
                           n4085);
   U1778 : BUF_X1 port map( A => n4082, Z => n17879);
   U1779 : OAI21_X1 port map( B1 => n14059, B2 => n14072, A => n18040, ZN => 
                           n4082);
   U1780 : BUF_X1 port map( A => n4079, Z => n17901);
   U1781 : OAI21_X1 port map( B1 => n14059, B2 => n14070, A => n18039, ZN => 
                           n4079);
   U1782 : OAI21_X1 port map( B1 => n14064, B2 => n14252, A => n18043, ZN => 
                           n4426);
   U1783 : OAI21_X1 port map( B1 => n14064, B2 => n14237, A => n18041, ZN => 
                           n4312);
   U1784 : INV_X1 port map( A => n14207, ZN => n14197);
   U1785 : NAND2_X1 port map( A1 => n14245, A2 => n14067, ZN => n14244);
   U1786 : INV_X1 port map( A => n14241, ZN => n14245);
   U1787 : NAND2_X1 port map( A1 => n14256, A2 => n14067, ZN => n14252);
   U1788 : INV_X1 port map( A => n14248, ZN => n14256);
   U1789 : NAND2_X1 port map( A1 => n14238, A2 => n14067, ZN => n14237);
   U1790 : INV_X1 port map( A => n14236, ZN => n14238);
   U1791 : NAND2_X1 port map( A1 => n14258, A2 => n14253, ZN => n14070);
   U1792 : NAND2_X1 port map( A1 => n14143, A2 => n14205, ZN => n14097);
   U1793 : NAND2_X1 port map( A1 => n14202, A2 => n14205, ZN => n14201);
   U1794 : NAND2_X1 port map( A1 => n14067, A2 => n14068, ZN => n14061);
   U1795 : INV_X1 port map( A => n14059, ZN => n14068);
   U1796 : NAND2_X1 port map( A1 => n14258, A2 => n14254, ZN => n14072);
   U1797 : INV_X1 port map( A => n14183, ZN => n14176);
   U1798 : AND2_X1 port map( A1 => n14000, A2 => n14001, ZN => n14004);
   U1799 : INV_X1 port map( A => n14096, ZN => n14087);
   U1800 : NAND2_X1 port map( A1 => n13946, A2 => n13932, ZN => n12575);
   U1801 : NAND2_X1 port map( A1 => n13926, A2 => n13932, ZN => n12550);
   U1802 : NAND2_X1 port map( A1 => n13936, A2 => n13932, ZN => n12606);
   U1803 : NAND2_X1 port map( A1 => n13955, A2 => n13932, ZN => n12621);
   U1804 : NAND2_X1 port map( A1 => n13969, A2 => n13932, ZN => n12622);
   U1805 : BUF_X1 port map( A => n10649, Z => n16489);
   U1806 : NAND2_X1 port map( A1 => n12465, A2 => n12452, ZN => n10592);
   U1807 : NAND2_X1 port map( A1 => n12455, A2 => n12452, ZN => n10624);
   U1808 : NAND2_X1 port map( A1 => n12477, A2 => n12452, ZN => n10644);
   U1809 : NAND2_X1 port map( A1 => n12488, A2 => n12452, ZN => n10646);
   U1810 : BUF_X1 port map( A => n10662, Z => n16468);
   U1811 : BUF_X1 port map( A => n10523, Z => n16672);
   U1812 : BUF_X1 port map( A => n10517, Z => n16684);
   U1813 : AND2_X1 port map( A1 => n12463, A2 => n12456, ZN => n12465);
   U1814 : AND2_X1 port map( A1 => n13944, A2 => n13937, ZN => n13946);
   U1815 : BUF_X1 port map( A => n10519, Z => n16681);
   U1816 : AND2_X1 port map( A1 => n12444, A2 => n12480, ZN => n12455);
   U1817 : AND2_X1 port map( A1 => n13921, A2 => n13961, ZN => n13936);
   U1818 : INV_X1 port map( A => n14253, ZN => n14062);
   U1819 : AND2_X1 port map( A1 => n13970, A2 => n13932, ZN => n13925);
   U1820 : AND2_X1 port map( A1 => n13957, A2 => n13937, ZN => n13960);
   U1821 : AND2_X1 port map( A1 => n12489, A2 => n12452, ZN => n12443);
   U1822 : AND2_X1 port map( A1 => n12474, A2 => n12456, ZN => n12479);
   U1823 : BUF_X1 port map( A => n10663, Z => n16465);
   U1824 : NAND2_X1 port map( A1 => n12451, A2 => n12479, ZN => n10626);
   U1825 : NAND2_X1 port map( A1 => n18044, A2 => n14000, ZN => n14001);
   U1826 : INV_X1 port map( A => n14254, ZN => n14063);
   U1827 : NAND2_X1 port map( A1 => n13927, A2 => n13960, ZN => n12607);
   U1828 : NAND2_X1 port map( A1 => n13935, A2 => n13969, ZN => n12617);
   U1829 : NAND2_X1 port map( A1 => n12454, A2 => n12488, ZN => n10639);
   U1830 : INV_X1 port map( A => n14134, ZN => n14094);
   U1831 : AND2_X1 port map( A1 => n12463, A2 => n12480, ZN => n12472);
   U1832 : AND2_X1 port map( A1 => n13944, A2 => n13961, ZN => n13953);
   U1833 : AND2_X1 port map( A1 => n13920, A2 => n13961, ZN => n13917);
   U1834 : AND2_X1 port map( A1 => n12439, A2 => n12480, ZN => n12436);
   U1835 : AND2_X1 port map( A1 => n13921, A2 => n13937, ZN => n13926);
   U1836 : INV_X1 port map( A => n14066, ZN => n14251);
   U1837 : NAND2_X1 port map( A1 => n12465, A2 => n12451, ZN => n10585);
   U1838 : NAND2_X1 port map( A1 => n12450, A2 => n12451, ZN => n10552);
   U1839 : NAND2_X1 port map( A1 => n12455, A2 => n12451, ZN => n10558);
   U1840 : NAND2_X1 port map( A1 => n12477, A2 => n12451, ZN => n10617);
   U1841 : NAND2_X1 port map( A1 => n12472, A2 => n12451, ZN => n10603);
   U1842 : NAND2_X1 port map( A1 => n12436, A2 => n12451, ZN => n10658);
   U1843 : NAND2_X1 port map( A1 => n13946, A2 => n13927, ZN => n12580);
   U1844 : NAND2_X1 port map( A1 => n13926, A2 => n13927, ZN => n12545);
   U1845 : NAND2_X1 port map( A1 => n13936, A2 => n13927, ZN => n12555);
   U1846 : NAND2_X1 port map( A1 => n13953, A2 => n13927, ZN => n12589);
   U1847 : NAND2_X1 port map( A1 => n13917, A2 => n13927, ZN => n12631);
   U1848 : AND2_X1 port map( A1 => n12475, A2 => n12454, ZN => n12445);
   U1849 : AND2_X1 port map( A1 => n13961, A2 => n13957, ZN => n13969);
   U1850 : AND2_X1 port map( A1 => n12480, A2 => n12474, ZN => n12488);
   U1851 : INV_X1 port map( A => n14064, ZN => n14249);
   U1852 : AND2_X1 port map( A1 => n13958, A2 => n13927, ZN => n13929);
   U1853 : AND2_X1 port map( A1 => n13958, A2 => n13935, ZN => n13922);
   U1854 : NAND2_X1 port map( A1 => n12463, A2 => n12440, ZN => n10619);
   U1855 : NAND2_X1 port map( A1 => n12463, A2 => n12443, ZN => n10610);
   U1856 : AND2_X1 port map( A1 => n12444, A2 => n12456, ZN => n12450);
   U1857 : AND2_X1 port map( A1 => n12439, A2 => n12456, ZN => n12477);
   U1858 : INV_X1 port map( A => n14131, ZN => n14104);
   U1859 : NAND2_X1 port map( A1 => n13944, A2 => n13925, ZN => n12594);
   U1860 : NAND2_X1 port map( A1 => n13922, A2 => n13957, ZN => n12601);
   U1861 : NAND2_X1 port map( A1 => n13929, A2 => n13957, ZN => n12599);
   U1862 : NAND2_X1 port map( A1 => n13928, A2 => n13957, ZN => n12627);
   U1863 : NAND2_X1 port map( A1 => n13925, A2 => n13957, ZN => n12626);
   U1864 : NAND2_X1 port map( A1 => n13936, A2 => n13935, ZN => n12565);
   U1865 : NAND2_X1 port map( A1 => n13946, A2 => n13935, ZN => n12581);
   U1866 : NAND2_X1 port map( A1 => n13926, A2 => n13935, ZN => n12556);
   U1867 : NAND2_X1 port map( A1 => n13953, A2 => n13935, ZN => n12590);
   U1868 : NAND2_X1 port map( A1 => n13917, A2 => n13935, ZN => n12632);
   U1869 : NAND2_X1 port map( A1 => n12455, A2 => n12454, ZN => n10571);
   U1870 : NAND2_X1 port map( A1 => n12465, A2 => n12454, ZN => n10587);
   U1871 : NAND2_X1 port map( A1 => n12450, A2 => n12454, ZN => n10560);
   U1872 : NAND2_X1 port map( A1 => n12472, A2 => n12454, ZN => n10605);
   U1873 : NAND2_X1 port map( A1 => n12436, A2 => n12454, ZN => n10660);
   U1874 : NAND2_X1 port map( A1 => n12445, A2 => n12463, ZN => n10580);
   U1875 : NAND2_X1 port map( A1 => n12447, A2 => n12463, ZN => n10578);
   U1876 : AND2_X1 port map( A1 => n13958, A2 => n13932, ZN => n13931);
   U1877 : AND2_X1 port map( A1 => n12475, A2 => n12452, ZN => n12449);
   U1878 : NAND2_X1 port map( A1 => n12444, A2 => n12441, ZN => n10569);
   U1879 : NAND2_X1 port map( A1 => n12444, A2 => n12449, ZN => n10554);
   U1880 : NAND2_X1 port map( A1 => n12444, A2 => n12445, ZN => n10545);
   U1881 : NAND2_X1 port map( A1 => n13922, A2 => n13944, ZN => n12571);
   U1882 : NAND2_X1 port map( A1 => n13929, A2 => n13944, ZN => n12570);
   U1883 : INV_X1 port map( A => n14145, ZN => n14107);
   U1884 : NAND2_X1 port map( A1 => n12440, A2 => n12474, ZN => n10653);
   U1885 : NAND2_X1 port map( A1 => n12443, A2 => n12474, ZN => n10651);
   U1886 : NAND2_X1 port map( A1 => n14108, A2 => n14085, ZN => n4164);
   U1887 : NAND2_X1 port map( A1 => n13921, A2 => n13931, ZN => n12552);
   U1888 : NAND2_X1 port map( A1 => n13921, A2 => n13923, ZN => n12564);
   U1889 : AND2_X1 port map( A1 => n12489, A2 => n12451, ZN => n12441);
   U1890 : AND2_X1 port map( A1 => n13970, A2 => n13927, ZN => n13923);
   U1891 : AND2_X1 port map( A1 => n13917, A2 => n13932, ZN => n12577);
   U1892 : AND2_X1 port map( A1 => n13953, A2 => n13932, ZN => n12629);
   U1893 : AND2_X1 port map( A1 => n12436, A2 => n12452, ZN => n10589);
   U1894 : AND2_X1 port map( A1 => n12450, A2 => n12452, ZN => n10550);
   U1895 : AND2_X1 port map( A1 => n12472, A2 => n12452, ZN => n10656);
   U1896 : AND2_X1 port map( A1 => n13970, A2 => n13935, ZN => n13919);
   U1897 : AND2_X1 port map( A1 => n12489, A2 => n12454, ZN => n12438);
   U1898 : AND2_X1 port map( A1 => n12475, A2 => n12451, ZN => n12447);
   U1899 : AND2_X1 port map( A1 => n13920, A2 => n13937, ZN => n13955);
   U1900 : AND2_X1 port map( A1 => n12451, A2 => n12488, ZN => n10632);
   U1901 : AND2_X1 port map( A1 => n13927, A2 => n13969, ZN => n12612);
   U1902 : AND2_X1 port map( A1 => n13935, A2 => n13960, ZN => n12604);
   U1903 : AND2_X1 port map( A1 => n12454, A2 => n12479, ZN => n10622);
   U1904 : AND2_X1 port map( A1 => n12463, A2 => n12441, ZN => n10601);
   U1905 : AND2_X1 port map( A1 => n12463, A2 => n12438, ZN => n10607);
   U1906 : AND2_X1 port map( A1 => n13955, A2 => n13927, ZN => n12592);
   U1907 : AND2_X1 port map( A1 => n13955, A2 => n13935, ZN => n12618);
   U1908 : AND2_X1 port map( A1 => n12477, A2 => n12454, ZN => n10641);
   U1909 : AND2_X1 port map( A1 => n13944, A2 => n13923, ZN => n12587);
   U1910 : AND2_X1 port map( A1 => n13944, A2 => n13919, ZN => n12591);
   U1911 : AND2_X1 port map( A1 => n13944, A2 => n13928, ZN => n12596);
   U1912 : AND2_X1 port map( A1 => n12444, A2 => n12438, ZN => n10567);
   U1913 : AND2_X1 port map( A1 => n12444, A2 => n12440, ZN => n10575);
   U1914 : AND2_X1 port map( A1 => n12444, A2 => n12443, ZN => n10576);
   U1915 : AND2_X1 port map( A1 => n12444, A2 => n12447, ZN => n10542);
   U1916 : AND2_X1 port map( A1 => n12444, A2 => n12446, ZN => n10543);
   U1917 : AND2_X1 port map( A1 => n13921, A2 => n13919, ZN => n12562);
   U1918 : AND2_X1 port map( A1 => n13921, A2 => n13928, ZN => n12567);
   U1919 : AND2_X1 port map( A1 => n13921, A2 => n13925, ZN => n12568);
   U1920 : AND2_X1 port map( A1 => n13921, A2 => n13922, ZN => n12538);
   U1921 : AND2_X1 port map( A1 => n13921, A2 => n13929, ZN => n12542);
   U1922 : AND2_X1 port map( A1 => n13921, A2 => n13933, ZN => n12548);
   U1923 : AND2_X1 port map( A1 => n13931, A2 => n13957, ZN => n12603);
   U1924 : AND2_X1 port map( A1 => n13933, A2 => n13957, ZN => n12597);
   U1925 : AND2_X1 port map( A1 => n13923, A2 => n13957, ZN => n12613);
   U1926 : AND2_X1 port map( A1 => n13919, A2 => n13957, ZN => n12623);
   U1927 : AND2_X1 port map( A1 => n12446, A2 => n12463, ZN => n10582);
   U1928 : AND2_X1 port map( A1 => n12449, A2 => n12463, ZN => n10583);
   U1929 : AND2_X1 port map( A1 => n13933, A2 => n13944, ZN => n12572);
   U1930 : AND2_X1 port map( A1 => n13931, A2 => n13944, ZN => n12573);
   U1931 : AND2_X1 port map( A1 => n12445, A2 => n12474, ZN => n10614);
   U1932 : AND2_X1 port map( A1 => n12446, A2 => n12474, ZN => n10615);
   U1933 : AND2_X1 port map( A1 => n12449, A2 => n12474, ZN => n10621);
   U1934 : AND2_X1 port map( A1 => n12447, A2 => n12474, ZN => n10608);
   U1935 : AND2_X1 port map( A1 => n12441, A2 => n12474, ZN => n10633);
   U1936 : AND2_X1 port map( A1 => n12438, A2 => n12474, ZN => n10648);
   U1937 : AND2_X1 port map( A1 => n14108, A2 => n14087, ZN => n4162);
   U1938 : BUF_X1 port map( A => n4462, Z => n16877);
   U1939 : OAI21_X1 port map( B1 => n14059, B2 => n14226, A => n18044, ZN => 
                           n4462);
   U1940 : BUF_X1 port map( A => n4459, Z => n16887);
   U1941 : OAI21_X1 port map( B1 => n14059, B2 => n14222, A => n18044, ZN => 
                           n4459);
   U1942 : BUF_X1 port map( A => n4451, Z => n16910);
   U1943 : OAI21_X1 port map( B1 => n14059, B2 => n14218, A => n18044, ZN => 
                           n4451);
   U1944 : OAI21_X1 port map( B1 => n14059, B2 => n14215, A => n18043, ZN => 
                           n4448);
   U1945 : BUF_X1 port map( A => n4382, Z => n17137);
   U1946 : OAI21_X1 port map( B1 => n14073, B2 => n14241, A => n18042, ZN => 
                           n4382);
   U1947 : BUF_X1 port map( A => n4376, Z => n17160);
   U1948 : OAI21_X1 port map( B1 => n14070, B2 => n14241, A => n18042, ZN => 
                           n4376);
   U1949 : BUF_X1 port map( A => n4438, Z => n16944);
   U1950 : OAI21_X1 port map( B1 => n14073, B2 => n14248, A => n18043, ZN => 
                           n4438);
   U1951 : BUF_X1 port map( A => n4435, Z => n16956);
   U1952 : OAI21_X1 port map( B1 => n14072, B2 => n14248, A => n18043, ZN => 
                           n4435);
   U1953 : BUF_X1 port map( A => n4432, Z => n16966);
   U1954 : OAI21_X1 port map( B1 => n14070, B2 => n14248, A => n18043, ZN => 
                           n4432);
   U1955 : BUF_X1 port map( A => n4373, Z => n17170);
   U1956 : OAI21_X1 port map( B1 => n14066, B2 => n14244, A => n18042, ZN => 
                           n4373);
   U1957 : BUF_X1 port map( A => n4429, Z => n16976);
   U1958 : OAI21_X1 port map( B1 => n14066, B2 => n14252, A => n18043, ZN => 
                           n4429);
   U1959 : BUF_X1 port map( A => n4370, Z => n17182);
   U1960 : OAI21_X1 port map( B1 => n14064, B2 => n14244, A => n18042, ZN => 
                           n4370);
   U1961 : AND2_X1 port map( A1 => n13958, A2 => n13918, ZN => n13933);
   U1962 : AND2_X1 port map( A1 => n12475, A2 => n12437, ZN => n12446);
   U1963 : INV_X1 port map( A => n14133, ZN => n14022);
   U1964 : BUF_X1 port map( A => n10425, Z => n16707);
   U1965 : BUF_X1 port map( A => n10315, Z => n16716);
   U1966 : BUF_X1 port map( A => n11868, Z => n16454);
   U1967 : INV_X1 port map( A => n14180, ZN => n14182);
   U1968 : INV_X1 port map( A => n14204, ZN => n14208);
   U1969 : BUF_X1 port map( A => n10425, Z => n16708);
   U1970 : BUF_X1 port map( A => n10315, Z => n16717);
   U1971 : BUF_X1 port map( A => n11868, Z => n16455);
   U1972 : BUF_X1 port map( A => n10511, Z => n16688);
   U1973 : BUF_X1 port map( A => n4273, Z => n17533);
   U1974 : BUF_X1 port map( A => n4270, Z => n17547);
   U1975 : BUF_X1 port map( A => n4267, Z => n17561);
   U1976 : BUF_X1 port map( A => n10511, Z => n16689);
   U1977 : BUF_X1 port map( A => n4273, Z => n17532);
   U1978 : BUF_X1 port map( A => n4270, Z => n17546);
   U1979 : BUF_X1 port map( A => n4267, Z => n17560);
   U1980 : BUF_X1 port map( A => n4273, Z => n17531);
   U1981 : BUF_X1 port map( A => n4270, Z => n17545);
   U1982 : BUF_X1 port map( A => n4267, Z => n17559);
   U1983 : BUF_X1 port map( A => n4262, Z => n17573);
   U1984 : BUF_X1 port map( A => n4259, Z => n17588);
   U1985 : BUF_X1 port map( A => n4262, Z => n17574);
   U1986 : BUF_X1 port map( A => n4259, Z => n17587);
   U1987 : BUF_X1 port map( A => n4259, Z => n17586);
   U1988 : BUF_X1 port map( A => n4256, Z => n17602);
   U1989 : BUF_X1 port map( A => n4251, Z => n17616);
   U1990 : BUF_X1 port map( A => n4256, Z => n17601);
   U1991 : BUF_X1 port map( A => n4251, Z => n17615);
   U1992 : BUF_X1 port map( A => n4256, Z => n17600);
   U1993 : BUF_X1 port map( A => n4251, Z => n17614);
   U1994 : BUF_X1 port map( A => n4090, Z => n17822);
   U1995 : BUF_X1 port map( A => n10511, Z => n16690);
   U1996 : BUF_X1 port map( A => n4262, Z => n17575);
   U1997 : INV_X1 port map( A => n18032, ZN => n18054);
   U1998 : INV_X1 port map( A => n18032, ZN => n18055);
   U1999 : BUF_X1 port map( A => n12302, Z => n16439);
   U2000 : BUF_X1 port map( A => n12302, Z => n16440);
   U2001 : BUF_X1 port map( A => n12302, Z => n16441);
   U2002 : BUF_X1 port map( A => n12149, Z => n16445);
   U2003 : BUF_X1 port map( A => n12149, Z => n16446);
   U2004 : BUF_X1 port map( A => n12149, Z => n16447);
   U2005 : BUF_X1 port map( A => n11996, Z => n16451);
   U2006 : BUF_X1 port map( A => n11996, Z => n16452);
   U2007 : BUF_X1 port map( A => n11996, Z => n16453);
   U2008 : BUF_X1 port map( A => n10400, Z => n16714);
   U2009 : BUF_X1 port map( A => n10400, Z => n16713);
   U2010 : BUF_X1 port map( A => n11843, Z => n16461);
   U2011 : BUF_X1 port map( A => n11843, Z => n16460);
   U2012 : BUF_X1 port map( A => n10290, Z => n16723);
   U2013 : BUF_X1 port map( A => n10290, Z => n16722);
   U2014 : BUF_X1 port map( A => n11843, Z => n16462);
   U2015 : BUF_X1 port map( A => n10290, Z => n16724);
   U2016 : BUF_X1 port map( A => n10400, Z => n16715);
   U2017 : BUF_X1 port map( A => n4090, Z => n17821);
   U2018 : BUF_X1 port map( A => n4090, Z => n17820);
   U2019 : NOR3_X1 port map( A1 => n14174, A2 => N9924, A3 => n14173, ZN => 
                           n14151);
   U2020 : NAND4_X1 port map( A1 => N9924, A2 => n14173, A3 => n14174, A4 => 
                           n14020, ZN => n14096);
   U2021 : NAND3_X1 port map( A1 => n14247, A2 => n14234, A3 => n14240, ZN => 
                           n14248);
   U2022 : NOR2_X1 port map( A1 => n17825, A2 => n14005, ZN => n14034);
   U2023 : NAND3_X1 port map( A1 => n14240, A2 => n14247, A3 => N276, ZN => 
                           n14059);
   U2024 : NOR3_X1 port map( A1 => n14006, A2 => n14231, A3 => n14266, ZN => 
                           n14240);
   U2025 : INV_X1 port map( A => n14232, ZN => n14266);
   U2026 : NOR3_X1 port map( A1 => N9922, A2 => N9924, A3 => n14174, ZN => 
                           n14091);
   U2027 : NAND4_X1 port map( A1 => n14231, A2 => n14232, A3 => n14233, A4 => 
                           n14234, ZN => n12415);
   U2028 : BUF_X1 port map( A => n12527, Z => n16413);
   U2029 : BUF_X1 port map( A => n12527, Z => n16412);
   U2030 : BUF_X1 port map( A => n10525, Z => n16665);
   U2031 : BUF_X1 port map( A => n10525, Z => n16664);
   U2032 : BUF_X1 port map( A => n12527, Z => n16414);
   U2033 : BUF_X1 port map( A => n10525, Z => n16666);
   U2034 : OAI22_X1 port map( A1 => n14135, A2 => n14136, B1 => n14096, B2 => 
                           n14131, ZN => n4153);
   U2035 : INV_X1 port map( A => n14129, ZN => n14135);
   U2036 : OAI22_X1 port map( A1 => n14144, A2 => n14136, B1 => n14145, B2 => 
                           n14096, ZN => n4161);
   U2037 : OAI22_X1 port map( A1 => n14172, A2 => n14142, B1 => n14089, B2 => 
                           n14096, ZN => n4195);
   U2038 : OAI22_X1 port map( A1 => n14172, A2 => n14101, B1 => n14098, B2 => 
                           n14096, ZN => n4198);
   U2039 : OAI22_X1 port map( A1 => n14181, A2 => n14208, B1 => n14207, B2 => 
                           n14184, ZN => n4232);
   U2040 : OAI22_X1 port map( A1 => n14208, A2 => n14185, B1 => n14207, B2 => 
                           n14186, ZN => n4233);
   U2041 : OAI22_X1 port map( A1 => n14185, A2 => n14182, B1 => n14183, B2 => 
                           n14186, ZN => n4206);
   U2042 : OAI22_X1 port map( A1 => n14181, A2 => n14182, B1 => n14183, B2 => 
                           n14184, ZN => n4207);
   U2043 : OAI22_X1 port map( A1 => n14163, A2 => n14115, B1 => n14164, B2 => 
                           n14117, ZN => n4188);
   U2044 : OAI22_X1 port map( A1 => n14163, A2 => n14122, B1 => n14164, B2 => 
                           n14123, ZN => n4219);
   U2045 : NAND2_X1 port map( A1 => N9925, A2 => n14197, ZN => n14164);
   U2046 : OAI22_X1 port map( A1 => n14120, A2 => n14159, B1 => n14121, B2 => 
                           n14160, ZN => n4220);
   U2047 : OAI22_X1 port map( A1 => n14124, A2 => n14116, B1 => n14125, B2 => 
                           n14118, ZN => n4141);
   U2048 : OAI22_X1 port map( A1 => n14159, A2 => n14116, B1 => n14160, B2 => 
                           n14118, ZN => n4181);
   U2049 : OAI22_X1 port map( A1 => n14122, A2 => n14116, B1 => n14123, B2 => 
                           n14118, ZN => n4239);
   U2050 : OAI22_X1 port map( A1 => n14122, A2 => n14166, B1 => n14123, B2 => 
                           n14167, ZN => n4189);
   U2051 : OAI22_X1 port map( A1 => n14159, A2 => n14166, B1 => n14160, B2 => 
                           n14167, ZN => n4225);
   U2052 : OAI22_X1 port map( A1 => n14122, A2 => n14120, B1 => n14123, B2 => 
                           n14121, ZN => n4142);
   U2053 : OAI22_X1 port map( A1 => n14098, A2 => n14099, B1 => n14100, B2 => 
                           n14101, ZN => n4114);
   U2054 : NOR2_X1 port map( A1 => n14259, A2 => N275, ZN => n14250);
   U2055 : AOI22_X1 port map( A1 => n14140, A2 => n14141, B1 => n14105, B2 => 
                           n14086, ZN => n4168);
   U2056 : INV_X1 port map( A => n14142, ZN => n14141);
   U2057 : AOI22_X1 port map( A1 => n14140, A2 => n14171, B1 => n14105, B2 => 
                           n14158, ZN => n4200);
   U2058 : INV_X1 port map( A => n14101, ZN => n14171);
   U2059 : NOR2_X1 port map( A1 => n14257, A2 => N274, ZN => n14067);
   U2060 : NOR2_X1 port map( A1 => n14263, A2 => N273, ZN => n14253);
   U2061 : NOR2_X1 port map( A1 => n14262, A2 => N273, ZN => n14254);
   U2062 : OAI21_X1 port map( B1 => n14005, B2 => n14006, A => n18039, ZN => 
                           n14000);
   U2063 : OAI221_X1 port map( B1 => n14220, B2 => n12413, C1 => n14058, C2 => 
                           n12415, A => n18036, ZN => n4273);
   U2064 : OAI221_X1 port map( B1 => n14217, B2 => n12413, C1 => n12415, C2 => 
                           n14228, A => n18035, ZN => n4270);
   U2065 : OAI221_X1 port map( B1 => n14213, B2 => n12413, C1 => n12415, C2 => 
                           n14226, A => n18035, ZN => n4267);
   U2066 : OAI221_X1 port map( B1 => n12412, B2 => n12413, C1 => n12414, C2 => 
                           n12415, A => n18035, ZN => n10511);
   U2067 : OAI221_X1 port map( B1 => n14214, B2 => n14220, C1 => n12415, C2 => 
                           n14221, A => n18035, ZN => n4259);
   U2068 : OAI221_X1 port map( B1 => n14214, B2 => n12412, C1 => n12415, C2 => 
                           n14222, A => n18035, ZN => n4262);
   U2069 : OAI221_X1 port map( B1 => n14214, B2 => n14217, C1 => n12415, C2 => 
                           n14218, A => n18035, ZN => n4256);
   U2070 : OAI221_X1 port map( B1 => n14213, B2 => n14214, C1 => n12415, C2 => 
                           n14215, A => n18035, ZN => n4251);
   U2071 : NOR2_X1 port map( A1 => N275, A2 => N274, ZN => n14260);
   U2072 : NAND4_X1 port map( A1 => N9922, A2 => N9924, A3 => n14174, A4 => 
                           n14020, ZN => n14099);
   U2073 : NOR2_X1 port map( A1 => N9641, A2 => N9909, ZN => n14133);
   U2074 : INV_X1 port map( A => N9925, ZN => n14205);
   U2075 : AOI22_X1 port map( A1 => n14170, A2 => n14180, B1 => n14176, B2 => 
                           n14092, ZN => n4209);
   U2076 : AOI22_X1 port map( A1 => n14204, A2 => n14170, B1 => n14197, B2 => 
                           n14092, ZN => n4237);
   U2077 : NAND2_X1 port map( A1 => N9925, A2 => n14138, ZN => n14134);
   U2078 : AOI21_X1 port map( B1 => n14105, B2 => n14088, A => n14200, ZN => 
                           n4228);
   U2079 : AND3_X1 port map( A1 => n14147, A2 => n14140, A3 => n14179, ZN => 
                           n14200);
   U2080 : AND3_X1 port map( A1 => N46302, A2 => n13962, A3 => N46303, ZN => 
                           n13957);
   U2081 : AOI21_X1 port map( B1 => n14103, B2 => n14105, A => n14199, ZN => 
                           n4230);
   U2082 : AND3_X1 port map( A1 => n14194, A2 => n14140, A3 => n14147, ZN => 
                           n14199);
   U2083 : AND3_X1 port map( A1 => n12481, A2 => n12499, A3 => N45789, ZN => 
                           n12463);
   U2084 : NAND2_X1 port map( A1 => n13998, A2 => n13997, ZN => n14007);
   U2085 : NAND2_X1 port map( A1 => n14091, A2 => N9925, ZN => n14118);
   U2086 : NAND2_X1 port map( A1 => n14176, A2 => N9925, ZN => n14167);
   U2087 : NAND2_X1 port map( A1 => n14151, A2 => N9925, ZN => n14121);
   U2088 : NOR3_X1 port map( A1 => n16414, A2 => n13981, A3 => n13983, ZN => 
                           n13987);
   U2089 : NOR3_X1 port map( A1 => n16666, A2 => n12500, A3 => n12502, ZN => 
                           n12506);
   U2090 : AOI21_X1 port map( B1 => n14085, B2 => n14104, A => n14127, ZN => 
                           n4159);
   U2091 : AND3_X1 port map( A1 => n14128, A2 => n14129, A3 => n14130, ZN => 
                           n14127);
   U2092 : AOI21_X1 port map( B1 => n14085, B2 => n14094, A => n14132, ZN => 
                           n4157);
   U2093 : AND3_X1 port map( A1 => n14128, A2 => n14133, A3 => n14130, ZN => 
                           n14132);
   U2094 : AOI21_X1 port map( B1 => n14176, B2 => n14152, A => n14177, ZN => 
                           n4211);
   U2095 : AND3_X1 port map( A1 => n14178, A2 => n14179, A3 => n14180, ZN => 
                           n14177);
   U2096 : AOI21_X1 port map( B1 => n14197, B2 => n14152, A => n14206, ZN => 
                           n4235);
   U2097 : AND3_X1 port map( A1 => n14178, A2 => n14179, A3 => n14204, ZN => 
                           n14206);
   U2098 : AND3_X1 port map( A1 => n13962, A2 => n13980, A3 => N46303, ZN => 
                           n13944);
   U2099 : AND3_X1 port map( A1 => n12481, A2 => n12482, A3 => N45788, ZN => 
                           n12444);
   U2100 : AND3_X1 port map( A1 => N45788, A2 => n12481, A3 => N45789, ZN => 
                           n12474);
   U2101 : INV_X1 port map( A => n14165, ZN => n4191);
   U2102 : OAI22_X1 port map( A1 => n14163, A2 => n14159, B1 => n14164, B2 => 
                           n14160, ZN => n14165);
   U2103 : NOR2_X1 port map( A1 => n14020, A2 => n14178, ZN => n14147);
   U2104 : NOR2_X1 port map( A1 => N9921, A2 => N9923, ZN => n14138);
   U2105 : NAND2_X1 port map( A1 => datain(30), A2 => n18039, ZN => n4058);
   U2106 : NAND2_X1 port map( A1 => datain(31), A2 => n18039, ZN => n10510);
   U2107 : NAND2_X1 port map( A1 => datain(24), A2 => n18038, ZN => n5040);
   U2108 : NAND2_X1 port map( A1 => datain(26), A2 => n18038, ZN => n4791);
   U2109 : NAND2_X1 port map( A1 => datain(28), A2 => n18038, ZN => n4533);
   U2110 : NAND2_X1 port map( A1 => datain(7), A2 => n18033, ZN => n7537);
   U2111 : NAND2_X1 port map( A1 => datain(8), A2 => n18037, ZN => n7428);
   U2112 : NAND2_X1 port map( A1 => datain(9), A2 => n18034, ZN => n7319);
   U2113 : NAND2_X1 port map( A1 => datain(10), A2 => n18033, ZN => n7205);
   U2114 : NAND2_X1 port map( A1 => datain(11), A2 => n18034, ZN => n7096);
   U2115 : NAND2_X1 port map( A1 => datain(12), A2 => n18033, ZN => n6987);
   U2116 : NAND2_X1 port map( A1 => datain(13), A2 => n18037, ZN => n6878);
   U2117 : NAND2_X1 port map( A1 => datain(14), A2 => n18034, ZN => n6769);
   U2118 : NAND2_X1 port map( A1 => datain(15), A2 => n18033, ZN => n6635);
   U2119 : NAND2_X1 port map( A1 => datain(16), A2 => n18037, ZN => n6448);
   U2120 : NAND2_X1 port map( A1 => datain(17), A2 => n18037, ZN => n6261);
   U2121 : NAND2_X1 port map( A1 => datain(18), A2 => n18038, ZN => n6076);
   U2122 : NAND2_X1 port map( A1 => datain(19), A2 => n18037, ZN => n5889);
   U2123 : NAND2_X1 port map( A1 => datain(20), A2 => n18034, ZN => n5717);
   U2124 : NAND2_X1 port map( A1 => datain(21), A2 => n18033, ZN => n5530);
   U2125 : NAND2_X1 port map( A1 => datain(22), A2 => n18034, ZN => n5343);
   U2126 : NAND2_X1 port map( A1 => datain(23), A2 => n18038, ZN => n5157);
   U2127 : NAND2_X1 port map( A1 => datain(25), A2 => n18037, ZN => n4924);
   U2128 : NAND2_X1 port map( A1 => datain(27), A2 => n18034, ZN => n4664);
   U2129 : NAND2_X1 port map( A1 => datain(29), A2 => n18038, ZN => n4278);
   U2130 : AND3_X1 port map( A1 => n13962, A2 => n13963, A3 => N46302, ZN => 
                           n13921);
   U2131 : OAI221_X1 port map( B1 => n17836, B2 => n14296, C1 => n17854, C2 => 
                           n16461, A => n18034, ZN => n8030);
   U2132 : OAI221_X1 port map( B1 => n17858, B2 => n14997, C1 => n17876, C2 => 
                           n16461, A => n18034, ZN => n8031);
   U2133 : OAI221_X1 port map( B1 => n17880, B2 => n15361, C1 => n17898, C2 => 
                           n16461, A => n18034, ZN => n8032);
   U2134 : OAI221_X1 port map( B1 => n17902, B2 => n14635, C1 => n17920, C2 => 
                           n16461, A => n18034, ZN => n8033);
   U2135 : OAI221_X1 port map( B1 => n17923, B2 => n15353, C1 => n17941, C2 => 
                           n16461, A => n18034, ZN => n8034);
   U2136 : OAI221_X1 port map( B1 => n17944, B2 => n14863, C1 => n17962, C2 => 
                           n16461, A => n18034, ZN => n8035);
   U2137 : OAI221_X1 port map( B1 => n17965, B2 => n15240, C1 => n17983, C2 => 
                           n16461, A => n18034, ZN => n8036);
   U2138 : OAI221_X1 port map( B1 => n17836, B2 => n14297, C1 => n17854, C2 => 
                           n16714, A => n18036, ZN => n8158);
   U2139 : OAI221_X1 port map( B1 => n17858, B2 => n14998, C1 => n17875, C2 => 
                           n16714, A => n18036, ZN => n8159);
   U2140 : OAI221_X1 port map( B1 => n17880, B2 => n15362, C1 => n17897, C2 => 
                           n16714, A => n18036, ZN => n8160);
   U2141 : OAI221_X1 port map( B1 => n17902, B2 => n14636, C1 => n17920, C2 => 
                           n16714, A => n18036, ZN => n8161);
   U2142 : OAI221_X1 port map( B1 => n17923, B2 => n15354, C1 => n17940, C2 => 
                           n16714, A => n18037, ZN => n8162);
   U2143 : OAI221_X1 port map( B1 => n17944, B2 => n14864, C1 => n17962, C2 => 
                           n16714, A => n18033, ZN => n8163);
   U2144 : OAI221_X1 port map( B1 => n17965, B2 => n15241, C1 => n17983, C2 => 
                           n16714, A => n18034, ZN => n8164);
   U2145 : OAI221_X1 port map( B1 => n17836, B2 => n14298, C1 => n17853, C2 => 
                           n16723, A => n18037, ZN => n8230);
   U2146 : OAI221_X1 port map( B1 => n17858, B2 => n14999, C1 => n17876, C2 => 
                           n16723, A => n18034, ZN => n8231);
   U2147 : OAI221_X1 port map( B1 => n17880, B2 => n15364, C1 => n17898, C2 => 
                           n16723, A => n18037, ZN => n8232);
   U2148 : OAI221_X1 port map( B1 => n17902, B2 => n14637, C1 => n17919, C2 => 
                           n16723, A => n18038, ZN => n8233);
   U2149 : OAI221_X1 port map( B1 => n17923, B2 => n15355, C1 => n17941, C2 => 
                           n16723, A => n18037, ZN => n8234);
   U2150 : OAI221_X1 port map( B1 => n17944, B2 => n14865, C1 => n17961, C2 => 
                           n16723, A => n18038, ZN => n8235);
   U2151 : OAI221_X1 port map( B1 => n17965, B2 => n15242, C1 => n17982, C2 => 
                           n16723, A => n18034, ZN => n8236);
   U2152 : OAI221_X1 port map( B1 => n17170, B2 => n12016, C1 => n17179, C2 => 
                           n16460, A => n18033, ZN => n8050);
   U2153 : OAI221_X1 port map( B1 => n17182, B2 => n12340, C1 => n17190, C2 => 
                           n16460, A => n18033, ZN => n8051);
   U2154 : OAI221_X1 port map( B1 => n17192, B2 => n14282, C1 => n17200, C2 => 
                           n16460, A => n18033, ZN => n8052);
   U2155 : OAI221_X1 port map( B1 => n16944, B2 => n11905, C1 => n16953, C2 => 
                           n16461, A => n18034, ZN => n8039);
   U2156 : OAI221_X1 port map( B1 => n16956, B2 => n14641, C1 => n16964, C2 => 
                           n16460, A => n18033, ZN => n8040);
   U2157 : OAI221_X1 port map( B1 => n16966, B2 => n15356, C1 => n16974, C2 => 
                           n16460, A => n18033, ZN => n8041);
   U2158 : OAI221_X1 port map( B1 => n16976, B2 => n14861, C1 => n16984, C2 => 
                           n16460, A => n18033, ZN => n8042);
   U2159 : OAI221_X1 port map( B1 => n16999, B2 => n14292, C1 => n17007, C2 => 
                           n16460, A => n18033, ZN => n8044);
   U2160 : OAI221_X1 port map( B1 => n17137, B2 => n14638, C1 => n17145, C2 => 
                           n16460, A => n18033, ZN => n8047);
   U2161 : OAI221_X1 port map( B1 => n17160, B2 => n14989, C1 => n17168, C2 => 
                           n16460, A => n18033, ZN => n8049);
   U2162 : OAI221_X1 port map( B1 => n16877, B2 => n14866, C1 => n16885, C2 => 
                           n16713, A => n18037, ZN => n8169);
   U2163 : OAI221_X1 port map( B1 => n16887, B2 => n15351, C1 => n16895, C2 => 
                           n16713, A => n18038, ZN => n8170);
   U2164 : OAI221_X1 port map( B1 => n16910, B2 => n14294, C1 => n16918, C2 => 
                           n16713, A => n18034, ZN => n8172);
   U2165 : OAI221_X1 port map( B1 => n4382, B2 => n14639, C1 => n17145, C2 => 
                           n16713, A => n18038, ZN => n8175);
   U2166 : OAI221_X1 port map( B1 => n4376, B2 => n14990, C1 => n17168, C2 => 
                           n16713, A => n18033, ZN => n8177);
   U2167 : OAI221_X1 port map( B1 => n4373, B2 => n12017, C1 => n17179, C2 => 
                           n16713, A => n18037, ZN => n8178);
   U2168 : OAI221_X1 port map( B1 => n4370, B2 => n12341, C1 => n17190, C2 => 
                           n16713, A => n18037, ZN => n8179);
   U2169 : OAI221_X1 port map( B1 => n4367, B2 => n14283, C1 => n17200, C2 => 
                           n16713, A => n18037, ZN => n8180);
   U2170 : OAI221_X1 port map( B1 => n16877, B2 => n14867, C1 => n16885, C2 => 
                           n16722, A => n18038, ZN => n8241);
   U2171 : OAI221_X1 port map( B1 => n16887, B2 => n15352, C1 => n16895, C2 => 
                           n16722, A => n18037, ZN => n8242);
   U2172 : OAI221_X1 port map( B1 => n16910, B2 => n14295, C1 => n16918, C2 => 
                           n16722, A => n18038, ZN => n8244);
   U2173 : OAI221_X1 port map( B1 => n16944, B2 => n11906, C1 => n16953, C2 => 
                           n16722, A => n18033, ZN => n8247);
   U2174 : OAI221_X1 port map( B1 => n16956, B2 => n14642, C1 => n16964, C2 => 
                           n16722, A => n18038, ZN => n8248);
   U2175 : OAI221_X1 port map( B1 => n16966, B2 => n15357, C1 => n16974, C2 => 
                           n16722, A => n18037, ZN => n8249);
   U2176 : OAI221_X1 port map( B1 => n4429, B2 => n14862, C1 => n16984, C2 => 
                           n16722, A => n18038, ZN => n8250);
   U2177 : OAI221_X1 port map( B1 => n16999, B2 => n14293, C1 => n17007, C2 => 
                           n16722, A => n18034, ZN => n8252);
   U2178 : OAI22_X1 port map( A1 => n16681, A2 => n14960, B1 => n16678, B2 => 
                           n14284, ZN => n12419);
   U2179 : OAI22_X1 port map( A1 => n16681, A2 => n14961, B1 => n16678, B2 => 
                           n14285, ZN => n12262);
   U2180 : OAI22_X1 port map( A1 => n16681, A2 => n14962, B1 => n16678, B2 => 
                           n14286, ZN => n12109);
   U2181 : OAI22_X1 port map( A1 => n16681, A2 => n14980, B1 => n16678, B2 => 
                           n14287, ZN => n11956);
   U2182 : OAI22_X1 port map( A1 => n14051, A2 => n16679, B1 => n16678, B2 => 
                           n14856, ZN => n10518);
   U2183 : OAI22_X1 port map( A1 => n17729, A2 => n15620, B1 => n17726, B2 => 
                           n12332, ZN => n5295);
   U2184 : OAI22_X1 port map( A1 => n17717, A2 => n15631, B1 => n17714, B2 => 
                           n11867, ZN => n5303);
   U2185 : OAI22_X1 port map( A1 => n17729, A2 => n15621, B1 => n17726, B2 => 
                           n12333, ZN => n5129);
   U2186 : OAI22_X1 port map( A1 => n17717, A2 => n15632, B1 => n17714, B2 => 
                           n11869, ZN => n5134);
   U2187 : OAI22_X1 port map( A1 => n17729, A2 => n15622, B1 => n17726, B2 => 
                           n12334, ZN => n5013);
   U2188 : OAI22_X1 port map( A1 => n17717, A2 => n15633, B1 => n17714, B2 => 
                           n11870, ZN => n5020);
   U2189 : OAI22_X1 port map( A1 => n17729, A2 => n15623, B1 => n17726, B2 => 
                           n12335, ZN => n4891);
   U2190 : OAI22_X1 port map( A1 => n17717, A2 => n15634, B1 => n17714, B2 => 
                           n11871, ZN => n4900);
   U2191 : OAI22_X1 port map( A1 => n17729, A2 => n15624, B1 => n17726, B2 => 
                           n12336, ZN => n4764);
   U2192 : OAI22_X1 port map( A1 => n17717, A2 => n15635, B1 => n17714, B2 => 
                           n11872, ZN => n4771);
   U2193 : OAI22_X1 port map( A1 => n17729, A2 => n15625, B1 => n17726, B2 => 
                           n12337, ZN => n4633);
   U2194 : OAI22_X1 port map( A1 => n17717, A2 => n15636, B1 => n17714, B2 => 
                           n11873, ZN => n4638);
   U2195 : OAI22_X1 port map( A1 => n17729, A2 => n15614, B1 => n17726, B2 => 
                           n12339, ZN => n4506);
   U2196 : OAI22_X1 port map( A1 => n17717, A2 => n15615, B1 => n17714, B2 => 
                           n11861, ZN => n4511);
   U2197 : OAI22_X1 port map( A1 => n17729, A2 => n15278, B1 => n17726, B2 => 
                           n12163, ZN => n4172);
   U2198 : OAI22_X1 port map( A1 => n17717, A2 => n15279, B1 => n17714, B2 => 
                           n11498, ZN => n4183);
   U2199 : OAI22_X1 port map( A1 => n16333, A2 => n15060, B1 => n16330, B2 => 
                           n12165, ZN => n12913);
   U2200 : OAI22_X1 port map( A1 => n16321, A2 => n15176, B1 => n16318, B2 => 
                           n14403, ZN => n12914);
   U2201 : OAI22_X1 port map( A1 => n16345, A2 => n12333, B1 => n16342, B2 => 
                           n11869, ZN => n12912);
   U2202 : OAI22_X1 port map( A1 => n16393, A2 => n14825, B1 => n16390, B2 => 
                           n11875, ZN => n12904);
   U2203 : OAI22_X1 port map( A1 => n16381, A2 => n15396, B1 => n16378, B2 => 
                           n14414, ZN => n12905);
   U2204 : OAI22_X1 port map( A1 => n16333, A2 => n15061, B1 => n16330, B2 => 
                           n12166, ZN => n12871);
   U2205 : OAI22_X1 port map( A1 => n16321, A2 => n15177, B1 => n16318, B2 => 
                           n14404, ZN => n12872);
   U2206 : OAI22_X1 port map( A1 => n16345, A2 => n12334, B1 => n16342, B2 => 
                           n11870, ZN => n12870);
   U2207 : OAI22_X1 port map( A1 => n16393, A2 => n14826, B1 => n16390, B2 => 
                           n11876, ZN => n12862);
   U2208 : OAI22_X1 port map( A1 => n16381, A2 => n15397, B1 => n16378, B2 => 
                           n14415, ZN => n12863);
   U2209 : OAI22_X1 port map( A1 => n16333, A2 => n15062, B1 => n16330, B2 => 
                           n12167, ZN => n12829);
   U2210 : OAI22_X1 port map( A1 => n16321, A2 => n15178, B1 => n16318, B2 => 
                           n14405, ZN => n12830);
   U2211 : OAI22_X1 port map( A1 => n16345, A2 => n12335, B1 => n16342, B2 => 
                           n11871, ZN => n12828);
   U2212 : OAI22_X1 port map( A1 => n16393, A2 => n14827, B1 => n16390, B2 => 
                           n11877, ZN => n12820);
   U2213 : OAI22_X1 port map( A1 => n16381, A2 => n15398, B1 => n16378, B2 => 
                           n14416, ZN => n12821);
   U2214 : OAI22_X1 port map( A1 => n16333, A2 => n15063, B1 => n16330, B2 => 
                           n12168, ZN => n12787);
   U2215 : OAI22_X1 port map( A1 => n16321, A2 => n15179, B1 => n16318, B2 => 
                           n14406, ZN => n12788);
   U2216 : OAI22_X1 port map( A1 => n16345, A2 => n12336, B1 => n16342, B2 => 
                           n11872, ZN => n12786);
   U2217 : OAI22_X1 port map( A1 => n16393, A2 => n14828, B1 => n16390, B2 => 
                           n11878, ZN => n12778);
   U2218 : OAI22_X1 port map( A1 => n16381, A2 => n15399, B1 => n16378, B2 => 
                           n14417, ZN => n12779);
   U2219 : OAI22_X1 port map( A1 => n16333, A2 => n15064, B1 => n16330, B2 => 
                           n12169, ZN => n12745);
   U2220 : OAI22_X1 port map( A1 => n16321, A2 => n15180, B1 => n16318, B2 => 
                           n14407, ZN => n12746);
   U2221 : OAI22_X1 port map( A1 => n16345, A2 => n12337, B1 => n16342, B2 => 
                           n11873, ZN => n12744);
   U2222 : OAI22_X1 port map( A1 => n16393, A2 => n14829, B1 => n16390, B2 => 
                           n11879, ZN => n12736);
   U2223 : OAI22_X1 port map( A1 => n16381, A2 => n15400, B1 => n16378, B2 => 
                           n14418, ZN => n12737);
   U2224 : OAI22_X1 port map( A1 => n16333, A2 => n15054, B1 => n16330, B2 => 
                           n12170, ZN => n12703);
   U2225 : OAI22_X1 port map( A1 => n16321, A2 => n15169, B1 => n16318, B2 => 
                           n14396, ZN => n12704);
   U2226 : OAI22_X1 port map( A1 => n16345, A2 => n12339, B1 => n16342, B2 => 
                           n11861, ZN => n12702);
   U2227 : OAI22_X1 port map( A1 => n16393, A2 => n14830, B1 => n16390, B2 => 
                           n11880, ZN => n12694);
   U2228 : OAI22_X1 port map( A1 => n16381, A2 => n15390, B1 => n16378, B2 => 
                           n14397, ZN => n12695);
   U2229 : OAI22_X1 port map( A1 => n16333, A2 => n14869, B1 => n16330, B2 => 
                           n12160, ZN => n12660);
   U2230 : OAI22_X1 port map( A1 => n16321, A2 => n14872, B1 => n16318, B2 => 
                           n14056, ZN => n12661);
   U2231 : OAI22_X1 port map( A1 => n16345, A2 => n12163, B1 => n16342, B2 => 
                           n11498, ZN => n12659);
   U2232 : OAI22_X1 port map( A1 => n16393, A2 => n14822, B1 => n16390, B2 => 
                           n11541, ZN => n12650);
   U2233 : OAI22_X1 port map( A1 => n16381, A2 => n15273, B1 => n16378, B2 => 
                           n14057, ZN => n12651);
   U2234 : OAI22_X1 port map( A1 => n16333, A2 => n15041, B1 => n16330, B2 => 
                           n12194, ZN => n12574);
   U2235 : OAI22_X1 port map( A1 => n16321, A2 => n15156, B1 => n16318, B2 => 
                           n14370, ZN => n12579);
   U2236 : OAI22_X1 port map( A1 => n16345, A2 => n12314, B1 => n16342, B2 => 
                           n11845, ZN => n12569);
   U2237 : OAI22_X1 port map( A1 => n16393, A2 => n14853, B1 => n16390, B2 => 
                           n11903, ZN => n12544);
   U2238 : OAI22_X1 port map( A1 => n16381, A2 => n15377, B1 => n16378, B2 => 
                           n14371, ZN => n12549);
   U2239 : OAI22_X1 port map( A1 => n16585, A2 => n15176, B1 => n16582, B2 => 
                           n14403, ZN => n10963);
   U2240 : OAI22_X1 port map( A1 => n16573, A2 => n15060, B1 => n16570, B2 => 
                           n12165, ZN => n10964);
   U2241 : OAI22_X1 port map( A1 => n16597, A2 => n12333, B1 => n16594, B2 => 
                           n11869, ZN => n10962);
   U2242 : OAI22_X1 port map( A1 => n16633, A2 => n14825, B1 => n16630, B2 => 
                           n14414, ZN => n10955);
   U2243 : OAI22_X1 port map( A1 => n16645, A2 => n14599, B1 => n16642, B2 => 
                           n11875, ZN => n10954);
   U2244 : OAI22_X1 port map( A1 => n16585, A2 => n15177, B1 => n16582, B2 => 
                           n14404, ZN => n10920);
   U2245 : OAI22_X1 port map( A1 => n16573, A2 => n15061, B1 => n16570, B2 => 
                           n12166, ZN => n10921);
   U2246 : OAI22_X1 port map( A1 => n16597, A2 => n12334, B1 => n16594, B2 => 
                           n11870, ZN => n10919);
   U2247 : OAI22_X1 port map( A1 => n16633, A2 => n14826, B1 => n16630, B2 => 
                           n14415, ZN => n10912);
   U2248 : OAI22_X1 port map( A1 => n16645, A2 => n14600, B1 => n16642, B2 => 
                           n11876, ZN => n10911);
   U2249 : OAI22_X1 port map( A1 => n16585, A2 => n15178, B1 => n16582, B2 => 
                           n14405, ZN => n10877);
   U2250 : OAI22_X1 port map( A1 => n16573, A2 => n15062, B1 => n16570, B2 => 
                           n12167, ZN => n10878);
   U2251 : OAI22_X1 port map( A1 => n16597, A2 => n12335, B1 => n16594, B2 => 
                           n11871, ZN => n10876);
   U2252 : OAI22_X1 port map( A1 => n16633, A2 => n14827, B1 => n16630, B2 => 
                           n14416, ZN => n10869);
   U2253 : OAI22_X1 port map( A1 => n16645, A2 => n14601, B1 => n16642, B2 => 
                           n11877, ZN => n10868);
   U2254 : OAI22_X1 port map( A1 => n16585, A2 => n15179, B1 => n16582, B2 => 
                           n14406, ZN => n10834);
   U2255 : OAI22_X1 port map( A1 => n16573, A2 => n15063, B1 => n16570, B2 => 
                           n12168, ZN => n10835);
   U2256 : OAI22_X1 port map( A1 => n16597, A2 => n12336, B1 => n16594, B2 => 
                           n11872, ZN => n10833);
   U2257 : OAI22_X1 port map( A1 => n16633, A2 => n14828, B1 => n16630, B2 => 
                           n14417, ZN => n10826);
   U2258 : OAI22_X1 port map( A1 => n16645, A2 => n14602, B1 => n16642, B2 => 
                           n11878, ZN => n10825);
   U2259 : OAI22_X1 port map( A1 => n16585, A2 => n15180, B1 => n16582, B2 => 
                           n14407, ZN => n10791);
   U2260 : OAI22_X1 port map( A1 => n16573, A2 => n15064, B1 => n16570, B2 => 
                           n12169, ZN => n10792);
   U2261 : OAI22_X1 port map( A1 => n16597, A2 => n12337, B1 => n16594, B2 => 
                           n11873, ZN => n10790);
   U2262 : OAI22_X1 port map( A1 => n16633, A2 => n14829, B1 => n16630, B2 => 
                           n14418, ZN => n10783);
   U2263 : OAI22_X1 port map( A1 => n16645, A2 => n14603, B1 => n16642, B2 => 
                           n11879, ZN => n10782);
   U2264 : OAI22_X1 port map( A1 => n16585, A2 => n15169, B1 => n16582, B2 => 
                           n14396, ZN => n10748);
   U2265 : OAI22_X1 port map( A1 => n16573, A2 => n15054, B1 => n16570, B2 => 
                           n12170, ZN => n10749);
   U2266 : OAI22_X1 port map( A1 => n16597, A2 => n12339, B1 => n16594, B2 => 
                           n11861, ZN => n10747);
   U2267 : OAI22_X1 port map( A1 => n16633, A2 => n14830, B1 => n16630, B2 => 
                           n14397, ZN => n10740);
   U2268 : OAI22_X1 port map( A1 => n16645, A2 => n14604, B1 => n16642, B2 => 
                           n11880, ZN => n10739);
   U2269 : OAI22_X1 port map( A1 => n16585, A2 => n14872, B1 => n16582, B2 => 
                           n14056, ZN => n10695);
   U2270 : OAI22_X1 port map( A1 => n16573, A2 => n14869, B1 => n16570, B2 => 
                           n12160, ZN => n10698);
   U2271 : OAI22_X1 port map( A1 => n16597, A2 => n12163, B1 => n16594, B2 => 
                           n11498, ZN => n10694);
   U2272 : OAI22_X1 port map( A1 => n16633, A2 => n14822, B1 => n16630, B2 => 
                           n14057, ZN => n10683);
   U2273 : OAI22_X1 port map( A1 => n16645, A2 => n14299, B1 => n16642, B2 => 
                           n11541, ZN => n10682);
   U2274 : OAI22_X1 port map( A1 => n16585, A2 => n15156, B1 => n16582, B2 => 
                           n14370, ZN => n10584);
   U2275 : OAI22_X1 port map( A1 => n16573, A2 => n15041, B1 => n16570, B2 => 
                           n12194, ZN => n10591);
   U2276 : OAI22_X1 port map( A1 => n16597, A2 => n12314, B1 => n16594, B2 => 
                           n11845, ZN => n10577);
   U2277 : OAI22_X1 port map( A1 => n16633, A2 => n14853, B1 => n16630, B2 => 
                           n14371, ZN => n10551);
   U2278 : OAI22_X1 port map( A1 => n16645, A2 => n14627, B1 => n16642, B2 => 
                           n11903, ZN => n10544);
   U2279 : OAI22_X1 port map( A1 => n17765, A2 => n15420, B1 => n17762, B2 => 
                           n14505, ZN => n5292);
   U2280 : OAI22_X1 port map( A1 => n17753, A2 => n14049, B1 => n17750, B2 => 
                           n12040, ZN => n5293);
   U2281 : OAI22_X1 port map( A1 => n17681, A2 => n14568, B1 => n17678, B2 => 
                           n12015, ZN => n5307);
   U2282 : OAI22_X1 port map( A1 => n17705, A2 => n15654, B1 => n17702, B2 => 
                           n14663, ZN => n5304);
   U2283 : OAI22_X1 port map( A1 => n17765, A2 => n15421, B1 => n17762, B2 => 
                           n14471, ZN => n5124);
   U2284 : OAI22_X1 port map( A1 => n17753, A2 => n12349, B1 => n17750, B2 => 
                           n12041, ZN => n5125);
   U2285 : OAI22_X1 port map( A1 => n17681, A2 => n14540, B1 => n17678, B2 => 
                           n11907, ZN => n5137);
   U2286 : OAI22_X1 port map( A1 => n17705, A2 => n15655, B1 => n17702, B2 => 
                           n14664, ZN => n5135);
   U2287 : OAI22_X1 port map( A1 => n17765, A2 => n15422, B1 => n17762, B2 => 
                           n14472, ZN => n5010);
   U2288 : OAI22_X1 port map( A1 => n17753, A2 => n12350, B1 => n17750, B2 => 
                           n12042, ZN => n5011);
   U2289 : OAI22_X1 port map( A1 => n17681, A2 => n14541, B1 => n17678, B2 => 
                           n11945, ZN => n5023);
   U2290 : OAI22_X1 port map( A1 => n17705, A2 => n15656, B1 => n17702, B2 => 
                           n14665, ZN => n5021);
   U2291 : OAI22_X1 port map( A1 => n17765, A2 => n15423, B1 => n17762, B2 => 
                           n14473, ZN => n4888);
   U2292 : OAI22_X1 port map( A1 => n17753, A2 => n12351, B1 => n17750, B2 => 
                           n12043, ZN => n4889);
   U2293 : OAI22_X1 port map( A1 => n17681, A2 => n14542, B1 => n17678, B2 => 
                           n11946, ZN => n4903);
   U2294 : OAI22_X1 port map( A1 => n17705, A2 => n15657, B1 => n17702, B2 => 
                           n14666, ZN => n4901);
   U2295 : OAI22_X1 port map( A1 => n17765, A2 => n15424, B1 => n17762, B2 => 
                           n14474, ZN => n4761);
   U2296 : OAI22_X1 port map( A1 => n17753, A2 => n12352, B1 => n17750, B2 => 
                           n12044, ZN => n4762);
   U2297 : OAI22_X1 port map( A1 => n17681, A2 => n14543, B1 => n17678, B2 => 
                           n11947, ZN => n4774);
   U2298 : OAI22_X1 port map( A1 => n17705, A2 => n15658, B1 => n17702, B2 => 
                           n14667, ZN => n4772);
   U2299 : OAI22_X1 port map( A1 => n17765, A2 => n15425, B1 => n17762, B2 => 
                           n14475, ZN => n4630);
   U2300 : OAI22_X1 port map( A1 => n17753, A2 => n12353, B1 => n17750, B2 => 
                           n12045, ZN => n4631);
   U2301 : OAI22_X1 port map( A1 => n17681, A2 => n14544, B1 => n17678, B2 => 
                           n11948, ZN => n4641);
   U2302 : OAI22_X1 port map( A1 => n17705, A2 => n15659, B1 => n17702, B2 => 
                           n14668, ZN => n4639);
   U2303 : OAI22_X1 port map( A1 => n17765, A2 => n15426, B1 => n17762, B2 => 
                           n14476, ZN => n4501);
   U2304 : OAI22_X1 port map( A1 => n17753, A2 => n12354, B1 => n17750, B2 => 
                           n12046, ZN => n4502);
   U2305 : OAI22_X1 port map( A1 => n17681, A2 => n14545, B1 => n17678, B2 => 
                           n11949, ZN => n4514);
   U2306 : OAI22_X1 port map( A1 => n17705, A2 => n15660, B1 => n17702, B2 => 
                           n14644, ZN => n4512);
   U2307 : OAI22_X1 port map( A1 => n17765, A2 => n15272, B1 => n17762, B2 => 
                           n14065, ZN => n4145);
   U2308 : OAI22_X1 port map( A1 => n17753, A2 => n12197, B1 => n17750, B2 => 
                           n11904, ZN => n4156);
   U2309 : OAI22_X1 port map( A1 => n17681, A2 => n14279, B1 => n17678, B2 => 
                           n11670, ZN => n4208);
   U2310 : OAI22_X1 port map( A1 => n17705, A2 => n15316, B1 => n17702, B2 => 
                           n14633, ZN => n4190);
   U2311 : NOR2_X1 port map( A1 => n14209, A2 => N9921, ZN => n14202);
   U2312 : OAI221_X1 port map( B1 => n17322, B2 => n15284, C1 => n17321, C2 => 
                           n16462, A => n18035, ZN => n8014);
   U2313 : OAI221_X1 port map( B1 => n17335, B2 => n11627, C1 => n17334, C2 => 
                           n16462, A => n18035, ZN => n8015);
   U2314 : OAI221_X1 port map( B1 => n17348, B2 => n14994, C1 => n17347, C2 => 
                           n16462, A => n18035, ZN => n8016);
   U2315 : OAI221_X1 port map( B1 => n17361, B2 => n15365, C1 => n17360, C2 => 
                           n16462, A => n18035, ZN => n8017);
   U2316 : OAI221_X1 port map( B1 => n17374, B2 => n14291, C1 => n17373, C2 => 
                           n16462, A => n18035, ZN => n8018);
   U2317 : OAI221_X1 port map( B1 => n17387, B2 => n14640, C1 => n17386, C2 => 
                           n16461, A => n18034, ZN => n8019);
   U2318 : OAI221_X1 port map( B1 => n17400, B2 => n14288, C1 => n17399, C2 => 
                           n16461, A => n18034, ZN => n8020);
   U2319 : OAI221_X1 port map( B1 => n17413, B2 => n15003, C1 => n17412, C2 => 
                           n16461, A => n18034, ZN => n8021);
   U2320 : OAI221_X1 port map( B1 => n16936, B2 => n14536, C1 => n16935, C2 => 
                           n16461, A => n18034, ZN => n8038);
   U2321 : OAI221_X1 port map( B1 => n17009, B2 => n14995, C1 => n17017, C2 => 
                           n16460, A => n18033, ZN => n8045);
   U2322 : OAI221_X1 port map( B1 => n16693, B2 => n14868, C1 => n16692, C2 => 
                           n10285, A => n18036, ZN => n8059);
   U2323 : OAI221_X1 port map( B1 => n17129, B2 => n15367, C1 => n17128, C2 => 
                           n16460, A => n18033, ZN => n8046);
   U2324 : OAI221_X1 port map( B1 => n17202, B2 => n15001, C1 => n17210, C2 => 
                           n16460, A => n18033, ZN => n8053);
   U2325 : OAI221_X1 port map( B1 => n17231, B2 => n15350, C1 => n17230, C2 => 
                           n16715, A => n18036, ZN => n8135);
   U2326 : OAI221_X1 port map( B1 => n17244, B2 => n12195, C1 => n17243, C2 => 
                           n16715, A => n18036, ZN => n8136);
   U2327 : OAI221_X1 port map( B1 => n17257, B2 => n14823, C1 => n17256, C2 => 
                           n16714, A => n18036, ZN => n8137);
   U2328 : OAI221_X1 port map( B1 => n17283, B2 => n14289, C1 => n17282, C2 => 
                           n16714, A => n18036, ZN => n8139);
   U2329 : OAI221_X1 port map( B1 => n17296, B2 => n14569, C1 => n17295, C2 => 
                           n16714, A => n18036, ZN => n8140);
   U2330 : OAI221_X1 port map( B1 => n17309, B2 => n15366, C1 => n17308, C2 => 
                           n16714, A => n18036, ZN => n8141);
   U2331 : OAI221_X1 port map( B1 => n18005, B2 => n12050, C1 => n18004, C2 => 
                           n16714, A => n18034, ZN => n8166);
   U2332 : OAI221_X1 port map( B1 => n18018, B2 => n14538, C1 => n18017, C2 => 
                           n16713, A => n18033, ZN => n8167);
   U2333 : OAI221_X1 port map( B1 => n16920, B2 => n15359, C1 => n16928, C2 => 
                           n16713, A => n18037, ZN => n8173);
   U2334 : OAI221_X1 port map( B1 => n17129, B2 => n15368, C1 => n17127, C2 => 
                           n16713, A => n18033, ZN => n8174);
   U2335 : OAI221_X1 port map( B1 => n4362, B2 => n15002, C1 => n17210, C2 => 
                           n16713, A => n18038, ZN => n8181);
   U2336 : OAI221_X1 port map( B1 => n17025, B2 => n12162, C1 => n17024, C2 => 
                           n16724, A => n18037, ZN => n8190);
   U2337 : OAI221_X1 port map( B1 => n17038, B2 => n14993, C1 => n17037, C2 => 
                           n16724, A => n18037, ZN => n8191);
   U2338 : OAI221_X1 port map( B1 => n17051, B2 => n14290, C1 => n17050, C2 => 
                           n16724, A => n18037, ZN => n8192);
   U2339 : OAI221_X1 port map( B1 => n17064, B2 => n15000, C1 => n17063, C2 => 
                           n16724, A => n18038, ZN => n8193);
   U2340 : OAI221_X1 port map( B1 => n17077, B2 => n15363, C1 => n17076, C2 => 
                           n16723, A => n18037, ZN => n8194);
   U2341 : OAI221_X1 port map( B1 => n17090, B2 => n15358, C1 => n17089, C2 => 
                           n16723, A => n18033, ZN => n8195);
   U2342 : OAI221_X1 port map( B1 => n17103, B2 => n11584, C1 => n17102, C2 => 
                           n16723, A => n18037, ZN => n8196);
   U2343 : OAI221_X1 port map( B1 => n17116, B2 => n12308, C1 => n17115, C2 => 
                           n16723, A => n18033, ZN => n8197);
   U2344 : OAI221_X1 port map( B1 => n18005, B2 => n12051, C1 => n18003, C2 => 
                           n16723, A => n18038, ZN => n8238);
   U2345 : OAI221_X1 port map( B1 => n18018, B2 => n14539, C1 => n18016, C2 => 
                           n16722, A => n18037, ZN => n8239);
   U2346 : OAI221_X1 port map( B1 => n16920, B2 => n15360, C1 => n16928, C2 => 
                           n16722, A => n18038, ZN => n8245);
   U2347 : OAI221_X1 port map( B1 => n16936, B2 => n14537, C1 => n16934, C2 => 
                           n16722, A => n18038, ZN => n8246);
   U2348 : OAI221_X1 port map( B1 => n4420, B2 => n14996, C1 => n17017, C2 => 
                           n16722, A => n18038, ZN => n8253);
   U2349 : OAI221_X1 port map( B1 => n17578, B2 => n14053, C1 => n17577, C2 => 
                           n10285, A => n18037, ZN => n8257);
   U2350 : OAI22_X1 port map( A1 => n14983, A2 => n16429, B1 => n14273, B2 => 
                           n16426, ZN => n12892);
   U2351 : OAI22_X1 port map( A1 => n14984, A2 => n16429, B1 => n14274, B2 => 
                           n16426, ZN => n12850);
   U2352 : OAI22_X1 port map( A1 => n14985, A2 => n16429, B1 => n14275, B2 => 
                           n16426, ZN => n12808);
   U2353 : OAI22_X1 port map( A1 => n14986, A2 => n16429, B1 => n14276, B2 => 
                           n16426, ZN => n12766);
   U2354 : OAI22_X1 port map( A1 => n14987, A2 => n16429, B1 => n14277, B2 => 
                           n16426, ZN => n12724);
   U2355 : OAI22_X1 port map( A1 => n14988, A2 => n16429, B1 => n14278, B2 => 
                           n16426, ZN => n12682);
   U2356 : OAI22_X1 port map( A1 => n14860, A2 => n16429, B1 => n14052, B2 => 
                           n16426, ZN => n12638);
   U2357 : OAI22_X1 port map( A1 => n14051, A2 => n16429, B1 => n14856, B2 => 
                           n16426, ZN => n12521);
   U2358 : OAI22_X1 port map( A1 => n16681, A2 => n14963, B1 => n14071, B2 => 
                           n16678, ZN => n11803);
   U2359 : OAI22_X1 port map( A1 => n16681, A2 => n14964, B1 => n14212, B2 => 
                           n16678, ZN => n11760);
   U2360 : OAI22_X1 port map( A1 => n16680, A2 => n14868, B1 => n14053, B2 => 
                           n16678, ZN => n11717);
   U2361 : OAI22_X1 port map( A1 => n16331, A2 => n15037, B1 => n16328, B2 => 
                           n12171, ZN => n13945);
   U2362 : OAI22_X1 port map( A1 => n16319, A2 => n15152, B1 => n16316, B2 => 
                           n14359, ZN => n13947);
   U2363 : OAI22_X1 port map( A1 => n16343, A2 => n12309, B1 => n16340, B2 => 
                           n11713, ZN => n13943);
   U2364 : OAI22_X1 port map( A1 => n16391, A2 => n14831, B1 => n16388, B2 => 
                           n11881, ZN => n13924);
   U2365 : OAI22_X1 port map( A1 => n16379, A2 => n15373, B1 => n16376, B2 => 
                           n14362, ZN => n13930);
   U2366 : OAI22_X1 port map( A1 => n16331, A2 => n15035, B1 => n16328, B2 => 
                           n12172, ZN => n13879);
   U2367 : OAI22_X1 port map( A1 => n16319, A2 => n15153, B1 => n16316, B2 => 
                           n14363, ZN => n13880);
   U2368 : OAI22_X1 port map( A1 => n16343, A2 => n12310, B1 => n16340, B2 => 
                           n11756, ZN => n13878);
   U2369 : OAI22_X1 port map( A1 => n16391, A2 => n14832, B1 => n16388, B2 => 
                           n11882, ZN => n13870);
   U2370 : OAI22_X1 port map( A1 => n16379, A2 => n15371, B1 => n16376, B2 => 
                           n14360, ZN => n13871);
   U2371 : OAI22_X1 port map( A1 => n16331, A2 => n15036, B1 => n16328, B2 => 
                           n12173, ZN => n13837);
   U2372 : OAI22_X1 port map( A1 => n16319, A2 => n15151, B1 => n16316, B2 => 
                           n14361, ZN => n13838);
   U2373 : OAI22_X1 port map( A1 => n16343, A2 => n12311, B1 => n16340, B2 => 
                           n11799, ZN => n13836);
   U2374 : OAI22_X1 port map( A1 => n16391, A2 => n14833, B1 => n16388, B2 => 
                           n11883, ZN => n13828);
   U2375 : OAI22_X1 port map( A1 => n16379, A2 => n15372, B1 => n16376, B2 => 
                           n14364, ZN => n13829);
   U2376 : OAI22_X1 port map( A1 => n16331, A2 => n15038, B1 => n16328, B2 => 
                           n12174, ZN => n13795);
   U2377 : OAI22_X1 port map( A1 => n16319, A2 => n15154, B1 => n16316, B2 => 
                           n14365, ZN => n13796);
   U2378 : OAI22_X1 port map( A1 => n16343, A2 => n12312, B1 => n16340, B2 => 
                           n11842, ZN => n13794);
   U2379 : OAI22_X1 port map( A1 => n16391, A2 => n14834, B1 => n16388, B2 => 
                           n11627, ZN => n13786);
   U2380 : OAI22_X1 port map( A1 => n16379, A2 => n15374, B1 => n16376, B2 => 
                           n14366, ZN => n13787);
   U2381 : OAI22_X1 port map( A1 => n16331, A2 => n15039, B1 => n16328, B2 => 
                           n12175, ZN => n13753);
   U2382 : OAI22_X1 port map( A1 => n16319, A2 => n15155, B1 => n16316, B2 => 
                           n14367, ZN => n13754);
   U2383 : OAI22_X1 port map( A1 => n16343, A2 => n12313, B1 => n16340, B2 => 
                           n11844, ZN => n13752);
   U2384 : OAI22_X1 port map( A1 => n16391, A2 => n14823, B1 => n16388, B2 => 
                           n11884, ZN => n13744);
   U2385 : OAI22_X1 port map( A1 => n16379, A2 => n15350, B1 => n16376, B2 => 
                           n14289, ZN => n13745);
   U2386 : OAI22_X1 port map( A1 => n16331, A2 => n14993, B1 => n16328, B2 => 
                           n12162, ZN => n13711);
   U2387 : OAI22_X1 port map( A1 => n16319, A2 => n15000, B1 => n16316, B2 => 
                           n14290, ZN => n13712);
   U2388 : OAI22_X1 port map( A1 => n16343, A2 => n12308, B1 => n16340, B2 => 
                           n11584, ZN => n13710);
   U2389 : OAI22_X1 port map( A1 => n16391, A2 => n14835, B1 => n16388, B2 => 
                           n11885, ZN => n13702);
   U2390 : OAI22_X1 port map( A1 => n16379, A2 => n15375, B1 => n16376, B2 => 
                           n14368, ZN => n13703);
   U2391 : OAI22_X1 port map( A1 => n16331, A2 => n15040, B1 => n16328, B2 => 
                           n12176, ZN => n13669);
   U2392 : OAI22_X1 port map( A1 => n16319, A2 => n15157, B1 => n16316, B2 => 
                           n14369, ZN => n13670);
   U2393 : OAI22_X1 port map( A1 => n16343, A2 => n12315, B1 => n16340, B2 => 
                           n11846, ZN => n13668);
   U2394 : OAI22_X1 port map( A1 => n16391, A2 => n14836, B1 => n16388, B2 => 
                           n11886, ZN => n13660);
   U2395 : OAI22_X1 port map( A1 => n16379, A2 => n15376, B1 => n16376, B2 => 
                           n14372, ZN => n13661);
   U2396 : OAI22_X1 port map( A1 => n16331, A2 => n15042, B1 => n16328, B2 => 
                           n12177, ZN => n13627);
   U2397 : OAI22_X1 port map( A1 => n16319, A2 => n15158, B1 => n16316, B2 => 
                           n14373, ZN => n13628);
   U2398 : OAI22_X1 port map( A1 => n16343, A2 => n12316, B1 => n16340, B2 => 
                           n11847, ZN => n13626);
   U2399 : OAI22_X1 port map( A1 => n16391, A2 => n14837, B1 => n16388, B2 => 
                           n11887, ZN => n13618);
   U2400 : OAI22_X1 port map( A1 => n16379, A2 => n15378, B1 => n16376, B2 => 
                           n14374, ZN => n13619);
   U2401 : OAI22_X1 port map( A1 => n16331, A2 => n15043, B1 => n16328, B2 => 
                           n12178, ZN => n13585);
   U2402 : OAI22_X1 port map( A1 => n16319, A2 => n15159, B1 => n16316, B2 => 
                           n14375, ZN => n13586);
   U2403 : OAI22_X1 port map( A1 => n16343, A2 => n12317, B1 => n16340, B2 => 
                           n11849, ZN => n13584);
   U2404 : OAI22_X1 port map( A1 => n16391, A2 => n14838, B1 => n16388, B2 => 
                           n11888, ZN => n13576);
   U2405 : OAI22_X1 port map( A1 => n16379, A2 => n15379, B1 => n16376, B2 => 
                           n14376, ZN => n13577);
   U2406 : OAI22_X1 port map( A1 => n16331, A2 => n15044, B1 => n16328, B2 => 
                           n12179, ZN => n13543);
   U2407 : OAI22_X1 port map( A1 => n16319, A2 => n15160, B1 => n16316, B2 => 
                           n14377, ZN => n13544);
   U2408 : OAI22_X1 port map( A1 => n16343, A2 => n12318, B1 => n16340, B2 => 
                           n11850, ZN => n13542);
   U2409 : OAI22_X1 port map( A1 => n16391, A2 => n14839, B1 => n16388, B2 => 
                           n11889, ZN => n13534);
   U2410 : OAI22_X1 port map( A1 => n16379, A2 => n15380, B1 => n16376, B2 => 
                           n14378, ZN => n13535);
   U2411 : OAI22_X1 port map( A1 => n16331, A2 => n15045, B1 => n16328, B2 => 
                           n12180, ZN => n13501);
   U2412 : OAI22_X1 port map( A1 => n16319, A2 => n15161, B1 => n16316, B2 => 
                           n14379, ZN => n13502);
   U2413 : OAI22_X1 port map( A1 => n16343, A2 => n12319, B1 => n16340, B2 => 
                           n11851, ZN => n13500);
   U2414 : OAI22_X1 port map( A1 => n16391, A2 => n14840, B1 => n16388, B2 => 
                           n11890, ZN => n13492);
   U2415 : OAI22_X1 port map( A1 => n16379, A2 => n15381, B1 => n16376, B2 => 
                           n14380, ZN => n13493);
   U2416 : OAI22_X1 port map( A1 => n16331, A2 => n15046, B1 => n16328, B2 => 
                           n12181, ZN => n13459);
   U2417 : OAI22_X1 port map( A1 => n16319, A2 => n15162, B1 => n16316, B2 => 
                           n14381, ZN => n13460);
   U2418 : OAI22_X1 port map( A1 => n16343, A2 => n12320, B1 => n16340, B2 => 
                           n11852, ZN => n13458);
   U2419 : OAI22_X1 port map( A1 => n16391, A2 => n14841, B1 => n16388, B2 => 
                           n11891, ZN => n13450);
   U2420 : OAI22_X1 port map( A1 => n16379, A2 => n15382, B1 => n16376, B2 => 
                           n14382, ZN => n13451);
   U2421 : OAI22_X1 port map( A1 => n16332, A2 => n15047, B1 => n16329, B2 => 
                           n12182, ZN => n13417);
   U2422 : OAI22_X1 port map( A1 => n16320, A2 => n15163, B1 => n16317, B2 => 
                           n14383, ZN => n13418);
   U2423 : OAI22_X1 port map( A1 => n16344, A2 => n12321, B1 => n16341, B2 => 
                           n11854, ZN => n13416);
   U2424 : OAI22_X1 port map( A1 => n16392, A2 => n14842, B1 => n16389, B2 => 
                           n11892, ZN => n13408);
   U2425 : OAI22_X1 port map( A1 => n16380, A2 => n15383, B1 => n16377, B2 => 
                           n14384, ZN => n13409);
   U2426 : OAI22_X1 port map( A1 => n16332, A2 => n15048, B1 => n16329, B2 => 
                           n12183, ZN => n13375);
   U2427 : OAI22_X1 port map( A1 => n16320, A2 => n15164, B1 => n16317, B2 => 
                           n14385, ZN => n13376);
   U2428 : OAI22_X1 port map( A1 => n16344, A2 => n12322, B1 => n16341, B2 => 
                           n11855, ZN => n13374);
   U2429 : OAI22_X1 port map( A1 => n16392, A2 => n14843, B1 => n16389, B2 => 
                           n11893, ZN => n13366);
   U2430 : OAI22_X1 port map( A1 => n16380, A2 => n15384, B1 => n16377, B2 => 
                           n14386, ZN => n13367);
   U2431 : OAI22_X1 port map( A1 => n16332, A2 => n15049, B1 => n16329, B2 => 
                           n12185, ZN => n13333);
   U2432 : OAI22_X1 port map( A1 => n16320, A2 => n15165, B1 => n16317, B2 => 
                           n14387, ZN => n13334);
   U2433 : OAI22_X1 port map( A1 => n16344, A2 => n12323, B1 => n16341, B2 => 
                           n11856, ZN => n13332);
   U2434 : OAI22_X1 port map( A1 => n16392, A2 => n14844, B1 => n16389, B2 => 
                           n11894, ZN => n13324);
   U2435 : OAI22_X1 port map( A1 => n16380, A2 => n15385, B1 => n16377, B2 => 
                           n14388, ZN => n13325);
   U2436 : OAI22_X1 port map( A1 => n16332, A2 => n15050, B1 => n16329, B2 => 
                           n12186, ZN => n13291);
   U2437 : OAI22_X1 port map( A1 => n16320, A2 => n15166, B1 => n16317, B2 => 
                           n14389, ZN => n13292);
   U2438 : OAI22_X1 port map( A1 => n16344, A2 => n12324, B1 => n16341, B2 => 
                           n11857, ZN => n13290);
   U2439 : OAI22_X1 port map( A1 => n16392, A2 => n14845, B1 => n16389, B2 => 
                           n11895, ZN => n13282);
   U2440 : OAI22_X1 port map( A1 => n16380, A2 => n15386, B1 => n16377, B2 => 
                           n14390, ZN => n13283);
   U2441 : OAI22_X1 port map( A1 => n16332, A2 => n15051, B1 => n16329, B2 => 
                           n12187, ZN => n13249);
   U2442 : OAI22_X1 port map( A1 => n16320, A2 => n15167, B1 => n16317, B2 => 
                           n14391, ZN => n13250);
   U2443 : OAI22_X1 port map( A1 => n16344, A2 => n12325, B1 => n16341, B2 => 
                           n11858, ZN => n13248);
   U2444 : OAI22_X1 port map( A1 => n16392, A2 => n14846, B1 => n16389, B2 => 
                           n11896, ZN => n13240);
   U2445 : OAI22_X1 port map( A1 => n16380, A2 => n15387, B1 => n16377, B2 => 
                           n14392, ZN => n13241);
   U2446 : OAI22_X1 port map( A1 => n16332, A2 => n15052, B1 => n16329, B2 => 
                           n12188, ZN => n13207);
   U2447 : OAI22_X1 port map( A1 => n16320, A2 => n15168, B1 => n16317, B2 => 
                           n14393, ZN => n13208);
   U2448 : OAI22_X1 port map( A1 => n16344, A2 => n12326, B1 => n16341, B2 => 
                           n11860, ZN => n13206);
   U2449 : OAI22_X1 port map( A1 => n16392, A2 => n14847, B1 => n16389, B2 => 
                           n11897, ZN => n13198);
   U2450 : OAI22_X1 port map( A1 => n16380, A2 => n15388, B1 => n16377, B2 => 
                           n14394, ZN => n13199);
   U2451 : OAI22_X1 port map( A1 => n16332, A2 => n15053, B1 => n16329, B2 => 
                           n12189, ZN => n13165);
   U2452 : OAI22_X1 port map( A1 => n16320, A2 => n15170, B1 => n16317, B2 => 
                           n14395, ZN => n13166);
   U2453 : OAI22_X1 port map( A1 => n16344, A2 => n12327, B1 => n16341, B2 => 
                           n11862, ZN => n13164);
   U2454 : OAI22_X1 port map( A1 => n16392, A2 => n14848, B1 => n16389, B2 => 
                           n11898, ZN => n13156);
   U2455 : OAI22_X1 port map( A1 => n16380, A2 => n15389, B1 => n16377, B2 => 
                           n14408, ZN => n13157);
   U2456 : OAI22_X1 port map( A1 => n16332, A2 => n15055, B1 => n16329, B2 => 
                           n12190, ZN => n13123);
   U2457 : OAI22_X1 port map( A1 => n16320, A2 => n15171, B1 => n16317, B2 => 
                           n14398, ZN => n13124);
   U2458 : OAI22_X1 port map( A1 => n16344, A2 => n12328, B1 => n16341, B2 => 
                           n11863, ZN => n13122);
   U2459 : OAI22_X1 port map( A1 => n16392, A2 => n14849, B1 => n16389, B2 => 
                           n11899, ZN => n13114);
   U2460 : OAI22_X1 port map( A1 => n16380, A2 => n15391, B1 => n16377, B2 => 
                           n14409, ZN => n13115);
   U2461 : OAI22_X1 port map( A1 => n16332, A2 => n15056, B1 => n16329, B2 => 
                           n12191, ZN => n13081);
   U2462 : OAI22_X1 port map( A1 => n16320, A2 => n15172, B1 => n16317, B2 => 
                           n14399, ZN => n13082);
   U2463 : OAI22_X1 port map( A1 => n16344, A2 => n12329, B1 => n16341, B2 => 
                           n11864, ZN => n13080);
   U2464 : OAI22_X1 port map( A1 => n16392, A2 => n14850, B1 => n16389, B2 => 
                           n11900, ZN => n13072);
   U2465 : OAI22_X1 port map( A1 => n16380, A2 => n15392, B1 => n16377, B2 => 
                           n14410, ZN => n13073);
   U2466 : OAI22_X1 port map( A1 => n16332, A2 => n15057, B1 => n16329, B2 => 
                           n12192, ZN => n13039);
   U2467 : OAI22_X1 port map( A1 => n16320, A2 => n15173, B1 => n16317, B2 => 
                           n14400, ZN => n13040);
   U2468 : OAI22_X1 port map( A1 => n16344, A2 => n12330, B1 => n16341, B2 => 
                           n11865, ZN => n13038);
   U2469 : OAI22_X1 port map( A1 => n16392, A2 => n14851, B1 => n16389, B2 => 
                           n11901, ZN => n13030);
   U2470 : OAI22_X1 port map( A1 => n16380, A2 => n15393, B1 => n16377, B2 => 
                           n14411, ZN => n13031);
   U2471 : OAI22_X1 port map( A1 => n16332, A2 => n15058, B1 => n16329, B2 => 
                           n12193, ZN => n12997);
   U2472 : OAI22_X1 port map( A1 => n16320, A2 => n15174, B1 => n16317, B2 => 
                           n14401, ZN => n12998);
   U2473 : OAI22_X1 port map( A1 => n16344, A2 => n12331, B1 => n16341, B2 => 
                           n11866, ZN => n12996);
   U2474 : OAI22_X1 port map( A1 => n16392, A2 => n14852, B1 => n16389, B2 => 
                           n11902, ZN => n12988);
   U2475 : OAI22_X1 port map( A1 => n16380, A2 => n15394, B1 => n16377, B2 => 
                           n14412, ZN => n12989);
   U2476 : OAI22_X1 port map( A1 => n16332, A2 => n15059, B1 => n16329, B2 => 
                           n12164, ZN => n12955);
   U2477 : OAI22_X1 port map( A1 => n16320, A2 => n15175, B1 => n16317, B2 => 
                           n14402, ZN => n12956);
   U2478 : OAI22_X1 port map( A1 => n16344, A2 => n12332, B1 => n16341, B2 => 
                           n11867, ZN => n12954);
   U2479 : OAI22_X1 port map( A1 => n16392, A2 => n14824, B1 => n16389, B2 => 
                           n11874, ZN => n12946);
   U2480 : OAI22_X1 port map( A1 => n16380, A2 => n15395, B1 => n16377, B2 => 
                           n14413, ZN => n12947);
   U2481 : OAI22_X1 port map( A1 => n16583, A2 => n15152, B1 => n16580, B2 => 
                           n14359, ZN => n12464);
   U2482 : OAI22_X1 port map( A1 => n16571, A2 => n15037, B1 => n16568, B2 => 
                           n12171, ZN => n12466);
   U2483 : OAI22_X1 port map( A1 => n16595, A2 => n12309, B1 => n16592, B2 => 
                           n11713, ZN => n12462);
   U2484 : OAI22_X1 port map( A1 => n16631, A2 => n14831, B1 => n16628, B2 => 
                           n14362, ZN => n12448);
   U2485 : OAI22_X1 port map( A1 => n16643, A2 => n14605, B1 => n16640, B2 => 
                           n11881, ZN => n12442);
   U2486 : OAI22_X1 port map( A1 => n16583, A2 => n15153, B1 => n16580, B2 => 
                           n14363, ZN => n12283);
   U2487 : OAI22_X1 port map( A1 => n16571, A2 => n15035, B1 => n16568, B2 => 
                           n12172, ZN => n12284);
   U2488 : OAI22_X1 port map( A1 => n16595, A2 => n12310, B1 => n16592, B2 => 
                           n11756, ZN => n12282);
   U2489 : OAI22_X1 port map( A1 => n16631, A2 => n14832, B1 => n16628, B2 => 
                           n14360, ZN => n12275);
   U2490 : OAI22_X1 port map( A1 => n16643, A2 => n14606, B1 => n16640, B2 => 
                           n11882, ZN => n12274);
   U2491 : OAI22_X1 port map( A1 => n16583, A2 => n15151, B1 => n16580, B2 => 
                           n14361, ZN => n12130);
   U2492 : OAI22_X1 port map( A1 => n16571, A2 => n15036, B1 => n16568, B2 => 
                           n12173, ZN => n12131);
   U2493 : OAI22_X1 port map( A1 => n16595, A2 => n12311, B1 => n16592, B2 => 
                           n11799, ZN => n12129);
   U2494 : OAI22_X1 port map( A1 => n16631, A2 => n14833, B1 => n16628, B2 => 
                           n14364, ZN => n12122);
   U2495 : OAI22_X1 port map( A1 => n16643, A2 => n14607, B1 => n16640, B2 => 
                           n11883, ZN => n12121);
   U2496 : OAI22_X1 port map( A1 => n16583, A2 => n15154, B1 => n16580, B2 => 
                           n14365, ZN => n11977);
   U2497 : OAI22_X1 port map( A1 => n16571, A2 => n15038, B1 => n16568, B2 => 
                           n12174, ZN => n11978);
   U2498 : OAI22_X1 port map( A1 => n16595, A2 => n12312, B1 => n16592, B2 => 
                           n11842, ZN => n11976);
   U2499 : OAI22_X1 port map( A1 => n16631, A2 => n14834, B1 => n16628, B2 => 
                           n14366, ZN => n11969);
   U2500 : OAI22_X1 port map( A1 => n16643, A2 => n14608, B1 => n16640, B2 => 
                           n11627, ZN => n11968);
   U2501 : OAI22_X1 port map( A1 => n16583, A2 => n15155, B1 => n16580, B2 => 
                           n14367, ZN => n11824);
   U2502 : OAI22_X1 port map( A1 => n16571, A2 => n15039, B1 => n16568, B2 => 
                           n12175, ZN => n11825);
   U2503 : OAI22_X1 port map( A1 => n16595, A2 => n12313, B1 => n16592, B2 => 
                           n11844, ZN => n11823);
   U2504 : OAI22_X1 port map( A1 => n16631, A2 => n14823, B1 => n16628, B2 => 
                           n14289, ZN => n11816);
   U2505 : OAI22_X1 port map( A1 => n16643, A2 => n14569, B1 => n16640, B2 => 
                           n11884, ZN => n11815);
   U2506 : OAI22_X1 port map( A1 => n16583, A2 => n15000, B1 => n16580, B2 => 
                           n14290, ZN => n11781);
   U2507 : OAI22_X1 port map( A1 => n16571, A2 => n14993, B1 => n16568, B2 => 
                           n12162, ZN => n11782);
   U2508 : OAI22_X1 port map( A1 => n16595, A2 => n12308, B1 => n16592, B2 => 
                           n11584, ZN => n11780);
   U2509 : OAI22_X1 port map( A1 => n16631, A2 => n14835, B1 => n16628, B2 => 
                           n14368, ZN => n11773);
   U2510 : OAI22_X1 port map( A1 => n16643, A2 => n14609, B1 => n16640, B2 => 
                           n11885, ZN => n11772);
   U2511 : OAI22_X1 port map( A1 => n16583, A2 => n15157, B1 => n16580, B2 => 
                           n14369, ZN => n11738);
   U2512 : OAI22_X1 port map( A1 => n16571, A2 => n15040, B1 => n16568, B2 => 
                           n12176, ZN => n11739);
   U2513 : OAI22_X1 port map( A1 => n16595, A2 => n12315, B1 => n16592, B2 => 
                           n11846, ZN => n11737);
   U2514 : OAI22_X1 port map( A1 => n16631, A2 => n14836, B1 => n16628, B2 => 
                           n14372, ZN => n11730);
   U2515 : OAI22_X1 port map( A1 => n16643, A2 => n14610, B1 => n16640, B2 => 
                           n11886, ZN => n11729);
   U2516 : OAI22_X1 port map( A1 => n16583, A2 => n15158, B1 => n16580, B2 => 
                           n14373, ZN => n11695);
   U2517 : OAI22_X1 port map( A1 => n16571, A2 => n15042, B1 => n16568, B2 => 
                           n12177, ZN => n11696);
   U2518 : OAI22_X1 port map( A1 => n16595, A2 => n12316, B1 => n16592, B2 => 
                           n11847, ZN => n11694);
   U2519 : OAI22_X1 port map( A1 => n16631, A2 => n14837, B1 => n16628, B2 => 
                           n14374, ZN => n11687);
   U2520 : OAI22_X1 port map( A1 => n16643, A2 => n14611, B1 => n16640, B2 => 
                           n11887, ZN => n11686);
   U2521 : OAI22_X1 port map( A1 => n16583, A2 => n15159, B1 => n16580, B2 => 
                           n14375, ZN => n11652);
   U2522 : OAI22_X1 port map( A1 => n16571, A2 => n15043, B1 => n16568, B2 => 
                           n12178, ZN => n11653);
   U2523 : OAI22_X1 port map( A1 => n16595, A2 => n12317, B1 => n16592, B2 => 
                           n11849, ZN => n11651);
   U2524 : OAI22_X1 port map( A1 => n16631, A2 => n14838, B1 => n16628, B2 => 
                           n14376, ZN => n11644);
   U2525 : OAI22_X1 port map( A1 => n16643, A2 => n14612, B1 => n16640, B2 => 
                           n11888, ZN => n11643);
   U2526 : OAI22_X1 port map( A1 => n16583, A2 => n15160, B1 => n16580, B2 => 
                           n14377, ZN => n11609);
   U2527 : OAI22_X1 port map( A1 => n16571, A2 => n15044, B1 => n16568, B2 => 
                           n12179, ZN => n11610);
   U2528 : OAI22_X1 port map( A1 => n16595, A2 => n12318, B1 => n16592, B2 => 
                           n11850, ZN => n11608);
   U2529 : OAI22_X1 port map( A1 => n16631, A2 => n14839, B1 => n16628, B2 => 
                           n14378, ZN => n11601);
   U2530 : OAI22_X1 port map( A1 => n16643, A2 => n14613, B1 => n16640, B2 => 
                           n11889, ZN => n11600);
   U2531 : OAI22_X1 port map( A1 => n16583, A2 => n15161, B1 => n16580, B2 => 
                           n14379, ZN => n11566);
   U2532 : OAI22_X1 port map( A1 => n16571, A2 => n15045, B1 => n16568, B2 => 
                           n12180, ZN => n11567);
   U2533 : OAI22_X1 port map( A1 => n16595, A2 => n12319, B1 => n16592, B2 => 
                           n11851, ZN => n11565);
   U2534 : OAI22_X1 port map( A1 => n16631, A2 => n14840, B1 => n16628, B2 => 
                           n14380, ZN => n11558);
   U2535 : OAI22_X1 port map( A1 => n16643, A2 => n14614, B1 => n16640, B2 => 
                           n11890, ZN => n11557);
   U2536 : OAI22_X1 port map( A1 => n16583, A2 => n15162, B1 => n16580, B2 => 
                           n14381, ZN => n11523);
   U2537 : OAI22_X1 port map( A1 => n16571, A2 => n15046, B1 => n16568, B2 => 
                           n12181, ZN => n11524);
   U2538 : OAI22_X1 port map( A1 => n16595, A2 => n12320, B1 => n16592, B2 => 
                           n11852, ZN => n11522);
   U2539 : OAI22_X1 port map( A1 => n16631, A2 => n14841, B1 => n16628, B2 => 
                           n14382, ZN => n11515);
   U2540 : OAI22_X1 port map( A1 => n16643, A2 => n14615, B1 => n16640, B2 => 
                           n11891, ZN => n11514);
   U2541 : OAI22_X1 port map( A1 => n16584, A2 => n15163, B1 => n16581, B2 => 
                           n14383, ZN => n11480);
   U2542 : OAI22_X1 port map( A1 => n16572, A2 => n15047, B1 => n16569, B2 => 
                           n12182, ZN => n11481);
   U2543 : OAI22_X1 port map( A1 => n16596, A2 => n12321, B1 => n16593, B2 => 
                           n11854, ZN => n11479);
   U2544 : OAI22_X1 port map( A1 => n16632, A2 => n14842, B1 => n16629, B2 => 
                           n14384, ZN => n11472);
   U2545 : OAI22_X1 port map( A1 => n16644, A2 => n14616, B1 => n16641, B2 => 
                           n11892, ZN => n11471);
   U2546 : OAI22_X1 port map( A1 => n16584, A2 => n15164, B1 => n16581, B2 => 
                           n14385, ZN => n11436);
   U2547 : OAI22_X1 port map( A1 => n16572, A2 => n15048, B1 => n16569, B2 => 
                           n12183, ZN => n11437);
   U2548 : OAI22_X1 port map( A1 => n16596, A2 => n12322, B1 => n16593, B2 => 
                           n11855, ZN => n11435);
   U2549 : OAI22_X1 port map( A1 => n16632, A2 => n14843, B1 => n16629, B2 => 
                           n14386, ZN => n11428);
   U2550 : OAI22_X1 port map( A1 => n16644, A2 => n14617, B1 => n16641, B2 => 
                           n11893, ZN => n11427);
   U2551 : OAI22_X1 port map( A1 => n16584, A2 => n15165, B1 => n16581, B2 => 
                           n14387, ZN => n11393);
   U2552 : OAI22_X1 port map( A1 => n16572, A2 => n15049, B1 => n16569, B2 => 
                           n12185, ZN => n11394);
   U2553 : OAI22_X1 port map( A1 => n16596, A2 => n12323, B1 => n16593, B2 => 
                           n11856, ZN => n11392);
   U2554 : OAI22_X1 port map( A1 => n16632, A2 => n14844, B1 => n16629, B2 => 
                           n14388, ZN => n11385);
   U2555 : OAI22_X1 port map( A1 => n16644, A2 => n14618, B1 => n16641, B2 => 
                           n11894, ZN => n11384);
   U2556 : OAI22_X1 port map( A1 => n16584, A2 => n15166, B1 => n16581, B2 => 
                           n14389, ZN => n11350);
   U2557 : OAI22_X1 port map( A1 => n16572, A2 => n15050, B1 => n16569, B2 => 
                           n12186, ZN => n11351);
   U2558 : OAI22_X1 port map( A1 => n16596, A2 => n12324, B1 => n16593, B2 => 
                           n11857, ZN => n11349);
   U2559 : OAI22_X1 port map( A1 => n16632, A2 => n14845, B1 => n16629, B2 => 
                           n14390, ZN => n11342);
   U2560 : OAI22_X1 port map( A1 => n16644, A2 => n14619, B1 => n16641, B2 => 
                           n11895, ZN => n11341);
   U2561 : OAI22_X1 port map( A1 => n16584, A2 => n15167, B1 => n16581, B2 => 
                           n14391, ZN => n11307);
   U2562 : OAI22_X1 port map( A1 => n16572, A2 => n15051, B1 => n16569, B2 => 
                           n12187, ZN => n11308);
   U2563 : OAI22_X1 port map( A1 => n16596, A2 => n12325, B1 => n16593, B2 => 
                           n11858, ZN => n11306);
   U2564 : OAI22_X1 port map( A1 => n16632, A2 => n14846, B1 => n16629, B2 => 
                           n14392, ZN => n11299);
   U2565 : OAI22_X1 port map( A1 => n16644, A2 => n14620, B1 => n16641, B2 => 
                           n11896, ZN => n11298);
   U2566 : OAI22_X1 port map( A1 => n16584, A2 => n15168, B1 => n16581, B2 => 
                           n14393, ZN => n11264);
   U2567 : OAI22_X1 port map( A1 => n16572, A2 => n15052, B1 => n16569, B2 => 
                           n12188, ZN => n11265);
   U2568 : OAI22_X1 port map( A1 => n16596, A2 => n12326, B1 => n16593, B2 => 
                           n11860, ZN => n11263);
   U2569 : OAI22_X1 port map( A1 => n16632, A2 => n14847, B1 => n16629, B2 => 
                           n14394, ZN => n11256);
   U2570 : OAI22_X1 port map( A1 => n16644, A2 => n14621, B1 => n16641, B2 => 
                           n11897, ZN => n11255);
   U2571 : OAI22_X1 port map( A1 => n16584, A2 => n15170, B1 => n16581, B2 => 
                           n14395, ZN => n11221);
   U2572 : OAI22_X1 port map( A1 => n16572, A2 => n15053, B1 => n16569, B2 => 
                           n12189, ZN => n11222);
   U2573 : OAI22_X1 port map( A1 => n16596, A2 => n12327, B1 => n16593, B2 => 
                           n11862, ZN => n11220);
   U2574 : OAI22_X1 port map( A1 => n16632, A2 => n14848, B1 => n16629, B2 => 
                           n14408, ZN => n11213);
   U2575 : OAI22_X1 port map( A1 => n16644, A2 => n14622, B1 => n16641, B2 => 
                           n11898, ZN => n11212);
   U2576 : OAI22_X1 port map( A1 => n16584, A2 => n15171, B1 => n16581, B2 => 
                           n14398, ZN => n11178);
   U2577 : OAI22_X1 port map( A1 => n16572, A2 => n15055, B1 => n16569, B2 => 
                           n12190, ZN => n11179);
   U2578 : OAI22_X1 port map( A1 => n16596, A2 => n12328, B1 => n16593, B2 => 
                           n11863, ZN => n11177);
   U2579 : OAI22_X1 port map( A1 => n16632, A2 => n14849, B1 => n16629, B2 => 
                           n14409, ZN => n11170);
   U2580 : OAI22_X1 port map( A1 => n16644, A2 => n14623, B1 => n16641, B2 => 
                           n11899, ZN => n11169);
   U2581 : OAI22_X1 port map( A1 => n16584, A2 => n15172, B1 => n16581, B2 => 
                           n14399, ZN => n11135);
   U2582 : OAI22_X1 port map( A1 => n16572, A2 => n15056, B1 => n16569, B2 => 
                           n12191, ZN => n11136);
   U2583 : OAI22_X1 port map( A1 => n16596, A2 => n12329, B1 => n16593, B2 => 
                           n11864, ZN => n11134);
   U2584 : OAI22_X1 port map( A1 => n16632, A2 => n14850, B1 => n16629, B2 => 
                           n14410, ZN => n11127);
   U2585 : OAI22_X1 port map( A1 => n16644, A2 => n14624, B1 => n16641, B2 => 
                           n11900, ZN => n11126);
   U2586 : OAI22_X1 port map( A1 => n16584, A2 => n15173, B1 => n16581, B2 => 
                           n14400, ZN => n11092);
   U2587 : OAI22_X1 port map( A1 => n16572, A2 => n15057, B1 => n16569, B2 => 
                           n12192, ZN => n11093);
   U2588 : OAI22_X1 port map( A1 => n16596, A2 => n12330, B1 => n16593, B2 => 
                           n11865, ZN => n11091);
   U2589 : OAI22_X1 port map( A1 => n16632, A2 => n14851, B1 => n16629, B2 => 
                           n14411, ZN => n11084);
   U2590 : OAI22_X1 port map( A1 => n16644, A2 => n14625, B1 => n16641, B2 => 
                           n11901, ZN => n11083);
   U2591 : OAI22_X1 port map( A1 => n16584, A2 => n15174, B1 => n16581, B2 => 
                           n14401, ZN => n11049);
   U2592 : OAI22_X1 port map( A1 => n16572, A2 => n15058, B1 => n16569, B2 => 
                           n12193, ZN => n11050);
   U2593 : OAI22_X1 port map( A1 => n16596, A2 => n12331, B1 => n16593, B2 => 
                           n11866, ZN => n11048);
   U2594 : OAI22_X1 port map( A1 => n16632, A2 => n14852, B1 => n16629, B2 => 
                           n14412, ZN => n11041);
   U2595 : OAI22_X1 port map( A1 => n16644, A2 => n14626, B1 => n16641, B2 => 
                           n11902, ZN => n11040);
   U2596 : OAI22_X1 port map( A1 => n16584, A2 => n15175, B1 => n16581, B2 => 
                           n14402, ZN => n11006);
   U2597 : OAI22_X1 port map( A1 => n16572, A2 => n15059, B1 => n16569, B2 => 
                           n12164, ZN => n11007);
   U2598 : OAI22_X1 port map( A1 => n16596, A2 => n12332, B1 => n16593, B2 => 
                           n11867, ZN => n11005);
   U2599 : OAI22_X1 port map( A1 => n16632, A2 => n14824, B1 => n16629, B2 => 
                           n14413, ZN => n10998);
   U2600 : OAI22_X1 port map( A1 => n16644, A2 => n14598, B1 => n16641, B2 => 
                           n11874, ZN => n10997);
   U2601 : OAI22_X1 port map( A1 => n17727, A2 => n15575, B1 => n17724, B2 => 
                           n12309, ZN => n12390);
   U2602 : OAI22_X1 port map( A1 => n17763, A2 => n15369, B1 => n17760, B2 => 
                           n14484, ZN => n12387);
   U2603 : OAI22_X1 port map( A1 => n17751, A2 => n12356, B1 => n17748, B2 => 
                           n12018, ZN => n12388);
   U2604 : OAI22_X1 port map( A1 => n17679, A2 => n14547, B1 => n17676, B2 => 
                           n11951, ZN => n12398);
   U2605 : OAI22_X1 port map( A1 => n17715, A2 => n15576, B1 => n17712, B2 => 
                           n11713, ZN => n12395);
   U2606 : OAI22_X1 port map( A1 => n17703, A2 => n15574, B1 => n17700, B2 => 
                           n14669, ZN => n12396);
   U2607 : OAI22_X1 port map( A1 => n17727, A2 => n15577, B1 => n17724, B2 => 
                           n12310, ZN => n12236);
   U2608 : OAI22_X1 port map( A1 => n17763, A2 => n15370, B1 => n17760, B2 => 
                           n14485, ZN => n12233);
   U2609 : OAI22_X1 port map( A1 => n17751, A2 => n12358, B1 => n17748, B2 => 
                           n12019, ZN => n12234);
   U2610 : OAI22_X1 port map( A1 => n17679, A2 => n14548, B1 => n17676, B2 => 
                           n11952, ZN => n12244);
   U2611 : OAI22_X1 port map( A1 => n17715, A2 => n15580, B1 => n17712, B2 => 
                           n11756, ZN => n12241);
   U2612 : OAI22_X1 port map( A1 => n17703, A2 => n15661, B1 => n17700, B2 => 
                           n14645, ZN => n12242);
   U2613 : OAI22_X1 port map( A1 => n17727, A2 => n15586, B1 => n17724, B2 => 
                           n12311, ZN => n12081);
   U2614 : OAI22_X1 port map( A1 => n17763, A2 => n15401, B1 => n17760, B2 => 
                           n14486, ZN => n12078);
   U2615 : OAI22_X1 port map( A1 => n17751, A2 => n12360, B1 => n17748, B2 => 
                           n12020, ZN => n12079);
   U2616 : OAI22_X1 port map( A1 => n17679, A2 => n14549, B1 => n17676, B2 => 
                           n11995, ZN => n12089);
   U2617 : OAI22_X1 port map( A1 => n17715, A2 => n15581, B1 => n17712, B2 => 
                           n11799, ZN => n12086);
   U2618 : OAI22_X1 port map( A1 => n17703, A2 => n15578, B1 => n17700, B2 => 
                           n14643, ZN => n12087);
   U2619 : OAI22_X1 port map( A1 => n17727, A2 => n15587, B1 => n17724, B2 => 
                           n12312, ZN => n11928);
   U2620 : OAI22_X1 port map( A1 => n17763, A2 => n15402, B1 => n17760, B2 => 
                           n14487, ZN => n11925);
   U2621 : OAI22_X1 port map( A1 => n17751, A2 => n12340, B1 => n17748, B2 => 
                           n12016, ZN => n11926);
   U2622 : OAI22_X1 port map( A1 => n17679, A2 => n14536, B1 => n17676, B2 => 
                           n11905, ZN => n11936);
   U2623 : OAI22_X1 port map( A1 => n17715, A2 => n15582, B1 => n17712, B2 => 
                           n11842, ZN => n11933);
   U2624 : OAI22_X1 port map( A1 => n17703, A2 => n15361, B1 => n17700, B2 => 
                           n14635, ZN => n11934);
   U2625 : OAI22_X1 port map( A1 => n17727, A2 => n15588, B1 => n17724, B2 => 
                           n12313, ZN => n10485);
   U2626 : OAI22_X1 port map( A1 => n17763, A2 => n15351, B1 => n17760, B2 => 
                           n14294, ZN => n10482);
   U2627 : OAI22_X1 port map( A1 => n17751, A2 => n12341, B1 => n17748, B2 => 
                           n12017, ZN => n10483);
   U2628 : OAI22_X1 port map( A1 => n17679, A2 => n14550, B1 => n17676, B2 => 
                           n11997, ZN => n10493);
   U2629 : OAI22_X1 port map( A1 => n17715, A2 => n15583, B1 => n17712, B2 => 
                           n11844, ZN => n10490);
   U2630 : OAI22_X1 port map( A1 => n17703, A2 => n15362, B1 => n17700, B2 => 
                           n14636, ZN => n10491);
   U2631 : OAI22_X1 port map( A1 => n17727, A2 => n15363, B1 => n17724, B2 => 
                           n12308, ZN => n10375);
   U2632 : OAI22_X1 port map( A1 => n17763, A2 => n15352, B1 => n17760, B2 => 
                           n14295, ZN => n10372);
   U2633 : OAI22_X1 port map( A1 => n17751, A2 => n12364, B1 => n17748, B2 => 
                           n12021, ZN => n10373);
   U2634 : OAI22_X1 port map( A1 => n17679, A2 => n14537, B1 => n17676, B2 => 
                           n11906, ZN => n10383);
   U2635 : OAI22_X1 port map( A1 => n17715, A2 => n15584, B1 => n17712, B2 => 
                           n11584, ZN => n10380);
   U2636 : OAI22_X1 port map( A1 => n17703, A2 => n15364, B1 => n17700, B2 => 
                           n14637, ZN => n10381);
   U2637 : OAI22_X1 port map( A1 => n17727, A2 => n15589, B1 => n17724, B2 => 
                           n12315, ZN => n10263);
   U2638 : OAI22_X1 port map( A1 => n17763, A2 => n15403, B1 => n17760, B2 => 
                           n14488, ZN => n10260);
   U2639 : OAI22_X1 port map( A1 => n17751, A2 => n12366, B1 => n17748, B2 => 
                           n12022, ZN => n10261);
   U2640 : OAI22_X1 port map( A1 => n17679, A2 => n14551, B1 => n17676, B2 => 
                           n11998, ZN => n10271);
   U2641 : OAI22_X1 port map( A1 => n17715, A2 => n15579, B1 => n17712, B2 => 
                           n11846, ZN => n10268);
   U2642 : OAI22_X1 port map( A1 => n17703, A2 => n15637, B1 => n17700, B2 => 
                           n14646, ZN => n10269);
   U2643 : OAI22_X1 port map( A1 => n17727, A2 => n15591, B1 => n17724, B2 => 
                           n12316, ZN => n7627);
   U2644 : OAI22_X1 port map( A1 => n17763, A2 => n15404, B1 => n17760, B2 => 
                           n14489, ZN => n7624);
   U2645 : OAI22_X1 port map( A1 => n17751, A2 => n12368, B1 => n17748, B2 => 
                           n12023, ZN => n7625);
   U2646 : OAI22_X1 port map( A1 => n17679, A2 => n14552, B1 => n17676, B2 => 
                           n11999, ZN => n7635);
   U2647 : OAI22_X1 port map( A1 => n17715, A2 => n15592, B1 => n17712, B2 => 
                           n11847, ZN => n7632);
   U2648 : OAI22_X1 port map( A1 => n17703, A2 => n15638, B1 => n17700, B2 => 
                           n14647, ZN => n7633);
   U2649 : OAI22_X1 port map( A1 => n17727, A2 => n15593, B1 => n17724, B2 => 
                           n12317, ZN => n7512);
   U2650 : OAI22_X1 port map( A1 => n17763, A2 => n15405, B1 => n17760, B2 => 
                           n14490, ZN => n7509);
   U2651 : OAI22_X1 port map( A1 => n17751, A2 => n12407, B1 => n17748, B2 => 
                           n12024, ZN => n7510);
   U2652 : OAI22_X1 port map( A1 => n17679, A2 => n14553, B1 => n17676, B2 => 
                           n12000, ZN => n7520);
   U2653 : OAI22_X1 port map( A1 => n17715, A2 => n15594, B1 => n17712, B2 => 
                           n11849, ZN => n7517);
   U2654 : OAI22_X1 port map( A1 => n17703, A2 => n15639, B1 => n17700, B2 => 
                           n14648, ZN => n7518);
   U2655 : OAI22_X1 port map( A1 => n17727, A2 => n15595, B1 => n17724, B2 => 
                           n12318, ZN => n7403);
   U2656 : OAI22_X1 port map( A1 => n17763, A2 => n15406, B1 => n17760, B2 => 
                           n14491, ZN => n7400);
   U2657 : OAI22_X1 port map( A1 => n17751, A2 => n12409, B1 => n17748, B2 => 
                           n12025, ZN => n7401);
   U2658 : OAI22_X1 port map( A1 => n17679, A2 => n14554, B1 => n17676, B2 => 
                           n12001, ZN => n7411);
   U2659 : OAI22_X1 port map( A1 => n17715, A2 => n15596, B1 => n17712, B2 => 
                           n11850, ZN => n7408);
   U2660 : OAI22_X1 port map( A1 => n17703, A2 => n15640, B1 => n17700, B2 => 
                           n14649, ZN => n7409);
   U2661 : OAI22_X1 port map( A1 => n17727, A2 => n15597, B1 => n17724, B2 => 
                           n12319, ZN => n7294);
   U2662 : OAI22_X1 port map( A1 => n17763, A2 => n15407, B1 => n17760, B2 => 
                           n14492, ZN => n7291);
   U2663 : OAI22_X1 port map( A1 => n17751, A2 => n12411, B1 => n17748, B2 => 
                           n12026, ZN => n7292);
   U2664 : OAI22_X1 port map( A1 => n17679, A2 => n14555, B1 => n17676, B2 => 
                           n12002, ZN => n7302);
   U2665 : OAI22_X1 port map( A1 => n17715, A2 => n15598, B1 => n17712, B2 => 
                           n11851, ZN => n7299);
   U2666 : OAI22_X1 port map( A1 => n17703, A2 => n15641, B1 => n17700, B2 => 
                           n14650, ZN => n7300);
   U2667 : OAI22_X1 port map( A1 => n17728, A2 => n15599, B1 => n17725, B2 => 
                           n12320, ZN => n7180);
   U2668 : OAI22_X1 port map( A1 => n17764, A2 => n15408, B1 => n17761, B2 => 
                           n14493, ZN => n7177);
   U2669 : OAI22_X1 port map( A1 => n17752, A2 => n12600, B1 => n17749, B2 => 
                           n12027, ZN => n7178);
   U2670 : OAI22_X1 port map( A1 => n17680, A2 => n14556, B1 => n17677, B2 => 
                           n12003, ZN => n7188);
   U2671 : OAI22_X1 port map( A1 => n17716, A2 => n15600, B1 => n17713, B2 => 
                           n11852, ZN => n7185);
   U2672 : OAI22_X1 port map( A1 => n17704, A2 => n15642, B1 => n17701, B2 => 
                           n14651, ZN => n7186);
   U2673 : OAI22_X1 port map( A1 => n17728, A2 => n15601, B1 => n17725, B2 => 
                           n12321, ZN => n7071);
   U2674 : OAI22_X1 port map( A1 => n17764, A2 => n15409, B1 => n17761, B2 => 
                           n14494, ZN => n7068);
   U2675 : OAI22_X1 port map( A1 => n17752, A2 => n12652, B1 => n17749, B2 => 
                           n12028, ZN => n7069);
   U2676 : OAI22_X1 port map( A1 => n17680, A2 => n14557, B1 => n17677, B2 => 
                           n12004, ZN => n7079);
   U2677 : OAI22_X1 port map( A1 => n17716, A2 => n15602, B1 => n17713, B2 => 
                           n11854, ZN => n7076);
   U2678 : OAI22_X1 port map( A1 => n17704, A2 => n15643, B1 => n17701, B2 => 
                           n14652, ZN => n7077);
   U2679 : OAI22_X1 port map( A1 => n17728, A2 => n15603, B1 => n17725, B2 => 
                           n12322, ZN => n6962);
   U2680 : OAI22_X1 port map( A1 => n17764, A2 => n15410, B1 => n17761, B2 => 
                           n14495, ZN => n6959);
   U2681 : OAI22_X1 port map( A1 => n17752, A2 => n13996, B1 => n17749, B2 => 
                           n12030, ZN => n6960);
   U2682 : OAI22_X1 port map( A1 => n17680, A2 => n14558, B1 => n17677, B2 => 
                           n12005, ZN => n6970);
   U2683 : OAI22_X1 port map( A1 => n17716, A2 => n15604, B1 => n17713, B2 => 
                           n11855, ZN => n6967);
   U2684 : OAI22_X1 port map( A1 => n17704, A2 => n15644, B1 => n17701, B2 => 
                           n14653, ZN => n6968);
   U2685 : OAI22_X1 port map( A1 => n17728, A2 => n15605, B1 => n17725, B2 => 
                           n12323, ZN => n6853);
   U2686 : OAI22_X1 port map( A1 => n17764, A2 => n15411, B1 => n17761, B2 => 
                           n14496, ZN => n6850);
   U2687 : OAI22_X1 port map( A1 => n17752, A2 => n14008, B1 => n17749, B2 => 
                           n12031, ZN => n6851);
   U2688 : OAI22_X1 port map( A1 => n17680, A2 => n14559, B1 => n17677, B2 => 
                           n12006, ZN => n6861);
   U2689 : OAI22_X1 port map( A1 => n17716, A2 => n15606, B1 => n17713, B2 => 
                           n11856, ZN => n6858);
   U2690 : OAI22_X1 port map( A1 => n17704, A2 => n15645, B1 => n17701, B2 => 
                           n14654, ZN => n6859);
   U2691 : OAI22_X1 port map( A1 => n17728, A2 => n15607, B1 => n17725, B2 => 
                           n12324, ZN => n6744);
   U2692 : OAI22_X1 port map( A1 => n17764, A2 => n15412, B1 => n17761, B2 => 
                           n14497, ZN => n6741);
   U2693 : OAI22_X1 port map( A1 => n17752, A2 => n14015, B1 => n17749, B2 => 
                           n12032, ZN => n6742);
   U2694 : OAI22_X1 port map( A1 => n17680, A2 => n14560, B1 => n17677, B2 => 
                           n12007, ZN => n6752);
   U2695 : OAI22_X1 port map( A1 => n17716, A2 => n15608, B1 => n17713, B2 => 
                           n11857, ZN => n6749);
   U2696 : OAI22_X1 port map( A1 => n17704, A2 => n15646, B1 => n17701, B2 => 
                           n14655, ZN => n6750);
   U2697 : OAI22_X1 port map( A1 => n17728, A2 => n15609, B1 => n17725, B2 => 
                           n12325, ZN => n6601);
   U2698 : OAI22_X1 port map( A1 => n17764, A2 => n15413, B1 => n17761, B2 => 
                           n14498, ZN => n6598);
   U2699 : OAI22_X1 port map( A1 => n17752, A2 => n14035, B1 => n17749, B2 => 
                           n12033, ZN => n6599);
   U2700 : OAI22_X1 port map( A1 => n17680, A2 => n14561, B1 => n17677, B2 => 
                           n12008, ZN => n6610);
   U2701 : OAI22_X1 port map( A1 => n17716, A2 => n15610, B1 => n17713, B2 => 
                           n11858, ZN => n6606);
   U2702 : OAI22_X1 port map( A1 => n17704, A2 => n15647, B1 => n17701, B2 => 
                           n14656, ZN => n6607);
   U2703 : OAI22_X1 port map( A1 => n17728, A2 => n15611, B1 => n17725, B2 => 
                           n12326, ZN => n6414);
   U2704 : OAI22_X1 port map( A1 => n17764, A2 => n15414, B1 => n17761, B2 => 
                           n14499, ZN => n6411);
   U2705 : OAI22_X1 port map( A1 => n17752, A2 => n14037, B1 => n17749, B2 => 
                           n12034, ZN => n6412);
   U2706 : OAI22_X1 port map( A1 => n17680, A2 => n14562, B1 => n17677, B2 => 
                           n12009, ZN => n6425);
   U2707 : OAI22_X1 port map( A1 => n17716, A2 => n15612, B1 => n17713, B2 => 
                           n11860, ZN => n6420);
   U2708 : OAI22_X1 port map( A1 => n17704, A2 => n15648, B1 => n17701, B2 => 
                           n14657, ZN => n6421);
   U2709 : OAI22_X1 port map( A1 => n17728, A2 => n15613, B1 => n17725, B2 => 
                           n12327, ZN => n6227);
   U2710 : OAI22_X1 port map( A1 => n17764, A2 => n15415, B1 => n17761, B2 => 
                           n14500, ZN => n6224);
   U2711 : OAI22_X1 port map( A1 => n17752, A2 => n14039, B1 => n17749, B2 => 
                           n12035, ZN => n6225);
   U2712 : OAI22_X1 port map( A1 => n17680, A2 => n14563, B1 => n17677, B2 => 
                           n12010, ZN => n6238);
   U2713 : OAI22_X1 port map( A1 => n17716, A2 => n15626, B1 => n17713, B2 => 
                           n11862, ZN => n6234);
   U2714 : OAI22_X1 port map( A1 => n17704, A2 => n15649, B1 => n17701, B2 => 
                           n14658, ZN => n6236);
   U2715 : OAI22_X1 port map( A1 => n17728, A2 => n15616, B1 => n17725, B2 => 
                           n12328, ZN => n6040);
   U2716 : OAI22_X1 port map( A1 => n17764, A2 => n15416, B1 => n17761, B2 => 
                           n14501, ZN => n6037);
   U2717 : OAI22_X1 port map( A1 => n17752, A2 => n14041, B1 => n17749, B2 => 
                           n12036, ZN => n6038);
   U2718 : OAI22_X1 port map( A1 => n17680, A2 => n14564, B1 => n17677, B2 => 
                           n12011, ZN => n6051);
   U2719 : OAI22_X1 port map( A1 => n17716, A2 => n15627, B1 => n17713, B2 => 
                           n11863, ZN => n6048);
   U2720 : OAI22_X1 port map( A1 => n17704, A2 => n15650, B1 => n17701, B2 => 
                           n14659, ZN => n6049);
   U2721 : OAI22_X1 port map( A1 => n17728, A2 => n15617, B1 => n17725, B2 => 
                           n12329, ZN => n5854);
   U2722 : OAI22_X1 port map( A1 => n17764, A2 => n15417, B1 => n17761, B2 => 
                           n14502, ZN => n5850);
   U2723 : OAI22_X1 port map( A1 => n17752, A2 => n14043, B1 => n17749, B2 => 
                           n12037, ZN => n5851);
   U2724 : OAI22_X1 port map( A1 => n17680, A2 => n14565, B1 => n17677, B2 => 
                           n12012, ZN => n5866);
   U2725 : OAI22_X1 port map( A1 => n17716, A2 => n15628, B1 => n17713, B2 => 
                           n11864, ZN => n5861);
   U2726 : OAI22_X1 port map( A1 => n17704, A2 => n15651, B1 => n17701, B2 => 
                           n14660, ZN => n5862);
   U2727 : OAI22_X1 port map( A1 => n17728, A2 => n15618, B1 => n17725, B2 => 
                           n12330, ZN => n5669);
   U2728 : OAI22_X1 port map( A1 => n17764, A2 => n15418, B1 => n17761, B2 => 
                           n14503, ZN => n5664);
   U2729 : OAI22_X1 port map( A1 => n17752, A2 => n14045, B1 => n17749, B2 => 
                           n12038, ZN => n5665);
   U2730 : OAI22_X1 port map( A1 => n17680, A2 => n14566, B1 => n17677, B2 => 
                           n12013, ZN => n5680);
   U2731 : OAI22_X1 port map( A1 => n17716, A2 => n15629, B1 => n17713, B2 => 
                           n11865, ZN => n5674);
   U2732 : OAI22_X1 port map( A1 => n17704, A2 => n15652, B1 => n17701, B2 => 
                           n14661, ZN => n5677);
   U2733 : OAI22_X1 port map( A1 => n17728, A2 => n15619, B1 => n17725, B2 => 
                           n12331, ZN => n5482);
   U2734 : OAI22_X1 port map( A1 => n17764, A2 => n15419, B1 => n17761, B2 => 
                           n14504, ZN => n5478);
   U2735 : OAI22_X1 port map( A1 => n17752, A2 => n14047, B1 => n17749, B2 => 
                           n12039, ZN => n5480);
   U2736 : OAI22_X1 port map( A1 => n17680, A2 => n14567, B1 => n17677, B2 => 
                           n12014, ZN => n5493);
   U2737 : OAI22_X1 port map( A1 => n17716, A2 => n15630, B1 => n17713, B2 => 
                           n11866, ZN => n5489);
   U2738 : OAI22_X1 port map( A1 => n17704, A2 => n15653, B1 => n17701, B2 => 
                           n14662, ZN => n5491);
   U2739 : OAI22_X1 port map( A1 => n17727, A2 => n15590, B1 => n17724, B2 => 
                           n12314, ZN => n14148);
   U2740 : OAI22_X1 port map( A1 => n17763, A2 => n15427, B1 => n17760, B2 => 
                           n14477, ZN => n14113);
   U2741 : OAI22_X1 port map( A1 => n17751, A2 => n12355, B1 => n17748, B2 => 
                           n12047, ZN => n14126);
   U2742 : OAI22_X1 port map( A1 => n17679, A2 => n14546, B1 => n17676, B2 => 
                           n11950, ZN => n14175);
   U2743 : OAI22_X1 port map( A1 => n17715, A2 => n15585, B1 => n17712, B2 => 
                           n11845, ZN => n14157);
   U2744 : OAI22_X1 port map( A1 => n17703, A2 => n15317, B1 => n17700, B2 => 
                           n14634, ZN => n14161);
   U2745 : OAI22_X1 port map( A1 => n14960, A2 => n16427, B1 => n14284, B2 => 
                           n16424, ZN => n13900);
   U2746 : OAI22_X1 port map( A1 => n14961, A2 => n16427, B1 => n14285, B2 => 
                           n16424, ZN => n13858);
   U2747 : OAI22_X1 port map( A1 => n14962, A2 => n16427, B1 => n14286, B2 => 
                           n16424, ZN => n13816);
   U2748 : OAI22_X1 port map( A1 => n14980, A2 => n16427, B1 => n14287, B2 => 
                           n16424, ZN => n13774);
   U2749 : OAI22_X1 port map( A1 => n14963, A2 => n16427, B1 => n14071, B2 => 
                           n16424, ZN => n13732);
   U2750 : OAI22_X1 port map( A1 => n14964, A2 => n16427, B1 => n14212, B2 => 
                           n16424, ZN => n13690);
   U2751 : OAI22_X1 port map( A1 => n14868, A2 => n16427, B1 => n14053, B2 => 
                           n16424, ZN => n13648);
   U2752 : OAI22_X1 port map( A1 => n14965, A2 => n16427, B1 => n14216, B2 => 
                           n16424, ZN => n13606);
   U2753 : OAI22_X1 port map( A1 => n14966, A2 => n16427, B1 => n14219, B2 => 
                           n16424, ZN => n13564);
   U2754 : OAI22_X1 port map( A1 => n14967, A2 => n16427, B1 => n14225, B2 => 
                           n16424, ZN => n13522);
   U2755 : OAI22_X1 port map( A1 => n14968, A2 => n16427, B1 => n14227, B2 => 
                           n16424, ZN => n13480);
   U2756 : OAI22_X1 port map( A1 => n14969, A2 => n16427, B1 => n14230, B2 => 
                           n16424, ZN => n13438);
   U2757 : OAI22_X1 port map( A1 => n14970, A2 => n16428, B1 => n14235, B2 => 
                           n16425, ZN => n13396);
   U2758 : OAI22_X1 port map( A1 => n14971, A2 => n16428, B1 => n14242, B2 => 
                           n16425, ZN => n13354);
   U2759 : OAI22_X1 port map( A1 => n14972, A2 => n16428, B1 => n14243, B2 => 
                           n16425, ZN => n13312);
   U2760 : OAI22_X1 port map( A1 => n14973, A2 => n16428, B1 => n14246, B2 => 
                           n16425, ZN => n13270);
   U2761 : OAI22_X1 port map( A1 => n14974, A2 => n16428, B1 => n14255, B2 => 
                           n16425, ZN => n13228);
   U2762 : OAI22_X1 port map( A1 => n14975, A2 => n16428, B1 => n14261, B2 => 
                           n16425, ZN => n13186);
   U2763 : OAI22_X1 port map( A1 => n14976, A2 => n16428, B1 => n14264, B2 => 
                           n16425, ZN => n13144);
   U2764 : OAI22_X1 port map( A1 => n14977, A2 => n16428, B1 => n14269, B2 => 
                           n16425, ZN => n13102);
   U2765 : OAI22_X1 port map( A1 => n14978, A2 => n16428, B1 => n14270, B2 => 
                           n16425, ZN => n13060);
   U2766 : OAI22_X1 port map( A1 => n14981, A2 => n16428, B1 => n14271, B2 => 
                           n16425, ZN => n13018);
   U2767 : OAI22_X1 port map( A1 => n14982, A2 => n16428, B1 => n14268, B2 => 
                           n16425, ZN => n12976);
   U2768 : OAI22_X1 port map( A1 => n14979, A2 => n16428, B1 => n14272, B2 => 
                           n16425, ZN => n12934);
   U2769 : OAI22_X1 port map( A1 => n16680, A2 => n14965, B1 => n14216, B2 => 
                           n16677, ZN => n11674);
   U2770 : OAI22_X1 port map( A1 => n16680, A2 => n14966, B1 => n14219, B2 => 
                           n16677, ZN => n11631);
   U2771 : OAI22_X1 port map( A1 => n16680, A2 => n14967, B1 => n14225, B2 => 
                           n16677, ZN => n11588);
   U2772 : OAI22_X1 port map( A1 => n16680, A2 => n14968, B1 => n14227, B2 => 
                           n16677, ZN => n11545);
   U2773 : OAI22_X1 port map( A1 => n16680, A2 => n14969, B1 => n14230, B2 => 
                           n16677, ZN => n11502);
   U2774 : OAI22_X1 port map( A1 => n16680, A2 => n14970, B1 => n14235, B2 => 
                           n16677, ZN => n11458);
   U2775 : OAI22_X1 port map( A1 => n16680, A2 => n14971, B1 => n14242, B2 => 
                           n16677, ZN => n11415);
   U2776 : OAI22_X1 port map( A1 => n16680, A2 => n14972, B1 => n14243, B2 => 
                           n16677, ZN => n11372);
   U2777 : OAI22_X1 port map( A1 => n16680, A2 => n14973, B1 => n14246, B2 => 
                           n16677, ZN => n11329);
   U2778 : OAI22_X1 port map( A1 => n16680, A2 => n14974, B1 => n14255, B2 => 
                           n16677, ZN => n11286);
   U2779 : OAI22_X1 port map( A1 => n16680, A2 => n14975, B1 => n14261, B2 => 
                           n16677, ZN => n11243);
   U2780 : OAI22_X1 port map( A1 => n16680, A2 => n14976, B1 => n14264, B2 => 
                           n16676, ZN => n11200);
   U2781 : OAI22_X1 port map( A1 => n16679, A2 => n14977, B1 => n14269, B2 => 
                           n16676, ZN => n11157);
   U2782 : OAI22_X1 port map( A1 => n16679, A2 => n14978, B1 => n14270, B2 => 
                           n16676, ZN => n11114);
   U2783 : OAI22_X1 port map( A1 => n16679, A2 => n14981, B1 => n14271, B2 => 
                           n16676, ZN => n11071);
   U2784 : OAI22_X1 port map( A1 => n16679, A2 => n14982, B1 => n14268, B2 => 
                           n16676, ZN => n11028);
   U2785 : OAI22_X1 port map( A1 => n16679, A2 => n14979, B1 => n14272, B2 => 
                           n16677, ZN => n10985);
   U2786 : OAI22_X1 port map( A1 => n16679, A2 => n14983, B1 => n14273, B2 => 
                           n16676, ZN => n10942);
   U2787 : OAI22_X1 port map( A1 => n16679, A2 => n14984, B1 => n14274, B2 => 
                           n16676, ZN => n10899);
   U2788 : OAI22_X1 port map( A1 => n16679, A2 => n14985, B1 => n14275, B2 => 
                           n16676, ZN => n10856);
   U2789 : OAI22_X1 port map( A1 => n16679, A2 => n14986, B1 => n14276, B2 => 
                           n16676, ZN => n10813);
   U2790 : OAI22_X1 port map( A1 => n16679, A2 => n14987, B1 => n14277, B2 => 
                           n16676, ZN => n10770);
   U2791 : OAI22_X1 port map( A1 => n16679, A2 => n14988, B1 => n14278, B2 => 
                           n16676, ZN => n10727);
   U2792 : OAI22_X1 port map( A1 => n16679, A2 => n14860, B1 => n14052, B2 => 
                           n16676, ZN => n10668);
   U2793 : NOR3_X1 port map( A1 => N9908, A2 => n14178, A3 => N9910, ZN => 
                           n14193);
   U2794 : INV_X1 port map( A => n14095, ZN => n14090);
   U2795 : OAI22_X1 port map( A1 => n16372, A2 => n15203, B1 => n16369, B2 => 
                           n12199, ZN => n12906);
   U2796 : OAI22_X1 port map( A1 => n16372, A2 => n15204, B1 => n16369, B2 => 
                           n12200, ZN => n12864);
   U2797 : OAI22_X1 port map( A1 => n16372, A2 => n15205, B1 => n16369, B2 => 
                           n12201, ZN => n12822);
   U2798 : OAI22_X1 port map( A1 => n16372, A2 => n15206, B1 => n16369, B2 => 
                           n12202, ZN => n12780);
   U2799 : OAI22_X1 port map( A1 => n16372, A2 => n15207, B1 => n16369, B2 => 
                           n12203, ZN => n12738);
   U2800 : OAI22_X1 port map( A1 => n16372, A2 => n15208, B1 => n16369, B2 => 
                           n12204, ZN => n12696);
   U2801 : OAI22_X1 port map( A1 => n16372, A2 => n14873, B1 => n16369, B2 => 
                           n12161, ZN => n12653);
   U2802 : OAI22_X1 port map( A1 => n16372, A2 => n15209, B1 => n16369, B2 => 
                           n12307, ZN => n12554);
   U2803 : OAI22_X1 port map( A1 => n16624, A2 => n15203, B1 => n16621, B2 => 
                           n12199, ZN => n10956);
   U2804 : OAI22_X1 port map( A1 => n16624, A2 => n15204, B1 => n16621, B2 => 
                           n12200, ZN => n10913);
   U2805 : OAI22_X1 port map( A1 => n16624, A2 => n15205, B1 => n16621, B2 => 
                           n12201, ZN => n10870);
   U2806 : OAI22_X1 port map( A1 => n16624, A2 => n15206, B1 => n16621, B2 => 
                           n12202, ZN => n10827);
   U2807 : OAI22_X1 port map( A1 => n16624, A2 => n15207, B1 => n16621, B2 => 
                           n12203, ZN => n10784);
   U2808 : OAI22_X1 port map( A1 => n16624, A2 => n15208, B1 => n16621, B2 => 
                           n12204, ZN => n10741);
   U2809 : OAI22_X1 port map( A1 => n16624, A2 => n14873, B1 => n16621, B2 => 
                           n12161, ZN => n10685);
   U2810 : OAI22_X1 port map( A1 => n16624, A2 => n15209, B1 => n16621, B2 => 
                           n12307, ZN => n10557);
   U2811 : NAND2_X1 port map( A1 => n14007, A2 => n14020, ZN => n14009);
   U2812 : BUF_X1 port map( A => n4240, Z => n17635);
   U2813 : BUF_X1 port map( A => n4240, Z => n17634);
   U2814 : BUF_X1 port map( A => n12527, Z => n16416);
   U2815 : BUF_X1 port map( A => n12527, Z => n16415);
   U2816 : BUF_X1 port map( A => n10525, Z => n16668);
   U2817 : BUF_X1 port map( A => n10525, Z => n16667);
   U2818 : OAI22_X1 port map( A1 => n16370, A2 => n15181, B1 => n16367, B2 => 
                           n12205, ZN => n13934);
   U2819 : OAI22_X1 port map( A1 => n16370, A2 => n15182, B1 => n16367, B2 => 
                           n12206, ZN => n13872);
   U2820 : OAI22_X1 port map( A1 => n16370, A2 => n15183, B1 => n16367, B2 => 
                           n12207, ZN => n13830);
   U2821 : OAI22_X1 port map( A1 => n16370, A2 => n15001, B1 => n16367, B2 => 
                           n12208, ZN => n13788);
   U2822 : OAI22_X1 port map( A1 => n16370, A2 => n15002, B1 => n16367, B2 => 
                           n12195, ZN => n13746);
   U2823 : OAI22_X1 port map( A1 => n16370, A2 => n15184, B1 => n16367, B2 => 
                           n12209, ZN => n13704);
   U2824 : OAI22_X1 port map( A1 => n16370, A2 => n15185, B1 => n16367, B2 => 
                           n12210, ZN => n13662);
   U2825 : OAI22_X1 port map( A1 => n16370, A2 => n15186, B1 => n16367, B2 => 
                           n12211, ZN => n13620);
   U2826 : OAI22_X1 port map( A1 => n16370, A2 => n15187, B1 => n16367, B2 => 
                           n12212, ZN => n13578);
   U2827 : OAI22_X1 port map( A1 => n16370, A2 => n15188, B1 => n16367, B2 => 
                           n12213, ZN => n13536);
   U2828 : OAI22_X1 port map( A1 => n16370, A2 => n15189, B1 => n16367, B2 => 
                           n12214, ZN => n13494);
   U2829 : OAI22_X1 port map( A1 => n16370, A2 => n15190, B1 => n16367, B2 => 
                           n12215, ZN => n13452);
   U2830 : OAI22_X1 port map( A1 => n16371, A2 => n15191, B1 => n16368, B2 => 
                           n12253, ZN => n13410);
   U2831 : OAI22_X1 port map( A1 => n16371, A2 => n15192, B1 => n16368, B2 => 
                           n12254, ZN => n13368);
   U2832 : OAI22_X1 port map( A1 => n16371, A2 => n15193, B1 => n16368, B2 => 
                           n12255, ZN => n13326);
   U2833 : OAI22_X1 port map( A1 => n16371, A2 => n15194, B1 => n16368, B2 => 
                           n12256, ZN => n13284);
   U2834 : OAI22_X1 port map( A1 => n16371, A2 => n15195, B1 => n16368, B2 => 
                           n12257, ZN => n13242);
   U2835 : OAI22_X1 port map( A1 => n16371, A2 => n15196, B1 => n16368, B2 => 
                           n12258, ZN => n13200);
   U2836 : OAI22_X1 port map( A1 => n16371, A2 => n15197, B1 => n16368, B2 => 
                           n12301, ZN => n13158);
   U2837 : OAI22_X1 port map( A1 => n16371, A2 => n15198, B1 => n16368, B2 => 
                           n12303, ZN => n13116);
   U2838 : OAI22_X1 port map( A1 => n16371, A2 => n15199, B1 => n16368, B2 => 
                           n12304, ZN => n13074);
   U2839 : OAI22_X1 port map( A1 => n16371, A2 => n15200, B1 => n16368, B2 => 
                           n12305, ZN => n13032);
   U2840 : OAI22_X1 port map( A1 => n16371, A2 => n15201, B1 => n16368, B2 => 
                           n12306, ZN => n12990);
   U2841 : OAI22_X1 port map( A1 => n16371, A2 => n15202, B1 => n16368, B2 => 
                           n12198, ZN => n12948);
   U2842 : OAI22_X1 port map( A1 => n16622, A2 => n15181, B1 => n16619, B2 => 
                           n12205, ZN => n12453);
   U2843 : OAI22_X1 port map( A1 => n16622, A2 => n15182, B1 => n16619, B2 => 
                           n12206, ZN => n12276);
   U2844 : OAI22_X1 port map( A1 => n16622, A2 => n15183, B1 => n16619, B2 => 
                           n12207, ZN => n12123);
   U2845 : OAI22_X1 port map( A1 => n16622, A2 => n15001, B1 => n16619, B2 => 
                           n12208, ZN => n11970);
   U2846 : OAI22_X1 port map( A1 => n16622, A2 => n15002, B1 => n16619, B2 => 
                           n12195, ZN => n11817);
   U2847 : OAI22_X1 port map( A1 => n16622, A2 => n15184, B1 => n16619, B2 => 
                           n12209, ZN => n11774);
   U2848 : OAI22_X1 port map( A1 => n16622, A2 => n15185, B1 => n16619, B2 => 
                           n12210, ZN => n11731);
   U2849 : OAI22_X1 port map( A1 => n16622, A2 => n15186, B1 => n16619, B2 => 
                           n12211, ZN => n11688);
   U2850 : OAI22_X1 port map( A1 => n16622, A2 => n15187, B1 => n16619, B2 => 
                           n12212, ZN => n11645);
   U2851 : OAI22_X1 port map( A1 => n16622, A2 => n15188, B1 => n16619, B2 => 
                           n12213, ZN => n11602);
   U2852 : OAI22_X1 port map( A1 => n16622, A2 => n15189, B1 => n16619, B2 => 
                           n12214, ZN => n11559);
   U2853 : OAI22_X1 port map( A1 => n16622, A2 => n15190, B1 => n16619, B2 => 
                           n12215, ZN => n11516);
   U2854 : OAI22_X1 port map( A1 => n16623, A2 => n15191, B1 => n16620, B2 => 
                           n12253, ZN => n11473);
   U2855 : OAI22_X1 port map( A1 => n16623, A2 => n15192, B1 => n16620, B2 => 
                           n12254, ZN => n11429);
   U2856 : OAI22_X1 port map( A1 => n16623, A2 => n15193, B1 => n16620, B2 => 
                           n12255, ZN => n11386);
   U2857 : OAI22_X1 port map( A1 => n16623, A2 => n15194, B1 => n16620, B2 => 
                           n12256, ZN => n11343);
   U2858 : OAI22_X1 port map( A1 => n16623, A2 => n15195, B1 => n16620, B2 => 
                           n12257, ZN => n11300);
   U2859 : OAI22_X1 port map( A1 => n16623, A2 => n15196, B1 => n16620, B2 => 
                           n12258, ZN => n11257);
   U2860 : OAI22_X1 port map( A1 => n16623, A2 => n15197, B1 => n16620, B2 => 
                           n12301, ZN => n11214);
   U2861 : OAI22_X1 port map( A1 => n16623, A2 => n15198, B1 => n16620, B2 => 
                           n12303, ZN => n11171);
   U2862 : OAI22_X1 port map( A1 => n16623, A2 => n15199, B1 => n16620, B2 => 
                           n12304, ZN => n11128);
   U2863 : OAI22_X1 port map( A1 => n16623, A2 => n15200, B1 => n16620, B2 => 
                           n12305, ZN => n11085);
   U2864 : OAI22_X1 port map( A1 => n16623, A2 => n15201, B1 => n16620, B2 => 
                           n12306, ZN => n11042);
   U2865 : OAI22_X1 port map( A1 => n16623, A2 => n15202, B1 => n16620, B2 => 
                           n12198, ZN => n10999);
   U2866 : NOR2_X1 port map( A1 => n12492, A2 => n12493, ZN => n10649);
   U2867 : NAND2_X1 port map( A1 => n14158, A2 => n14095, ZN => n4184);
   U2868 : NAND2_X1 port map( A1 => n14094, A2 => n14095, ZN => n4119);
   U2869 : NAND2_X1 port map( A1 => n14104, A2 => n14095, ZN => n4126);
   U2870 : NAND2_X1 port map( A1 => n14107, A2 => n14095, ZN => n4135);
   U2871 : NAND2_X1 port map( A1 => n14108, A2 => n14095, ZN => n4133);
   U2872 : NOR2_X1 port map( A1 => n14100, A2 => n14020, ZN => n14180);
   U2873 : NAND2_X1 port map( A1 => datain(6), A2 => n18038, ZN => n7652);
   U2874 : NAND2_X1 port map( A1 => n14137, A2 => N9925, ZN => n14131);
   U2875 : NAND2_X1 port map( A1 => n14202, A2 => N9925, ZN => n14145);
   U2876 : NAND2_X1 port map( A1 => n14263, A2 => N273, ZN => n14066);
   U2877 : NOR2_X1 port map( A1 => n14172, A2 => n14020, ZN => n14204);
   U2878 : BUF_X1 port map( A => n4223, Z => n17665);
   U2879 : BUF_X1 port map( A => n4223, Z => n17664);
   U2880 : BUF_X1 port map( A => n4202, Z => n17689);
   U2881 : BUF_X1 port map( A => n4202, Z => n17688);
   U2882 : BUF_X1 port map( A => n4240, Z => n17636);
   U2883 : NOR2_X1 port map( A1 => n13976, A2 => N46301, ZN => n13937);
   U2884 : NOR2_X1 port map( A1 => n12495, A2 => N45787, ZN => n12456);
   U2885 : NOR2_X1 port map( A1 => n13975, A2 => N46300, ZN => n13961);
   U2886 : NOR2_X1 port map( A1 => n12494, A2 => N45786, ZN => n12480);
   U2887 : NOR2_X1 port map( A1 => N46301, A2 => N46300, ZN => n13958);
   U2888 : NOR2_X1 port map( A1 => N45787, A2 => N45786, ZN => n12475);
   U2889 : NOR2_X1 port map( A1 => n14144, A2 => n14820, ZN => n14179);
   U2890 : OAI22_X1 port map( A1 => n16700, A2 => n14960, B1 => n16439, B2 => 
                           n16692, ZN => n7759);
   U2891 : OAI22_X1 port map( A1 => n17585, A2 => n14284, B1 => n16439, B2 => 
                           n17577, ZN => n7798);
   U2892 : OAI22_X1 port map( A1 => n17836, A2 => n14506, B1 => n16439, B2 => 
                           n17839, ZN => n7800);
   U2893 : OAI22_X1 port map( A1 => n17880, A2 => n15574, B1 => n16439, B2 => 
                           n17883, ZN => n7801);
   U2894 : OAI22_X1 port map( A1 => n17923, A2 => n15432, B1 => n16439, B2 => 
                           n17926, ZN => n7802);
   U2895 : OAI22_X1 port map( A1 => n17965, A2 => n15245, B1 => n16439, B2 => 
                           n17968, ZN => n7803);
   U2896 : OAI22_X1 port map( A1 => n18012, A2 => n12055, B1 => n16439, B2 => 
                           n18003, ZN => n7804);
   U2897 : OAI22_X1 port map( A1 => n16887, A2 => n15369, B1 => n16439, B2 => 
                           n16888, ZN => n7806);
   U2898 : OAI22_X1 port map( A1 => n16910, A2 => n14484, B1 => n16439, B2 => 
                           n16911, ZN => n7807);
   U2899 : OAI22_X1 port map( A1 => n16943, A2 => n14547, B1 => n16440, B2 => 
                           n16934, ZN => n7808);
   U2900 : OAI22_X1 port map( A1 => n16956, A2 => n14772, B1 => n16440, B2 => 
                           n16957, ZN => n7809);
   U2901 : OAI22_X1 port map( A1 => n16976, A2 => n14888, B1 => n16440, B2 => 
                           n16977, ZN => n7810);
   U2902 : OAI22_X1 port map( A1 => n16999, A2 => n14427, B1 => n16440, B2 => 
                           n17000, ZN => n7811);
   U2903 : OAI22_X1 port map( A1 => n17032, A2 => n12171, B1 => n16440, B2 => 
                           n17023, ZN => n7812);
   U2904 : OAI22_X1 port map( A1 => n17058, A2 => n14359, B1 => n16440, B2 => 
                           n17049, ZN => n7813);
   U2905 : OAI22_X1 port map( A1 => n17084, A2 => n15575, B1 => n16440, B2 => 
                           n17075, ZN => n7814);
   U2906 : OAI22_X1 port map( A1 => n17110, A2 => n11713, B1 => n16440, B2 => 
                           n17101, ZN => n7815);
   U2907 : OAI22_X1 port map( A1 => n17136, A2 => n15736, B1 => n16440, B2 => 
                           n17127, ZN => n7816);
   U2908 : OAI22_X1 port map( A1 => n17171, A2 => n12018, B1 => n16440, B2 => 
                           n17172, ZN => n7818);
   U2909 : OAI22_X1 port map( A1 => n17192, A2 => n14300, B1 => n16440, B2 => 
                           n17193, ZN => n7819);
   U2910 : OAI22_X1 port map( A1 => n17251, A2 => n12205, B1 => n16441, B2 => 
                           n17242, ZN => n7821);
   U2911 : OAI22_X1 port map( A1 => n17303, A2 => n14605, B1 => n16441, B2 => 
                           n17294, ZN => n7823);
   U2912 : OAI22_X1 port map( A1 => n17329, A2 => n15292, B1 => n16441, B2 => 
                           n17320, ZN => n7824);
   U2913 : OAI22_X1 port map( A1 => n17355, A2 => n15072, B1 => n16441, B2 => 
                           n17346, ZN => n7825);
   U2914 : OAI22_X1 port map( A1 => n17381, A2 => n14426, B1 => n16441, B2 => 
                           n17372, ZN => n7826);
   U2915 : OAI22_X1 port map( A1 => n17407, A2 => n14329, B1 => n16441, B2 => 
                           n17398, ZN => n7827);
   U2916 : OAI22_X1 port map( A1 => n17433, A2 => n15326, B1 => n16441, B2 => 
                           n17424, ZN => n7828);
   U2917 : OAI22_X1 port map( A1 => n17459, A2 => n14711, B1 => n16441, B2 => 
                           n17451, ZN => n7829);
   U2918 : OAI22_X1 port map( A1 => n17485, A2 => n15758, B1 => n16441, B2 => 
                           n17476, ZN => n7830);
   U2919 : OAI22_X1 port map( A1 => n17511, A2 => n15576, B1 => n16441, B2 => 
                           n17502, ZN => n7831);
   U2920 : OAI22_X1 port map( A1 => n16700, A2 => n14961, B1 => n16445, B2 => 
                           n16692, ZN => n7833);
   U2921 : OAI22_X1 port map( A1 => n17585, A2 => n14285, B1 => n16445, B2 => 
                           n17577, ZN => n7872);
   U2922 : OAI22_X1 port map( A1 => n17838, A2 => n14507, B1 => n16445, B2 => 
                           n17839, ZN => n7874);
   U2923 : OAI22_X1 port map( A1 => n17860, A2 => n15124, B1 => n16445, B2 => 
                           n17861, ZN => n7875);
   U2924 : OAI22_X1 port map( A1 => n17925, A2 => n15433, B1 => n16445, B2 => 
                           n17926, ZN => n7876);
   U2925 : OAI22_X1 port map( A1 => n17946, A2 => n14911, B1 => n16445, B2 => 
                           n17947, ZN => n7877);
   U2926 : OAI22_X1 port map( A1 => n18012, A2 => n12052, B1 => n16445, B2 => 
                           n18003, ZN => n7878);
   U2927 : OAI22_X1 port map( A1 => n18025, A2 => n14570, B1 => n16445, B2 => 
                           n18016, ZN => n7879);
   U2928 : OAI22_X1 port map( A1 => n16887, A2 => n15370, B1 => n16445, B2 => 
                           n16888, ZN => n7880);
   U2929 : OAI22_X1 port map( A1 => n16943, A2 => n14548, B1 => n16446, B2 => 
                           n16934, ZN => n7882);
   U2930 : OAI22_X1 port map( A1 => n16945, A2 => n11952, B1 => n16446, B2 => 
                           n16946, ZN => n7883);
   U2931 : OAI22_X1 port map( A1 => n16976, A2 => n14889, B1 => n16446, B2 => 
                           n16977, ZN => n7884);
   U2932 : OAI22_X1 port map( A1 => n17032, A2 => n12172, B1 => n16446, B2 => 
                           n17023, ZN => n7886);
   U2933 : OAI22_X1 port map( A1 => n17045, A2 => n15035, B1 => n16446, B2 => 
                           n17036, ZN => n7887);
   U2934 : OAI22_X1 port map( A1 => n17084, A2 => n15577, B1 => n16446, B2 => 
                           n17075, ZN => n7888);
   U2935 : OAI22_X1 port map( A1 => n17097, A2 => n15496, B1 => n16446, B2 => 
                           n17088, ZN => n7889);
   U2936 : OAI22_X1 port map( A1 => n17136, A2 => n15737, B1 => n16446, B2 => 
                           n17127, ZN => n7890);
   U2937 : OAI22_X1 port map( A1 => n17137, A2 => n14679, B1 => n16446, B2 => 
                           n17138, ZN => n7891);
   U2938 : OAI22_X1 port map( A1 => n17171, A2 => n12019, B1 => n16446, B2 => 
                           n17172, ZN => n7892);
   U2939 : OAI22_X1 port map( A1 => n17182, A2 => n12358, B1 => n16446, B2 => 
                           n17183, ZN => n7893);
   U2940 : OAI22_X1 port map( A1 => n17238, A2 => n15371, B1 => n16447, B2 => 
                           n17229, ZN => n7895);
   U2941 : OAI22_X1 port map( A1 => n17290, A2 => n14360, B1 => n16447, B2 => 
                           n17281, ZN => n7897);
   U2942 : OAI22_X1 port map( A1 => n17329, A2 => n15293, B1 => n16447, B2 => 
                           n17320, ZN => n7898);
   U2943 : OAI22_X1 port map( A1 => n17342, A2 => n11882, B1 => n16447, B2 => 
                           n17333, ZN => n7899);
   U2944 : OAI22_X1 port map( A1 => n17381, A2 => n14428, B1 => n16447, B2 => 
                           n17372, ZN => n7900);
   U2945 : OAI22_X1 port map( A1 => n17394, A2 => n14714, B1 => n16447, B2 => 
                           n17385, ZN => n7901);
   U2946 : OAI22_X1 port map( A1 => n17433, A2 => n15327, B1 => n16447, B2 => 
                           n17424, ZN => n7902);
   U2947 : OAI22_X1 port map( A1 => n17446, A2 => n12359, B1 => n16447, B2 => 
                           n17437, ZN => n7903);
   U2948 : OAI22_X1 port map( A1 => n17485, A2 => n15759, B1 => n16447, B2 => 
                           n17476, ZN => n7904);
   U2949 : OAI22_X1 port map( A1 => n17498, A2 => n14773, B1 => n16447, B2 => 
                           n17489, ZN => n7905);
   U2950 : OAI22_X1 port map( A1 => n16700, A2 => n14962, B1 => n16451, B2 => 
                           n16692, ZN => n7907);
   U2951 : OAI22_X1 port map( A1 => n17838, A2 => n14508, B1 => n16451, B2 => 
                           n17840, ZN => n7948);
   U2952 : OAI22_X1 port map( A1 => n17860, A2 => n15125, B1 => n16451, B2 => 
                           n17861, ZN => n7949);
   U2953 : OAI22_X1 port map( A1 => n17882, A2 => n15578, B1 => n16451, B2 => 
                           n17883, ZN => n7950);
   U2954 : OAI22_X1 port map( A1 => n17904, A2 => n14643, B1 => n16451, B2 => 
                           n17905, ZN => n7951);
   U2955 : OAI22_X1 port map( A1 => n18012, A2 => n12053, B1 => n16451, B2 => 
                           n18003, ZN => n7952);
   U2956 : OAI22_X1 port map( A1 => n18025, A2 => n14571, B1 => n16451, B2 => 
                           n18016, ZN => n7953);
   U2957 : OAI22_X1 port map( A1 => n16877, A2 => n14940, B1 => n16451, B2 => 
                           n16878, ZN => n7955);
   U2958 : OAI22_X1 port map( A1 => n16943, A2 => n14549, B1 => n16452, B2 => 
                           n16934, ZN => n7956);
   U2959 : OAI22_X1 port map( A1 => n16945, A2 => n11995, B1 => n16452, B2 => 
                           n16946, ZN => n7957);
   U2960 : OAI22_X1 port map( A1 => n16956, A2 => n14776, B1 => n16452, B2 => 
                           n16957, ZN => n7958);
   U2961 : OAI22_X1 port map( A1 => n16966, A2 => n15468, B1 => n16452, B2 => 
                           n16967, ZN => n7959);
   U2962 : OAI22_X1 port map( A1 => n17032, A2 => n12173, B1 => n16452, B2 => 
                           n17023, ZN => n7960);
   U2963 : OAI22_X1 port map( A1 => n17045, A2 => n15036, B1 => n16452, B2 => 
                           n17036, ZN => n7961);
   U2964 : OAI22_X1 port map( A1 => n17058, A2 => n14361, B1 => n16452, B2 => 
                           n17049, ZN => n7962);
   U2965 : OAI22_X1 port map( A1 => n17071, A2 => n15151, B1 => n16452, B2 => 
                           n17062, ZN => n7963);
   U2966 : OAI22_X1 port map( A1 => n17136, A2 => n15738, B1 => n16452, B2 => 
                           n17127, ZN => n7964);
   U2967 : OAI22_X1 port map( A1 => n17137, A2 => n14680, B1 => n16452, B2 => 
                           n17138, ZN => n7965);
   U2968 : OAI22_X1 port map( A1 => n17160, A2 => n15006, B1 => n16452, B2 => 
                           n17161, ZN => n7967);
   U2969 : OAI22_X1 port map( A1 => n17238, A2 => n15372, B1 => n16453, B2 => 
                           n17229, ZN => n7969);
   U2970 : OAI22_X1 port map( A1 => n17251, A2 => n12207, B1 => n16453, B2 => 
                           n17242, ZN => n7970);
   U2971 : OAI22_X1 port map( A1 => n17264, A2 => n14833, B1 => n16453, B2 => 
                           n17255, ZN => n7971);
   U2972 : OAI22_X1 port map( A1 => n17329, A2 => n15294, B1 => n16453, B2 => 
                           n17320, ZN => n7972);
   U2973 : OAI22_X1 port map( A1 => n17342, A2 => n11883, B1 => n16453, B2 => 
                           n17333, ZN => n7973);
   U2974 : OAI22_X1 port map( A1 => n17355, A2 => n15076, B1 => n16453, B2 => 
                           n17346, ZN => n7974);
   U2975 : OAI22_X1 port map( A1 => n17368, A2 => n15671, B1 => n16453, B2 => 
                           n17359, ZN => n7975);
   U2976 : OAI22_X1 port map( A1 => n17433, A2 => n15328, B1 => n16453, B2 => 
                           n17424, ZN => n7976);
   U2977 : OAI22_X1 port map( A1 => n17446, A2 => n12361, B1 => n16453, B2 => 
                           n17437, ZN => n7977);
   U2978 : OAI22_X1 port map( A1 => n17459, A2 => n14715, B1 => n16453, B2 => 
                           n17451, ZN => n7978);
   U2979 : OAI22_X1 port map( A1 => n17472, A2 => n15523, B1 => n16453, B2 => 
                           n17463, ZN => n7979);
   U2980 : OAI22_X1 port map( A1 => n17123, A2 => n12309, B1 => n17115, B2 => 
                           n16437, ZN => n7780);
   U2981 : OAI22_X1 port map( A1 => n17316, A2 => n15699, B1 => n17308, B2 => 
                           n16438, ZN => n7788);
   U2982 : OAI22_X1 port map( A1 => n17420, A2 => n15210, B1 => n17412, B2 => 
                           n16438, ZN => n7792);
   U2983 : OAI22_X1 port map( A1 => n17123, A2 => n12310, B1 => n17114, B2 => 
                           n16443, ZN => n7855);
   U2984 : OAI22_X1 port map( A1 => n17316, A2 => n15700, B1 => n17307, B2 => 
                           n16444, ZN => n7863);
   U2985 : OAI22_X1 port map( A1 => n17420, A2 => n15211, B1 => n17411, B2 => 
                           n16444, ZN => n7867);
   U2986 : OAI22_X1 port map( A1 => n17123, A2 => n12311, B1 => n17114, B2 => 
                           n16449, ZN => n7931);
   U2987 : OAI22_X1 port map( A1 => n17316, A2 => n15701, B1 => n17307, B2 => 
                           n16450, ZN => n7939);
   U2988 : OAI22_X1 port map( A1 => n17420, A2 => n15212, B1 => n17411, B2 => 
                           n16450, ZN => n7943);
   U2989 : OAI22_X1 port map( A1 => n17122, A2 => n12312, B1 => n17114, B2 => 
                           n16457, ZN => n8005);
   U2990 : OAI22_X1 port map( A1 => n17315, A2 => n15702, B1 => n17307, B2 => 
                           n16458, ZN => n8013);
   U2991 : OAI22_X1 port map( A1 => n17122, A2 => n12313, B1 => n17115, B2 => 
                           n16710, ZN => n8133);
   U2992 : OAI22_X1 port map( A1 => n17419, A2 => n15213, B1 => n17411, B2 => 
                           n16711, ZN => n8149);
   U2993 : OAI22_X1 port map( A1 => n17315, A2 => n15703, B1 => n17308, B2 => 
                           n16719, ZN => n8213);
   U2994 : OAI22_X1 port map( A1 => n17419, A2 => n15214, B1 => n17412, B2 => 
                           n16720, ZN => n8221);
   U2995 : OAI22_X1 port map( A1 => n17123, A2 => n12314, B1 => n17115, B2 => 
                           n16705, ZN => n10093);
   U2996 : OAI22_X1 port map( A1 => n17316, A2 => n15721, B1 => n17308, B2 => 
                           n16703, ZN => n10109);
   U2997 : OAI22_X1 port map( A1 => n17420, A2 => n15239, B1 => n17412, B2 => 
                           n16703, ZN => n10117);
   U2998 : NOR2_X1 port map( A1 => n13981, A2 => n13982, ZN => n13962);
   U2999 : INV_X1 port map( A => n13983, ZN => n13982);
   U3000 : NOR2_X1 port map( A1 => n12500, A2 => n12501, ZN => n12481);
   U3001 : INV_X1 port map( A => n12502, ZN => n12501);
   U3002 : OAI22_X1 port map( A1 => n17484, A2 => n15764, B1 => n17476, B2 => 
                           n16730, ZN => n8322);
   U3003 : OAI22_X1 port map( A1 => n17497, A2 => n14781, B1 => n17490, B2 => 
                           n16730, ZN => n8323);
   U3004 : OAI22_X1 port map( A1 => n17510, A2 => n15579, B1 => n17503, B2 => 
                           n16730, ZN => n8324);
   U3005 : OAI22_X1 port map( A1 => n17446, A2 => n12357, B1 => n17438, B2 => 
                           n16438, ZN => n7793);
   U3006 : OAI22_X1 port map( A1 => n17472, A2 => n15521, B1 => n17464, B2 => 
                           n16438, ZN => n7794);
   U3007 : OAI22_X1 port map( A1 => n17498, A2 => n14771, B1 => n17490, B2 => 
                           n16438, ZN => n7795);
   U3008 : OAI22_X1 port map( A1 => n17459, A2 => n14713, B1 => n17451, B2 => 
                           n16444, ZN => n7868);
   U3009 : OAI22_X1 port map( A1 => n17472, A2 => n15522, B1 => n17463, B2 => 
                           n16444, ZN => n7869);
   U3010 : OAI22_X1 port map( A1 => n17511, A2 => n15580, B1 => n17503, B2 => 
                           n16444, ZN => n7870);
   U3011 : OAI22_X1 port map( A1 => n17485, A2 => n15760, B1 => n17476, B2 => 
                           n16450, ZN => n7944);
   U3012 : OAI22_X1 port map( A1 => n17498, A2 => n14775, B1 => n17489, B2 => 
                           n16450, ZN => n7945);
   U3013 : OAI22_X1 port map( A1 => n17511, A2 => n15581, B1 => n17502, B2 => 
                           n16450, ZN => n7946);
   U3014 : OAI22_X1 port map( A1 => n17432, A2 => n15329, B1 => n17425, B2 => 
                           n16458, ZN => n8022);
   U3015 : OAI22_X1 port map( A1 => n17445, A2 => n12362, B1 => n17437, B2 => 
                           n16458, ZN => n8023);
   U3016 : OAI22_X1 port map( A1 => n17458, A2 => n14717, B1 => n17451, B2 => 
                           n16458, ZN => n8024);
   U3017 : OAI22_X1 port map( A1 => n17471, A2 => n15524, B1 => n17464, B2 => 
                           n16458, ZN => n8025);
   U3018 : OAI22_X1 port map( A1 => n17484, A2 => n15761, B1 => n17476, B2 => 
                           n16459, ZN => n8026);
   U3019 : OAI22_X1 port map( A1 => n17497, A2 => n14777, B1 => n17489, B2 => 
                           n16459, ZN => n8027);
   U3020 : OAI22_X1 port map( A1 => n17510, A2 => n15582, B1 => n17502, B2 => 
                           n16459, ZN => n8028);
   U3021 : OAI22_X1 port map( A1 => n17432, A2 => n15330, B1 => n17425, B2 => 
                           n16711, ZN => n8150);
   U3022 : OAI22_X1 port map( A1 => n17445, A2 => n12363, B1 => n17438, B2 => 
                           n16711, ZN => n8151);
   U3023 : OAI22_X1 port map( A1 => n17458, A2 => n14718, B1 => n17451, B2 => 
                           n16711, ZN => n8152);
   U3024 : OAI22_X1 port map( A1 => n17471, A2 => n15525, B1 => n17463, B2 => 
                           n16711, ZN => n8153);
   U3025 : OAI22_X1 port map( A1 => n17484, A2 => n15762, B1 => n17477, B2 => 
                           n16712, ZN => n8154);
   U3026 : OAI22_X1 port map( A1 => n17497, A2 => n14778, B1 => n17490, B2 => 
                           n16712, ZN => n8155);
   U3027 : OAI22_X1 port map( A1 => n17510, A2 => n15583, B1 => n17503, B2 => 
                           n16712, ZN => n8156);
   U3028 : OAI22_X1 port map( A1 => n17432, A2 => n15331, B1 => n17424, B2 => 
                           n16720, ZN => n8222);
   U3029 : OAI22_X1 port map( A1 => n17445, A2 => n12365, B1 => n17437, B2 => 
                           n16720, ZN => n8223);
   U3030 : OAI22_X1 port map( A1 => n17458, A2 => n14720, B1 => n17451, B2 => 
                           n16720, ZN => n8224);
   U3031 : OAI22_X1 port map( A1 => n17471, A2 => n15526, B1 => n17463, B2 => 
                           n16720, ZN => n8225);
   U3032 : OAI22_X1 port map( A1 => n17484, A2 => n15763, B1 => n17477, B2 => 
                           n16721, ZN => n8226);
   U3033 : OAI22_X1 port map( A1 => n17497, A2 => n14780, B1 => n17490, B2 => 
                           n16721, ZN => n8227);
   U3034 : OAI22_X1 port map( A1 => n17510, A2 => n15584, B1 => n17503, B2 => 
                           n16721, ZN => n8228);
   U3035 : OAI22_X1 port map( A1 => n17432, A2 => n15332, B1 => n17424, B2 => 
                           n16729, ZN => n8318);
   U3036 : OAI22_X1 port map( A1 => n17445, A2 => n12367, B1 => n17437, B2 => 
                           n16729, ZN => n8319);
   U3037 : OAI22_X1 port map( A1 => n17458, A2 => n14722, B1 => n17451, B2 => 
                           n16729, ZN => n8320);
   U3038 : OAI22_X1 port map( A1 => n17431, A2 => n15333, B1 => n17424, B2 => 
                           n16736, ZN => n8390);
   U3039 : OAI22_X1 port map( A1 => n17433, A2 => n15349, B1 => n17425, B2 => 
                           n16703, ZN => n10118);
   U3040 : OAI22_X1 port map( A1 => n17446, A2 => n12348, B1 => n17438, B2 => 
                           n16702, ZN => n10119);
   U3041 : OAI22_X1 port map( A1 => n17459, A2 => n15318, B1 => n17451, B2 => 
                           n16703, ZN => n10120);
   U3042 : OAI22_X1 port map( A1 => n17472, A2 => n15458, B1 => n17464, B2 => 
                           n16702, ZN => n10121);
   U3043 : OAI22_X1 port map( A1 => n17485, A2 => n15781, B1 => n17477, B2 => 
                           n16702, ZN => n10122);
   U3044 : OAI22_X1 port map( A1 => n17498, A2 => n14815, B1 => n17489, B2 => 
                           n16702, ZN => n10123);
   U3045 : OAI22_X1 port map( A1 => n17511, A2 => n15585, B1 => n17502, B2 => 
                           n16702, ZN => n10124);
   U3046 : OAI22_X1 port map( A1 => n17045, A2 => n15037, B1 => n17036, B2 => 
                           n16437, ZN => n7777);
   U3047 : OAI22_X1 port map( A1 => n17071, A2 => n15152, B1 => n17062, B2 => 
                           n16437, ZN => n7778);
   U3048 : OAI22_X1 port map( A1 => n17097, A2 => n15495, B1 => n17088, B2 => 
                           n16437, ZN => n7779);
   U3049 : OAI22_X1 port map( A1 => n17238, A2 => n15373, B1 => n17229, B2 => 
                           n16438, ZN => n7785);
   U3050 : OAI22_X1 port map( A1 => n17264, A2 => n14831, B1 => n17255, B2 => 
                           n16438, ZN => n7786);
   U3051 : OAI22_X1 port map( A1 => n17290, A2 => n14362, B1 => n17281, B2 => 
                           n16438, ZN => n7787);
   U3052 : OAI22_X1 port map( A1 => n17342, A2 => n11881, B1 => n17333, B2 => 
                           n16438, ZN => n7789);
   U3053 : OAI22_X1 port map( A1 => n17368, A2 => n15669, B1 => n17359, B2 => 
                           n16438, ZN => n7790);
   U3054 : OAI22_X1 port map( A1 => n17394, A2 => n14712, B1 => n17385, B2 => 
                           n16438, ZN => n7791);
   U3055 : OAI22_X1 port map( A1 => n17058, A2 => n14363, B1 => n17049, B2 => 
                           n16443, ZN => n7852);
   U3056 : OAI22_X1 port map( A1 => n17071, A2 => n15153, B1 => n17063, B2 => 
                           n16443, ZN => n7853);
   U3057 : OAI22_X1 port map( A1 => n17110, A2 => n11756, B1 => n17101, B2 => 
                           n16443, ZN => n7854);
   U3058 : OAI22_X1 port map( A1 => n17251, A2 => n12206, B1 => n17242, B2 => 
                           n16444, ZN => n7860);
   U3059 : OAI22_X1 port map( A1 => n17264, A2 => n14832, B1 => n17256, B2 => 
                           n16444, ZN => n7861);
   U3060 : OAI22_X1 port map( A1 => n17303, A2 => n14606, B1 => n17294, B2 => 
                           n16444, ZN => n7862);
   U3061 : OAI22_X1 port map( A1 => n17355, A2 => n15074, B1 => n17346, B2 => 
                           n16444, ZN => n7864);
   U3062 : OAI22_X1 port map( A1 => n17368, A2 => n15670, B1 => n17360, B2 => 
                           n16444, ZN => n7865);
   U3063 : OAI22_X1 port map( A1 => n17407, A2 => n14330, B1 => n17398, B2 => 
                           n16444, ZN => n7866);
   U3064 : OAI22_X1 port map( A1 => n17084, A2 => n15586, B1 => n17075, B2 => 
                           n16449, ZN => n7928);
   U3065 : OAI22_X1 port map( A1 => n17097, A2 => n15497, B1 => n17089, B2 => 
                           n16449, ZN => n7929);
   U3066 : OAI22_X1 port map( A1 => n17110, A2 => n11799, B1 => n17102, B2 => 
                           n16449, ZN => n7930);
   U3067 : OAI22_X1 port map( A1 => n17290, A2 => n14364, B1 => n17282, B2 => 
                           n16450, ZN => n7937);
   U3068 : OAI22_X1 port map( A1 => n17303, A2 => n14607, B1 => n17295, B2 => 
                           n16450, ZN => n7938);
   U3069 : OAI22_X1 port map( A1 => n17381, A2 => n14430, B1 => n17372, B2 => 
                           n16450, ZN => n7940);
   U3070 : OAI22_X1 port map( A1 => n17394, A2 => n14716, B1 => n17386, B2 => 
                           n16450, ZN => n7941);
   U3071 : OAI22_X1 port map( A1 => n17407, A2 => n14331, B1 => n17399, B2 => 
                           n16450, ZN => n7942);
   U3072 : OAI22_X1 port map( A1 => n17031, A2 => n12174, B1 => n17024, B2 => 
                           n16457, ZN => n7998);
   U3073 : OAI22_X1 port map( A1 => n17044, A2 => n15038, B1 => n17037, B2 => 
                           n16457, ZN => n7999);
   U3074 : OAI22_X1 port map( A1 => n17057, A2 => n14365, B1 => n17050, B2 => 
                           n16457, ZN => n8000);
   U3075 : OAI22_X1 port map( A1 => n17070, A2 => n15154, B1 => n17062, B2 => 
                           n16457, ZN => n8001);
   U3076 : OAI22_X1 port map( A1 => n17083, A2 => n15587, B1 => n17076, B2 => 
                           n16457, ZN => n8002);
   U3077 : OAI22_X1 port map( A1 => n17096, A2 => n15498, B1 => n17088, B2 => 
                           n16457, ZN => n8003);
   U3078 : OAI22_X1 port map( A1 => n17109, A2 => n11842, B1 => n17101, B2 => 
                           n16457, ZN => n8004);
   U3079 : OAI22_X1 port map( A1 => n17237, A2 => n15374, B1 => n17230, B2 => 
                           n16458, ZN => n8007);
   U3080 : OAI22_X1 port map( A1 => n17250, A2 => n12208, B1 => n17243, B2 => 
                           n16458, ZN => n8008);
   U3081 : OAI22_X1 port map( A1 => n17263, A2 => n14834, B1 => n17255, B2 => 
                           n16458, ZN => n8009);
   U3082 : OAI22_X1 port map( A1 => n17289, A2 => n14366, B1 => n17281, B2 => 
                           n16458, ZN => n8011);
   U3083 : OAI22_X1 port map( A1 => n17302, A2 => n14608, B1 => n17294, B2 => 
                           n16458, ZN => n8012);
   U3084 : OAI22_X1 port map( A1 => n17031, A2 => n12175, B1 => n17023, B2 => 
                           n16710, ZN => n8126);
   U3085 : OAI22_X1 port map( A1 => n17044, A2 => n15039, B1 => n17036, B2 => 
                           n16710, ZN => n8127);
   U3086 : OAI22_X1 port map( A1 => n17057, A2 => n14367, B1 => n17049, B2 => 
                           n16710, ZN => n8128);
   U3087 : OAI22_X1 port map( A1 => n17070, A2 => n15155, B1 => n17063, B2 => 
                           n16710, ZN => n8129);
   U3088 : OAI22_X1 port map( A1 => n17083, A2 => n15588, B1 => n17075, B2 => 
                           n16710, ZN => n8130);
   U3089 : OAI22_X1 port map( A1 => n17096, A2 => n15499, B1 => n17089, B2 => 
                           n16710, ZN => n8131);
   U3090 : OAI22_X1 port map( A1 => n17109, A2 => n11844, B1 => n17102, B2 => 
                           n16710, ZN => n8132);
   U3091 : OAI22_X1 port map( A1 => n17328, A2 => n15295, B1 => n17321, B2 => 
                           n16711, ZN => n8142);
   U3092 : OAI22_X1 port map( A1 => n17341, A2 => n11884, B1 => n17334, B2 => 
                           n16711, ZN => n8143);
   U3093 : OAI22_X1 port map( A1 => n17354, A2 => n15078, B1 => n17347, B2 => 
                           n16711, ZN => n8144);
   U3094 : OAI22_X1 port map( A1 => n17367, A2 => n15672, B1 => n17359, B2 => 
                           n16711, ZN => n8145);
   U3095 : OAI22_X1 port map( A1 => n17380, A2 => n14432, B1 => n17373, B2 => 
                           n16711, ZN => n8146);
   U3096 : OAI22_X1 port map( A1 => n17393, A2 => n14719, B1 => n17385, B2 => 
                           n16711, ZN => n8147);
   U3097 : OAI22_X1 port map( A1 => n17406, A2 => n14332, B1 => n17398, B2 => 
                           n16711, ZN => n8148);
   U3098 : OAI22_X1 port map( A1 => n17237, A2 => n15375, B1 => n17229, B2 => 
                           n16719, ZN => n8207);
   U3099 : OAI22_X1 port map( A1 => n17250, A2 => n12209, B1 => n17242, B2 => 
                           n16719, ZN => n8208);
   U3100 : OAI22_X1 port map( A1 => n17263, A2 => n14835, B1 => n17256, B2 => 
                           n16719, ZN => n8209);
   U3101 : OAI22_X1 port map( A1 => n17289, A2 => n14368, B1 => n17282, B2 => 
                           n16719, ZN => n8211);
   U3102 : OAI22_X1 port map( A1 => n17302, A2 => n14609, B1 => n17295, B2 => 
                           n16719, ZN => n8212);
   U3103 : OAI22_X1 port map( A1 => n17328, A2 => n15296, B1 => n17320, B2 => 
                           n16720, ZN => n8214);
   U3104 : OAI22_X1 port map( A1 => n17341, A2 => n11885, B1 => n17333, B2 => 
                           n16720, ZN => n8215);
   U3105 : OAI22_X1 port map( A1 => n17354, A2 => n15080, B1 => n17346, B2 => 
                           n16720, ZN => n8216);
   U3106 : OAI22_X1 port map( A1 => n17367, A2 => n15673, B1 => n17360, B2 => 
                           n16720, ZN => n8217);
   U3107 : OAI22_X1 port map( A1 => n17380, A2 => n14434, B1 => n17372, B2 => 
                           n16720, ZN => n8218);
   U3108 : OAI22_X1 port map( A1 => n17393, A2 => n14721, B1 => n17386, B2 => 
                           n16720, ZN => n8219);
   U3109 : OAI22_X1 port map( A1 => n17406, A2 => n14333, B1 => n17399, B2 => 
                           n16720, ZN => n8220);
   U3110 : OAI22_X1 port map( A1 => n17031, A2 => n12176, B1 => n17023, B2 => 
                           n16727, ZN => n8286);
   U3111 : OAI22_X1 port map( A1 => n17044, A2 => n15040, B1 => n17036, B2 => 
                           n16727, ZN => n8287);
   U3112 : OAI22_X1 port map( A1 => n17057, A2 => n14369, B1 => n17049, B2 => 
                           n16727, ZN => n8288);
   U3113 : OAI22_X1 port map( A1 => n17083, A2 => n15589, B1 => n17075, B2 => 
                           n16727, ZN => n8290);
   U3114 : OAI22_X1 port map( A1 => n17237, A2 => n15376, B1 => n17229, B2 => 
                           n16728, ZN => n8303);
   U3115 : OAI22_X1 port map( A1 => n17250, A2 => n12210, B1 => n17242, B2 => 
                           n16728, ZN => n8304);
   U3116 : OAI22_X1 port map( A1 => n17328, A2 => n15297, B1 => n17320, B2 => 
                           n16729, ZN => n8310);
   U3117 : OAI22_X1 port map( A1 => n17341, A2 => n11886, B1 => n17333, B2 => 
                           n16729, ZN => n8311);
   U3118 : OAI22_X1 port map( A1 => n17354, A2 => n15081, B1 => n17346, B2 => 
                           n16729, ZN => n8312);
   U3119 : OAI22_X1 port map( A1 => n17380, A2 => n14435, B1 => n17372, B2 => 
                           n16729, ZN => n8314);
   U3120 : OAI22_X1 port map( A1 => n17031, A2 => n12177, B1 => n17023, B2 => 
                           n16733, ZN => n8358);
   U3121 : OAI22_X1 port map( A1 => n17328, A2 => n15298, B1 => n17320, B2 => 
                           n16735, ZN => n8382);
   U3122 : OAI22_X1 port map( A1 => n17032, A2 => n12194, B1 => n17024, B2 => 
                           n16705, ZN => n10086);
   U3123 : OAI22_X1 port map( A1 => n17045, A2 => n15041, B1 => n17037, B2 => 
                           n16705, ZN => n10087);
   U3124 : OAI22_X1 port map( A1 => n17058, A2 => n14370, B1 => n17050, B2 => 
                           n16705, ZN => n10088);
   U3125 : OAI22_X1 port map( A1 => n17071, A2 => n15156, B1 => n17062, B2 => 
                           n16705, ZN => n10089);
   U3126 : OAI22_X1 port map( A1 => n17084, A2 => n15590, B1 => n17076, B2 => 
                           n16705, ZN => n10090);
   U3127 : OAI22_X1 port map( A1 => n17097, A2 => n15517, B1 => n17088, B2 => 
                           n16705, ZN => n10091);
   U3128 : OAI22_X1 port map( A1 => n17110, A2 => n11845, B1 => n17101, B2 => 
                           n16705, ZN => n10092);
   U3129 : OAI22_X1 port map( A1 => n17238, A2 => n15377, B1 => n17230, B2 => 
                           n16704, ZN => n10103);
   U3130 : OAI22_X1 port map( A1 => n17251, A2 => n12307, B1 => n17243, B2 => 
                           n16704, ZN => n10104);
   U3131 : OAI22_X1 port map( A1 => n17264, A2 => n14853, B1 => n17255, B2 => 
                           n16704, ZN => n10105);
   U3132 : OAI22_X1 port map( A1 => n17290, A2 => n14371, B1 => n17281, B2 => 
                           n16703, ZN => n10107);
   U3133 : OAI22_X1 port map( A1 => n17303, A2 => n14627, B1 => n17294, B2 => 
                           n16704, ZN => n10108);
   U3134 : OAI22_X1 port map( A1 => n17329, A2 => n15314, B1 => n17321, B2 => 
                           n16703, ZN => n10110);
   U3135 : OAI22_X1 port map( A1 => n17342, A2 => n11903, B1 => n17334, B2 => 
                           n16703, ZN => n10111);
   U3136 : OAI22_X1 port map( A1 => n17355, A2 => n15071, B1 => n17347, B2 => 
                           n16703, ZN => n10112);
   U3137 : OAI22_X1 port map( A1 => n17368, A2 => n15691, B1 => n17359, B2 => 
                           n16703, ZN => n10113);
   U3138 : OAI22_X1 port map( A1 => n17381, A2 => n14425, B1 => n17373, B2 => 
                           n16703, ZN => n10114);
   U3139 : OAI22_X1 port map( A1 => n17394, A2 => n14756, B1 => n17385, B2 => 
                           n16703, ZN => n10115);
   U3140 : OAI22_X1 port map( A1 => n17407, A2 => n14358, B1 => n17398, B2 => 
                           n16703, ZN => n10116);
   U3141 : OAI22_X1 port map( A1 => n17585, A2 => n14286, B1 => n17577, B2 => 
                           n16448, ZN => n7911);
   U3142 : OAI22_X1 port map( A1 => n17585, A2 => n14287, B1 => n17577, B2 => 
                           n16456, ZN => n7985);
   U3143 : OAI22_X1 port map( A1 => n16699, A2 => n14963, B1 => n16692, B2 => 
                           n16709, ZN => n8055);
   U3144 : OAI22_X1 port map( A1 => n16699, A2 => n14964, B1 => n16692, B2 => 
                           n16718, ZN => n8057);
   U3145 : OAI22_X1 port map( A1 => n16699, A2 => n14965, B1 => n16692, B2 => 
                           n16731, ZN => n8061);
   U3146 : OAI22_X1 port map( A1 => n16699, A2 => n14966, B1 => n16692, B2 => 
                           n16737, ZN => n8063);
   U3147 : OAI22_X1 port map( A1 => n17584, A2 => n14071, B1 => n17577, B2 => 
                           n16709, ZN => n8113);
   U3148 : OAI22_X1 port map( A1 => n17584, A2 => n14212, B1 => n17577, B2 => 
                           n16718, ZN => n8185);
   U3149 : OAI22_X1 port map( A1 => n16942, A2 => n14550, B1 => n16935, B2 => 
                           n16709, ZN => n8118);
   U3150 : OAI22_X1 port map( A1 => n17135, A2 => n15739, B1 => n17128, B2 => 
                           n16718, ZN => n8198);
   U3151 : OAI22_X1 port map( A1 => n16942, A2 => n14551, B1 => n16934, B2 => 
                           n16726, ZN => n8278);
   U3152 : OAI22_X1 port map( A1 => n17135, A2 => n15740, B1 => n17127, B2 => 
                           n16727, ZN => n8294);
   U3153 : OAI22_X1 port map( A1 => n16942, A2 => n14552, B1 => n16935, B2 => 
                           n16733, ZN => n8350);
   U3154 : OAI22_X1 port map( A1 => n17135, A2 => n15741, B1 => n17128, B2 => 
                           n16734, ZN => n8366);
   U3155 : OAI22_X1 port map( A1 => n16943, A2 => n14546, B1 => n16934, B2 => 
                           n16706, ZN => n10078);
   U3156 : OAI22_X1 port map( A1 => n17136, A2 => n15757, B1 => n17127, B2 => 
                           n16705, ZN => n10094);
   U3157 : OAI22_X1 port map( A1 => n18025, A2 => n14573, B1 => n18017, B2 => 
                           n16436, ZN => n7769);
   U3158 : OAI22_X1 port map( A1 => n18012, A2 => n12054, B1 => n18003, B2 => 
                           n16456, ZN => n7990);
   U3159 : OAI22_X1 port map( A1 => n18025, A2 => n14572, B1 => n18016, B2 => 
                           n16456, ZN => n7991);
   U3160 : OAI22_X1 port map( A1 => n18011, A2 => n12056, B1 => n18003, B2 => 
                           n16725, ZN => n8270);
   U3161 : OAI22_X1 port map( A1 => n18024, A2 => n14574, B1 => n18016, B2 => 
                           n16725, ZN => n8271);
   U3162 : OAI22_X1 port map( A1 => n18011, A2 => n12057, B1 => n18004, B2 => 
                           n16732, ZN => n8342);
   U3163 : OAI22_X1 port map( A1 => n17852, A2 => n18026, B1 => n17836, B2 => 
                           n14280, ZN => n9990);
   U3164 : OAI22_X1 port map( A1 => n17874, A2 => n18026, B1 => n17858, B2 => 
                           n14991, ZN => n9991);
   U3165 : OAI22_X1 port map( A1 => n17896, A2 => n18026, B1 => n17880, B2 => 
                           n15316, ZN => n9992);
   U3166 : OAI22_X1 port map( A1 => n17918, A2 => n18026, B1 => n17902, B2 => 
                           n14633, ZN => n9993);
   U3167 : OAI22_X1 port map( A1 => n17939, A2 => n18026, B1 => n17923, B2 => 
                           n15315, ZN => n9994);
   U3168 : OAI22_X1 port map( A1 => n17960, A2 => n18026, B1 => n17944, B2 => 
                           n14858, ZN => n9995);
   U3169 : OAI22_X1 port map( A1 => n17981, A2 => n18026, B1 => n17965, B2 => 
                           n15033, ZN => n9996);
   U3170 : OAI22_X1 port map( A1 => n17853, A2 => n16701, B1 => n17836, B2 => 
                           n14281, ZN => n10062);
   U3171 : OAI22_X1 port map( A1 => n17875, A2 => n16701, B1 => n17858, B2 => 
                           n14992, ZN => n10063);
   U3172 : OAI22_X1 port map( A1 => n17897, A2 => n16701, B1 => n17880, B2 => 
                           n15317, ZN => n10064);
   U3173 : OAI22_X1 port map( A1 => n17919, A2 => n16701, B1 => n17902, B2 => 
                           n14634, ZN => n10065);
   U3174 : OAI22_X1 port map( A1 => n17940, A2 => n16701, B1 => n17923, B2 => 
                           n14670, ZN => n10066);
   U3175 : OAI22_X1 port map( A1 => n17961, A2 => n16701, B1 => n17944, B2 => 
                           n14859, ZN => n10067);
   U3176 : OAI22_X1 port map( A1 => n17982, A2 => n16702, B1 => n17965, B2 => 
                           n15034, ZN => n10068);
   U3177 : OAI22_X1 port map( A1 => n16698, A2 => n14967, B1 => n16691, B2 => 
                           n16743, ZN => n8065);
   U3178 : OAI22_X1 port map( A1 => n16698, A2 => n14968, B1 => n16691, B2 => 
                           n16749, ZN => n8067);
   U3179 : OAI22_X1 port map( A1 => n16698, A2 => n14969, B1 => n16691, B2 => 
                           n16755, ZN => n8069);
   U3180 : OAI22_X1 port map( A1 => n16698, A2 => n14970, B1 => n16691, B2 => 
                           n16761, ZN => n8071);
   U3181 : OAI22_X1 port map( A1 => n16697, A2 => n14971, B1 => n16691, B2 => 
                           n16767, ZN => n8073);
   U3182 : OAI22_X1 port map( A1 => n16697, A2 => n14972, B1 => n16691, B2 => 
                           n16773, ZN => n8075);
   U3183 : OAI22_X1 port map( A1 => n16697, A2 => n14973, B1 => n16691, B2 => 
                           n16779, ZN => n8077);
   U3184 : OAI22_X1 port map( A1 => n16696, A2 => n14974, B1 => n16691, B2 => 
                           n16785, ZN => n8079);
   U3185 : OAI22_X1 port map( A1 => n16696, A2 => n14975, B1 => n16691, B2 => 
                           n16791, ZN => n8081);
   U3186 : OAI22_X1 port map( A1 => n16696, A2 => n14976, B1 => n16691, B2 => 
                           n16797, ZN => n8083);
   U3187 : OAI22_X1 port map( A1 => n16696, A2 => n14977, B1 => n16691, B2 => 
                           n16803, ZN => n8085);
   U3188 : OAI22_X1 port map( A1 => n16695, A2 => n14978, B1 => n16691, B2 => 
                           n16809, ZN => n8087);
   U3189 : OAI22_X1 port map( A1 => n16697, A2 => n14979, B1 => n16691, B2 => 
                           n16827, ZN => n8093);
   U3190 : OAI22_X1 port map( A1 => n17070, A2 => n15157, B1 => n17063, B2 => 
                           n16727, ZN => n8289);
   U3191 : OAI22_X1 port map( A1 => n17096, A2 => n15500, B1 => n17089, B2 => 
                           n16727, ZN => n8291);
   U3192 : OAI22_X1 port map( A1 => n17109, A2 => n11846, B1 => n17102, B2 => 
                           n16727, ZN => n8292);
   U3193 : OAI22_X1 port map( A1 => n17263, A2 => n14836, B1 => n17256, B2 => 
                           n16728, ZN => n8305);
   U3194 : OAI22_X1 port map( A1 => n17289, A2 => n14372, B1 => n17282, B2 => 
                           n16728, ZN => n8307);
   U3195 : OAI22_X1 port map( A1 => n17302, A2 => n14610, B1 => n17295, B2 => 
                           n16728, ZN => n8308);
   U3196 : OAI22_X1 port map( A1 => n17367, A2 => n15674, B1 => n17360, B2 => 
                           n16729, ZN => n8313);
   U3197 : OAI22_X1 port map( A1 => n17393, A2 => n14723, B1 => n17386, B2 => 
                           n16729, ZN => n8315);
   U3198 : OAI22_X1 port map( A1 => n17406, A2 => n14334, B1 => n17399, B2 => 
                           n16729, ZN => n8316);
   U3199 : OAI22_X1 port map( A1 => n17471, A2 => n15527, B1 => n17464, B2 => 
                           n16729, ZN => n8321);
   U3200 : OAI22_X1 port map( A1 => n17584, A2 => n14216, B1 => n17576, B2 => 
                           n16731, ZN => n8329);
   U3201 : OAI22_X1 port map( A1 => n18024, A2 => n14575, B1 => n18017, B2 => 
                           n16732, ZN => n8343);
   U3202 : OAI22_X1 port map( A1 => n17044, A2 => n15042, B1 => n17037, B2 => 
                           n16733, ZN => n8359);
   U3203 : OAI22_X1 port map( A1 => n17057, A2 => n14373, B1 => n17050, B2 => 
                           n16733, ZN => n8360);
   U3204 : OAI22_X1 port map( A1 => n17070, A2 => n15158, B1 => n17063, B2 => 
                           n16733, ZN => n8361);
   U3205 : OAI22_X1 port map( A1 => n17083, A2 => n15591, B1 => n17076, B2 => 
                           n16734, ZN => n8362);
   U3206 : OAI22_X1 port map( A1 => n17096, A2 => n15501, B1 => n17089, B2 => 
                           n16734, ZN => n8363);
   U3207 : OAI22_X1 port map( A1 => n17109, A2 => n11847, B1 => n17102, B2 => 
                           n16734, ZN => n8364);
   U3208 : OAI22_X1 port map( A1 => n17237, A2 => n15378, B1 => n17230, B2 => 
                           n16735, ZN => n8375);
   U3209 : OAI22_X1 port map( A1 => n17250, A2 => n12211, B1 => n17243, B2 => 
                           n16735, ZN => n8376);
   U3210 : OAI22_X1 port map( A1 => n17263, A2 => n14837, B1 => n17256, B2 => 
                           n16735, ZN => n8377);
   U3211 : OAI22_X1 port map( A1 => n17289, A2 => n14374, B1 => n17282, B2 => 
                           n16735, ZN => n8379);
   U3212 : OAI22_X1 port map( A1 => n17302, A2 => n14611, B1 => n17295, B2 => 
                           n16735, ZN => n8380);
   U3213 : OAI22_X1 port map( A1 => n17341, A2 => n11887, B1 => n17334, B2 => 
                           n16735, ZN => n8383);
   U3214 : OAI22_X1 port map( A1 => n17354, A2 => n15083, B1 => n17347, B2 => 
                           n16735, ZN => n8384);
   U3215 : OAI22_X1 port map( A1 => n17367, A2 => n15675, B1 => n17360, B2 => 
                           n16735, ZN => n8385);
   U3216 : OAI22_X1 port map( A1 => n17380, A2 => n14437, B1 => n17373, B2 => 
                           n16736, ZN => n8386);
   U3217 : OAI22_X1 port map( A1 => n17393, A2 => n14725, B1 => n17386, B2 => 
                           n16736, ZN => n8387);
   U3218 : OAI22_X1 port map( A1 => n17406, A2 => n14335, B1 => n17399, B2 => 
                           n16736, ZN => n8388);
   U3219 : OAI22_X1 port map( A1 => n17444, A2 => n12369, B1 => n17438, B2 => 
                           n16736, ZN => n8391);
   U3220 : OAI22_X1 port map( A1 => n17457, A2 => n14724, B1 => n17450, B2 => 
                           n16736, ZN => n8392);
   U3221 : OAI22_X1 port map( A1 => n17470, A2 => n15528, B1 => n17464, B2 => 
                           n16736, ZN => n8393);
   U3222 : OAI22_X1 port map( A1 => n17483, A2 => n15765, B1 => n17477, B2 => 
                           n16736, ZN => n8394);
   U3223 : OAI22_X1 port map( A1 => n17496, A2 => n14783, B1 => n17490, B2 => 
                           n16736, ZN => n8395);
   U3224 : OAI22_X1 port map( A1 => n17509, A2 => n15592, B1 => n17503, B2 => 
                           n16736, ZN => n8396);
   U3225 : OAI22_X1 port map( A1 => n17584, A2 => n14219, B1 => n17576, B2 => 
                           n16737, ZN => n8401);
   U3226 : OAI22_X1 port map( A1 => n18011, A2 => n12058, B1 => n18004, B2 => 
                           n16738, ZN => n8414);
   U3227 : OAI22_X1 port map( A1 => n18024, A2 => n14576, B1 => n18017, B2 => 
                           n16738, ZN => n8415);
   U3228 : OAI22_X1 port map( A1 => n16942, A2 => n14553, B1 => n16935, B2 => 
                           n16739, ZN => n8422);
   U3229 : OAI22_X1 port map( A1 => n17030, A2 => n12178, B1 => n17024, B2 => 
                           n16739, ZN => n8430);
   U3230 : OAI22_X1 port map( A1 => n17043, A2 => n15043, B1 => n17037, B2 => 
                           n16739, ZN => n8431);
   U3231 : OAI22_X1 port map( A1 => n17056, A2 => n14375, B1 => n17050, B2 => 
                           n16739, ZN => n8432);
   U3232 : OAI22_X1 port map( A1 => n17069, A2 => n15159, B1 => n17063, B2 => 
                           n16739, ZN => n8433);
   U3233 : OAI22_X1 port map( A1 => n17082, A2 => n15593, B1 => n17076, B2 => 
                           n16740, ZN => n8434);
   U3234 : OAI22_X1 port map( A1 => n17095, A2 => n15502, B1 => n17089, B2 => 
                           n16740, ZN => n8435);
   U3235 : OAI22_X1 port map( A1 => n17108, A2 => n11849, B1 => n17102, B2 => 
                           n16740, ZN => n8436);
   U3236 : OAI22_X1 port map( A1 => n17135, A2 => n15742, B1 => n17128, B2 => 
                           n16740, ZN => n8438);
   U3237 : OAI22_X1 port map( A1 => n17236, A2 => n15379, B1 => n17230, B2 => 
                           n16741, ZN => n8447);
   U3238 : OAI22_X1 port map( A1 => n17249, A2 => n12212, B1 => n17243, B2 => 
                           n16741, ZN => n8448);
   U3239 : OAI22_X1 port map( A1 => n17262, A2 => n14838, B1 => n17256, B2 => 
                           n16741, ZN => n8449);
   U3240 : OAI22_X1 port map( A1 => n17288, A2 => n14376, B1 => n17282, B2 => 
                           n16741, ZN => n8451);
   U3241 : OAI22_X1 port map( A1 => n17301, A2 => n14612, B1 => n17295, B2 => 
                           n16741, ZN => n8452);
   U3242 : OAI22_X1 port map( A1 => n17327, A2 => n15299, B1 => n17321, B2 => 
                           n16741, ZN => n8454);
   U3243 : OAI22_X1 port map( A1 => n17340, A2 => n11888, B1 => n17334, B2 => 
                           n16741, ZN => n8455);
   U3244 : OAI22_X1 port map( A1 => n17353, A2 => n15085, B1 => n17347, B2 => 
                           n16741, ZN => n8456);
   U3245 : OAI22_X1 port map( A1 => n17366, A2 => n15676, B1 => n17360, B2 => 
                           n16741, ZN => n8457);
   U3246 : OAI22_X1 port map( A1 => n17379, A2 => n14439, B1 => n17373, B2 => 
                           n16742, ZN => n8458);
   U3247 : OAI22_X1 port map( A1 => n17392, A2 => n14727, B1 => n17386, B2 => 
                           n16742, ZN => n8459);
   U3248 : OAI22_X1 port map( A1 => n17405, A2 => n14336, B1 => n17399, B2 => 
                           n16742, ZN => n8460);
   U3249 : OAI22_X1 port map( A1 => n17431, A2 => n15334, B1 => n17425, B2 => 
                           n16742, ZN => n8462);
   U3250 : OAI22_X1 port map( A1 => n17444, A2 => n12408, B1 => n17438, B2 => 
                           n16742, ZN => n8463);
   U3251 : OAI22_X1 port map( A1 => n17457, A2 => n14726, B1 => n17450, B2 => 
                           n16742, ZN => n8464);
   U3252 : OAI22_X1 port map( A1 => n17470, A2 => n15529, B1 => n17464, B2 => 
                           n16742, ZN => n8465);
   U3253 : OAI22_X1 port map( A1 => n17483, A2 => n15766, B1 => n17477, B2 => 
                           n16742, ZN => n8466);
   U3254 : OAI22_X1 port map( A1 => n17496, A2 => n14785, B1 => n17490, B2 => 
                           n16742, ZN => n8467);
   U3255 : OAI22_X1 port map( A1 => n17509, A2 => n15594, B1 => n17503, B2 => 
                           n16742, ZN => n8468);
   U3256 : OAI22_X1 port map( A1 => n17583, A2 => n14225, B1 => n17576, B2 => 
                           n16743, ZN => n8473);
   U3257 : OAI22_X1 port map( A1 => n18011, A2 => n12059, B1 => n18004, B2 => 
                           n16744, ZN => n8486);
   U3258 : OAI22_X1 port map( A1 => n18024, A2 => n14577, B1 => n18017, B2 => 
                           n16744, ZN => n8487);
   U3259 : OAI22_X1 port map( A1 => n16941, A2 => n14554, B1 => n16935, B2 => 
                           n16745, ZN => n8494);
   U3260 : OAI22_X1 port map( A1 => n17030, A2 => n12179, B1 => n17024, B2 => 
                           n16745, ZN => n8502);
   U3261 : OAI22_X1 port map( A1 => n17043, A2 => n15044, B1 => n17037, B2 => 
                           n16745, ZN => n8503);
   U3262 : OAI22_X1 port map( A1 => n17056, A2 => n14377, B1 => n17050, B2 => 
                           n16745, ZN => n8504);
   U3263 : OAI22_X1 port map( A1 => n17069, A2 => n15160, B1 => n17063, B2 => 
                           n16745, ZN => n8505);
   U3264 : OAI22_X1 port map( A1 => n17082, A2 => n15595, B1 => n17076, B2 => 
                           n16746, ZN => n8506);
   U3265 : OAI22_X1 port map( A1 => n17095, A2 => n15503, B1 => n17089, B2 => 
                           n16746, ZN => n8507);
   U3266 : OAI22_X1 port map( A1 => n17108, A2 => n11850, B1 => n17102, B2 => 
                           n16746, ZN => n8508);
   U3267 : OAI22_X1 port map( A1 => n17134, A2 => n15743, B1 => n17128, B2 => 
                           n16746, ZN => n8510);
   U3268 : OAI22_X1 port map( A1 => n17236, A2 => n15380, B1 => n17230, B2 => 
                           n16747, ZN => n8519);
   U3269 : OAI22_X1 port map( A1 => n17249, A2 => n12213, B1 => n17243, B2 => 
                           n16747, ZN => n8520);
   U3270 : OAI22_X1 port map( A1 => n17262, A2 => n14839, B1 => n17256, B2 => 
                           n16747, ZN => n8521);
   U3271 : OAI22_X1 port map( A1 => n17288, A2 => n14378, B1 => n17282, B2 => 
                           n16747, ZN => n8523);
   U3272 : OAI22_X1 port map( A1 => n17301, A2 => n14613, B1 => n17295, B2 => 
                           n16747, ZN => n8524);
   U3273 : OAI22_X1 port map( A1 => n17327, A2 => n15300, B1 => n17321, B2 => 
                           n16747, ZN => n8526);
   U3274 : OAI22_X1 port map( A1 => n17340, A2 => n11889, B1 => n17334, B2 => 
                           n16747, ZN => n8527);
   U3275 : OAI22_X1 port map( A1 => n17353, A2 => n15087, B1 => n17347, B2 => 
                           n16747, ZN => n8528);
   U3276 : OAI22_X1 port map( A1 => n17366, A2 => n15677, B1 => n17360, B2 => 
                           n16747, ZN => n8529);
   U3277 : OAI22_X1 port map( A1 => n17379, A2 => n14441, B1 => n17373, B2 => 
                           n16748, ZN => n8530);
   U3278 : OAI22_X1 port map( A1 => n17392, A2 => n14729, B1 => n17386, B2 => 
                           n16748, ZN => n8531);
   U3279 : OAI22_X1 port map( A1 => n17405, A2 => n14337, B1 => n17399, B2 => 
                           n16748, ZN => n8532);
   U3280 : OAI22_X1 port map( A1 => n17431, A2 => n15335, B1 => n17425, B2 => 
                           n16748, ZN => n8534);
   U3281 : OAI22_X1 port map( A1 => n17444, A2 => n12410, B1 => n17438, B2 => 
                           n16748, ZN => n8535);
   U3282 : OAI22_X1 port map( A1 => n17457, A2 => n14728, B1 => n17450, B2 => 
                           n16748, ZN => n8536);
   U3283 : OAI22_X1 port map( A1 => n17470, A2 => n15530, B1 => n17464, B2 => 
                           n16748, ZN => n8537);
   U3284 : OAI22_X1 port map( A1 => n17483, A2 => n15767, B1 => n17477, B2 => 
                           n16748, ZN => n8538);
   U3285 : OAI22_X1 port map( A1 => n17496, A2 => n14787, B1 => n17490, B2 => 
                           n16748, ZN => n8539);
   U3286 : OAI22_X1 port map( A1 => n17509, A2 => n15596, B1 => n17503, B2 => 
                           n16748, ZN => n8540);
   U3287 : OAI22_X1 port map( A1 => n17583, A2 => n14227, B1 => n17576, B2 => 
                           n16749, ZN => n8545);
   U3288 : OAI22_X1 port map( A1 => n18010, A2 => n12060, B1 => n18004, B2 => 
                           n16750, ZN => n8558);
   U3289 : OAI22_X1 port map( A1 => n18023, A2 => n14578, B1 => n18017, B2 => 
                           n16750, ZN => n8559);
   U3290 : OAI22_X1 port map( A1 => n16941, A2 => n14555, B1 => n16935, B2 => 
                           n16751, ZN => n8566);
   U3291 : OAI22_X1 port map( A1 => n17030, A2 => n12180, B1 => n17024, B2 => 
                           n16751, ZN => n8574);
   U3292 : OAI22_X1 port map( A1 => n17043, A2 => n15045, B1 => n17037, B2 => 
                           n16751, ZN => n8575);
   U3293 : OAI22_X1 port map( A1 => n17056, A2 => n14379, B1 => n17050, B2 => 
                           n16751, ZN => n8576);
   U3294 : OAI22_X1 port map( A1 => n17069, A2 => n15161, B1 => n17063, B2 => 
                           n16751, ZN => n8577);
   U3295 : OAI22_X1 port map( A1 => n17082, A2 => n15597, B1 => n17076, B2 => 
                           n16752, ZN => n8578);
   U3296 : OAI22_X1 port map( A1 => n17095, A2 => n15504, B1 => n17089, B2 => 
                           n16752, ZN => n8579);
   U3297 : OAI22_X1 port map( A1 => n17108, A2 => n11851, B1 => n17102, B2 => 
                           n16752, ZN => n8580);
   U3298 : OAI22_X1 port map( A1 => n17134, A2 => n15744, B1 => n17128, B2 => 
                           n16752, ZN => n8582);
   U3299 : OAI22_X1 port map( A1 => n17236, A2 => n15381, B1 => n17230, B2 => 
                           n16753, ZN => n8591);
   U3300 : OAI22_X1 port map( A1 => n17249, A2 => n12214, B1 => n17243, B2 => 
                           n16753, ZN => n8592);
   U3301 : OAI22_X1 port map( A1 => n17262, A2 => n14840, B1 => n17256, B2 => 
                           n16753, ZN => n8593);
   U3302 : OAI22_X1 port map( A1 => n17288, A2 => n14380, B1 => n17282, B2 => 
                           n16753, ZN => n8595);
   U3303 : OAI22_X1 port map( A1 => n17301, A2 => n14614, B1 => n17295, B2 => 
                           n16753, ZN => n8596);
   U3304 : OAI22_X1 port map( A1 => n17327, A2 => n15301, B1 => n17321, B2 => 
                           n16753, ZN => n8598);
   U3305 : OAI22_X1 port map( A1 => n17340, A2 => n11890, B1 => n17334, B2 => 
                           n16753, ZN => n8599);
   U3306 : OAI22_X1 port map( A1 => n17353, A2 => n15089, B1 => n17347, B2 => 
                           n16753, ZN => n8600);
   U3307 : OAI22_X1 port map( A1 => n17366, A2 => n15678, B1 => n17360, B2 => 
                           n16753, ZN => n8601);
   U3308 : OAI22_X1 port map( A1 => n17379, A2 => n14443, B1 => n17373, B2 => 
                           n16754, ZN => n8602);
   U3309 : OAI22_X1 port map( A1 => n17392, A2 => n14731, B1 => n17386, B2 => 
                           n16754, ZN => n8603);
   U3310 : OAI22_X1 port map( A1 => n17405, A2 => n14338, B1 => n17399, B2 => 
                           n16754, ZN => n8604);
   U3311 : OAI22_X1 port map( A1 => n17431, A2 => n15336, B1 => n17425, B2 => 
                           n16754, ZN => n8606);
   U3312 : OAI22_X1 port map( A1 => n17444, A2 => n12551, B1 => n17438, B2 => 
                           n16754, ZN => n8607);
   U3313 : OAI22_X1 port map( A1 => n17457, A2 => n14730, B1 => n17450, B2 => 
                           n16754, ZN => n8608);
   U3314 : OAI22_X1 port map( A1 => n17470, A2 => n15531, B1 => n17464, B2 => 
                           n16754, ZN => n8609);
   U3315 : OAI22_X1 port map( A1 => n17483, A2 => n15768, B1 => n17477, B2 => 
                           n16754, ZN => n8610);
   U3316 : OAI22_X1 port map( A1 => n17496, A2 => n14789, B1 => n17490, B2 => 
                           n16754, ZN => n8611);
   U3317 : OAI22_X1 port map( A1 => n17509, A2 => n15598, B1 => n17503, B2 => 
                           n16754, ZN => n8612);
   U3318 : OAI22_X1 port map( A1 => n17583, A2 => n14230, B1 => n17576, B2 => 
                           n16755, ZN => n8617);
   U3319 : OAI22_X1 port map( A1 => n18010, A2 => n12098, B1 => n18004, B2 => 
                           n16756, ZN => n8630);
   U3320 : OAI22_X1 port map( A1 => n18023, A2 => n14579, B1 => n18017, B2 => 
                           n16756, ZN => n8631);
   U3321 : OAI22_X1 port map( A1 => n16941, A2 => n14556, B1 => n16935, B2 => 
                           n16757, ZN => n8638);
   U3322 : OAI22_X1 port map( A1 => n17030, A2 => n12181, B1 => n17024, B2 => 
                           n16757, ZN => n8646);
   U3323 : OAI22_X1 port map( A1 => n17043, A2 => n15046, B1 => n17037, B2 => 
                           n16757, ZN => n8647);
   U3324 : OAI22_X1 port map( A1 => n17056, A2 => n14381, B1 => n17050, B2 => 
                           n16757, ZN => n8648);
   U3325 : OAI22_X1 port map( A1 => n17069, A2 => n15162, B1 => n17063, B2 => 
                           n16757, ZN => n8649);
   U3326 : OAI22_X1 port map( A1 => n17082, A2 => n15599, B1 => n17076, B2 => 
                           n16758, ZN => n8650);
   U3327 : OAI22_X1 port map( A1 => n17095, A2 => n15505, B1 => n17089, B2 => 
                           n16758, ZN => n8651);
   U3328 : OAI22_X1 port map( A1 => n17108, A2 => n11852, B1 => n17102, B2 => 
                           n16758, ZN => n8652);
   U3329 : OAI22_X1 port map( A1 => n17134, A2 => n15745, B1 => n17128, B2 => 
                           n16758, ZN => n8654);
   U3330 : OAI22_X1 port map( A1 => n17236, A2 => n15382, B1 => n17230, B2 => 
                           n16759, ZN => n8663);
   U3331 : OAI22_X1 port map( A1 => n17249, A2 => n12215, B1 => n17243, B2 => 
                           n16759, ZN => n8664);
   U3332 : OAI22_X1 port map( A1 => n17262, A2 => n14841, B1 => n17256, B2 => 
                           n16759, ZN => n8665);
   U3333 : OAI22_X1 port map( A1 => n17288, A2 => n14382, B1 => n17282, B2 => 
                           n16759, ZN => n8667);
   U3334 : OAI22_X1 port map( A1 => n17301, A2 => n14615, B1 => n17295, B2 => 
                           n16759, ZN => n8668);
   U3335 : OAI22_X1 port map( A1 => n17327, A2 => n15302, B1 => n17321, B2 => 
                           n16759, ZN => n8670);
   U3336 : OAI22_X1 port map( A1 => n17340, A2 => n11891, B1 => n17334, B2 => 
                           n16759, ZN => n8671);
   U3337 : OAI22_X1 port map( A1 => n17353, A2 => n15091, B1 => n17347, B2 => 
                           n16759, ZN => n8672);
   U3338 : OAI22_X1 port map( A1 => n17366, A2 => n15679, B1 => n17360, B2 => 
                           n16759, ZN => n8673);
   U3339 : OAI22_X1 port map( A1 => n17379, A2 => n14445, B1 => n17373, B2 => 
                           n16760, ZN => n8674);
   U3340 : OAI22_X1 port map( A1 => n17392, A2 => n14733, B1 => n17386, B2 => 
                           n16760, ZN => n8675);
   U3341 : OAI22_X1 port map( A1 => n17405, A2 => n14339, B1 => n17399, B2 => 
                           n16760, ZN => n8676);
   U3342 : OAI22_X1 port map( A1 => n17430, A2 => n15337, B1 => n17425, B2 => 
                           n16760, ZN => n8678);
   U3343 : OAI22_X1 port map( A1 => n17443, A2 => n12602, B1 => n17438, B2 => 
                           n16760, ZN => n8679);
   U3344 : OAI22_X1 port map( A1 => n17456, A2 => n14732, B1 => n17450, B2 => 
                           n16760, ZN => n8680);
   U3345 : OAI22_X1 port map( A1 => n17469, A2 => n15532, B1 => n17464, B2 => 
                           n16760, ZN => n8681);
   U3346 : OAI22_X1 port map( A1 => n17482, A2 => n15769, B1 => n17477, B2 => 
                           n16760, ZN => n8682);
   U3347 : OAI22_X1 port map( A1 => n17495, A2 => n14791, B1 => n17490, B2 => 
                           n16760, ZN => n8683);
   U3348 : OAI22_X1 port map( A1 => n17508, A2 => n15600, B1 => n17503, B2 => 
                           n16760, ZN => n8684);
   U3349 : OAI22_X1 port map( A1 => n17583, A2 => n14235, B1 => n17576, B2 => 
                           n16761, ZN => n8689);
   U3350 : OAI22_X1 port map( A1 => n18010, A2 => n12099, B1 => n18004, B2 => 
                           n16762, ZN => n8702);
   U3351 : OAI22_X1 port map( A1 => n18023, A2 => n14580, B1 => n18017, B2 => 
                           n16762, ZN => n8703);
   U3352 : OAI22_X1 port map( A1 => n16941, A2 => n14557, B1 => n16935, B2 => 
                           n16763, ZN => n8710);
   U3353 : OAI22_X1 port map( A1 => n17029, A2 => n12182, B1 => n17024, B2 => 
                           n16763, ZN => n8718);
   U3354 : OAI22_X1 port map( A1 => n17042, A2 => n15047, B1 => n17037, B2 => 
                           n16763, ZN => n8719);
   U3355 : OAI22_X1 port map( A1 => n17055, A2 => n14383, B1 => n17050, B2 => 
                           n16763, ZN => n8720);
   U3356 : OAI22_X1 port map( A1 => n17068, A2 => n15163, B1 => n17063, B2 => 
                           n16763, ZN => n8721);
   U3357 : OAI22_X1 port map( A1 => n17081, A2 => n15601, B1 => n17076, B2 => 
                           n16764, ZN => n8722);
   U3358 : OAI22_X1 port map( A1 => n17094, A2 => n15506, B1 => n17089, B2 => 
                           n16764, ZN => n8723);
   U3359 : OAI22_X1 port map( A1 => n17107, A2 => n11854, B1 => n17102, B2 => 
                           n16764, ZN => n8724);
   U3360 : OAI22_X1 port map( A1 => n17134, A2 => n15746, B1 => n17128, B2 => 
                           n16764, ZN => n8726);
   U3361 : OAI22_X1 port map( A1 => n17235, A2 => n15383, B1 => n17230, B2 => 
                           n16765, ZN => n8735);
   U3362 : OAI22_X1 port map( A1 => n17248, A2 => n12253, B1 => n17243, B2 => 
                           n16765, ZN => n8736);
   U3363 : OAI22_X1 port map( A1 => n17261, A2 => n14842, B1 => n17256, B2 => 
                           n16765, ZN => n8737);
   U3364 : OAI22_X1 port map( A1 => n17287, A2 => n14384, B1 => n17282, B2 => 
                           n16765, ZN => n8739);
   U3365 : OAI22_X1 port map( A1 => n17300, A2 => n14616, B1 => n17295, B2 => 
                           n16765, ZN => n8740);
   U3366 : OAI22_X1 port map( A1 => n17326, A2 => n15303, B1 => n17321, B2 => 
                           n16765, ZN => n8742);
   U3367 : OAI22_X1 port map( A1 => n17339, A2 => n11892, B1 => n17334, B2 => 
                           n16765, ZN => n8743);
   U3368 : OAI22_X1 port map( A1 => n17352, A2 => n15093, B1 => n17347, B2 => 
                           n16765, ZN => n8744);
   U3369 : OAI22_X1 port map( A1 => n17365, A2 => n15680, B1 => n17360, B2 => 
                           n16765, ZN => n8745);
   U3370 : OAI22_X1 port map( A1 => n17378, A2 => n14447, B1 => n17373, B2 => 
                           n16766, ZN => n8746);
   U3371 : OAI22_X1 port map( A1 => n17391, A2 => n14735, B1 => n17386, B2 => 
                           n16766, ZN => n8747);
   U3372 : OAI22_X1 port map( A1 => n17404, A2 => n14340, B1 => n17399, B2 => 
                           n16766, ZN => n8748);
   U3373 : OAI22_X1 port map( A1 => n17430, A2 => n15338, B1 => n17425, B2 => 
                           n16766, ZN => n8750);
   U3374 : OAI22_X1 port map( A1 => n17443, A2 => n12669, B1 => n17438, B2 => 
                           n16766, ZN => n8751);
   U3375 : OAI22_X1 port map( A1 => n17456, A2 => n14734, B1 => n17450, B2 => 
                           n16766, ZN => n8752);
   U3376 : OAI22_X1 port map( A1 => n17469, A2 => n15533, B1 => n17464, B2 => 
                           n16766, ZN => n8753);
   U3377 : OAI22_X1 port map( A1 => n17482, A2 => n15770, B1 => n17477, B2 => 
                           n16766, ZN => n8754);
   U3378 : OAI22_X1 port map( A1 => n17495, A2 => n14793, B1 => n17490, B2 => 
                           n16766, ZN => n8755);
   U3379 : OAI22_X1 port map( A1 => n17508, A2 => n15602, B1 => n17503, B2 => 
                           n16766, ZN => n8756);
   U3380 : OAI22_X1 port map( A1 => n17582, A2 => n14242, B1 => n17576, B2 => 
                           n16767, ZN => n8761);
   U3381 : OAI22_X1 port map( A1 => n18010, A2 => n12100, B1 => n18004, B2 => 
                           n16768, ZN => n8774);
   U3382 : OAI22_X1 port map( A1 => n18023, A2 => n14581, B1 => n18017, B2 => 
                           n16768, ZN => n8775);
   U3383 : OAI22_X1 port map( A1 => n16940, A2 => n14558, B1 => n16935, B2 => 
                           n16769, ZN => n8782);
   U3384 : OAI22_X1 port map( A1 => n17029, A2 => n12183, B1 => n17024, B2 => 
                           n16769, ZN => n8790);
   U3385 : OAI22_X1 port map( A1 => n17042, A2 => n15048, B1 => n17037, B2 => 
                           n16769, ZN => n8791);
   U3386 : OAI22_X1 port map( A1 => n17055, A2 => n14385, B1 => n17050, B2 => 
                           n16769, ZN => n8792);
   U3387 : OAI22_X1 port map( A1 => n17068, A2 => n15164, B1 => n17063, B2 => 
                           n16769, ZN => n8793);
   U3388 : OAI22_X1 port map( A1 => n17081, A2 => n15603, B1 => n17076, B2 => 
                           n16770, ZN => n8794);
   U3389 : OAI22_X1 port map( A1 => n17094, A2 => n15507, B1 => n17089, B2 => 
                           n16770, ZN => n8795);
   U3390 : OAI22_X1 port map( A1 => n17107, A2 => n11855, B1 => n17102, B2 => 
                           n16770, ZN => n8796);
   U3391 : OAI22_X1 port map( A1 => n17133, A2 => n15747, B1 => n17128, B2 => 
                           n16770, ZN => n8798);
   U3392 : OAI22_X1 port map( A1 => n17235, A2 => n15384, B1 => n17230, B2 => 
                           n16771, ZN => n8807);
   U3393 : OAI22_X1 port map( A1 => n17248, A2 => n12254, B1 => n17243, B2 => 
                           n16771, ZN => n8808);
   U3394 : OAI22_X1 port map( A1 => n17261, A2 => n14843, B1 => n17256, B2 => 
                           n16771, ZN => n8809);
   U3395 : OAI22_X1 port map( A1 => n17287, A2 => n14386, B1 => n17282, B2 => 
                           n16771, ZN => n8811);
   U3396 : OAI22_X1 port map( A1 => n17300, A2 => n14617, B1 => n17295, B2 => 
                           n16771, ZN => n8812);
   U3397 : OAI22_X1 port map( A1 => n17326, A2 => n15304, B1 => n17321, B2 => 
                           n16771, ZN => n8814);
   U3398 : OAI22_X1 port map( A1 => n17339, A2 => n11893, B1 => n17334, B2 => 
                           n16771, ZN => n8815);
   U3399 : OAI22_X1 port map( A1 => n17352, A2 => n15095, B1 => n17347, B2 => 
                           n16771, ZN => n8816);
   U3400 : OAI22_X1 port map( A1 => n17365, A2 => n15681, B1 => n17360, B2 => 
                           n16771, ZN => n8817);
   U3401 : OAI22_X1 port map( A1 => n17378, A2 => n14449, B1 => n17373, B2 => 
                           n16772, ZN => n8818);
   U3402 : OAI22_X1 port map( A1 => n17391, A2 => n14737, B1 => n17386, B2 => 
                           n16772, ZN => n8819);
   U3403 : OAI22_X1 port map( A1 => n17404, A2 => n14341, B1 => n17399, B2 => 
                           n16772, ZN => n8820);
   U3404 : OAI22_X1 port map( A1 => n17430, A2 => n15339, B1 => n17425, B2 => 
                           n16772, ZN => n8822);
   U3405 : OAI22_X1 port map( A1 => n17443, A2 => n13999, B1 => n17438, B2 => 
                           n16772, ZN => n8823);
   U3406 : OAI22_X1 port map( A1 => n17456, A2 => n14736, B1 => n17450, B2 => 
                           n16772, ZN => n8824);
   U3407 : OAI22_X1 port map( A1 => n17469, A2 => n15534, B1 => n17464, B2 => 
                           n16772, ZN => n8825);
   U3408 : OAI22_X1 port map( A1 => n17482, A2 => n15771, B1 => n17477, B2 => 
                           n16772, ZN => n8826);
   U3409 : OAI22_X1 port map( A1 => n17495, A2 => n14795, B1 => n17490, B2 => 
                           n16772, ZN => n8827);
   U3410 : OAI22_X1 port map( A1 => n17508, A2 => n15604, B1 => n17503, B2 => 
                           n16772, ZN => n8828);
   U3411 : OAI22_X1 port map( A1 => n17582, A2 => n14243, B1 => n17576, B2 => 
                           n16773, ZN => n8833);
   U3412 : OAI22_X1 port map( A1 => n18009, A2 => n12101, B1 => n18004, B2 => 
                           n16774, ZN => n8846);
   U3413 : OAI22_X1 port map( A1 => n18022, A2 => n14582, B1 => n18017, B2 => 
                           n16774, ZN => n8847);
   U3414 : OAI22_X1 port map( A1 => n16940, A2 => n14559, B1 => n16935, B2 => 
                           n16775, ZN => n8854);
   U3415 : OAI22_X1 port map( A1 => n17029, A2 => n12185, B1 => n17024, B2 => 
                           n16775, ZN => n8862);
   U3416 : OAI22_X1 port map( A1 => n17042, A2 => n15049, B1 => n17037, B2 => 
                           n16775, ZN => n8863);
   U3417 : OAI22_X1 port map( A1 => n17055, A2 => n14387, B1 => n17050, B2 => 
                           n16775, ZN => n8864);
   U3418 : OAI22_X1 port map( A1 => n17068, A2 => n15165, B1 => n17063, B2 => 
                           n16775, ZN => n8865);
   U3419 : OAI22_X1 port map( A1 => n17081, A2 => n15605, B1 => n17076, B2 => 
                           n16776, ZN => n8866);
   U3420 : OAI22_X1 port map( A1 => n17094, A2 => n15508, B1 => n17089, B2 => 
                           n16776, ZN => n8867);
   U3421 : OAI22_X1 port map( A1 => n17107, A2 => n11856, B1 => n17102, B2 => 
                           n16776, ZN => n8868);
   U3422 : OAI22_X1 port map( A1 => n17133, A2 => n15748, B1 => n17128, B2 => 
                           n16776, ZN => n8870);
   U3423 : OAI22_X1 port map( A1 => n17235, A2 => n15385, B1 => n17230, B2 => 
                           n16777, ZN => n8879);
   U3424 : OAI22_X1 port map( A1 => n17248, A2 => n12255, B1 => n17243, B2 => 
                           n16777, ZN => n8880);
   U3425 : OAI22_X1 port map( A1 => n17261, A2 => n14844, B1 => n17256, B2 => 
                           n16777, ZN => n8881);
   U3426 : OAI22_X1 port map( A1 => n17287, A2 => n14388, B1 => n17282, B2 => 
                           n16777, ZN => n8883);
   U3427 : OAI22_X1 port map( A1 => n17300, A2 => n14618, B1 => n17295, B2 => 
                           n16777, ZN => n8884);
   U3428 : OAI22_X1 port map( A1 => n17326, A2 => n15305, B1 => n17321, B2 => 
                           n16777, ZN => n8886);
   U3429 : OAI22_X1 port map( A1 => n17339, A2 => n11894, B1 => n17334, B2 => 
                           n16777, ZN => n8887);
   U3430 : OAI22_X1 port map( A1 => n17352, A2 => n15097, B1 => n17347, B2 => 
                           n16777, ZN => n8888);
   U3431 : OAI22_X1 port map( A1 => n17365, A2 => n15682, B1 => n17360, B2 => 
                           n16777, ZN => n8889);
   U3432 : OAI22_X1 port map( A1 => n17378, A2 => n14451, B1 => n17373, B2 => 
                           n16778, ZN => n8890);
   U3433 : OAI22_X1 port map( A1 => n17391, A2 => n14739, B1 => n17386, B2 => 
                           n16778, ZN => n8891);
   U3434 : OAI22_X1 port map( A1 => n17404, A2 => n14342, B1 => n17399, B2 => 
                           n16778, ZN => n8892);
   U3435 : OAI22_X1 port map( A1 => n17429, A2 => n15340, B1 => n17425, B2 => 
                           n16778, ZN => n8894);
   U3436 : OAI22_X1 port map( A1 => n17442, A2 => n14014, B1 => n17438, B2 => 
                           n16778, ZN => n8895);
   U3437 : OAI22_X1 port map( A1 => n17455, A2 => n14738, B1 => n17450, B2 => 
                           n16778, ZN => n8896);
   U3438 : OAI22_X1 port map( A1 => n17468, A2 => n15535, B1 => n17464, B2 => 
                           n16778, ZN => n8897);
   U3439 : OAI22_X1 port map( A1 => n17481, A2 => n15772, B1 => n17477, B2 => 
                           n16778, ZN => n8898);
   U3440 : OAI22_X1 port map( A1 => n17494, A2 => n14797, B1 => n17490, B2 => 
                           n16778, ZN => n8899);
   U3441 : OAI22_X1 port map( A1 => n17507, A2 => n15606, B1 => n17503, B2 => 
                           n16778, ZN => n8900);
   U3442 : OAI22_X1 port map( A1 => n17582, A2 => n14246, B1 => n17576, B2 => 
                           n16779, ZN => n8905);
   U3443 : OAI22_X1 port map( A1 => n18009, A2 => n12102, B1 => n18004, B2 => 
                           n16780, ZN => n8918);
   U3444 : OAI22_X1 port map( A1 => n18022, A2 => n14583, B1 => n18017, B2 => 
                           n16780, ZN => n8919);
   U3445 : OAI22_X1 port map( A1 => n16940, A2 => n14560, B1 => n16935, B2 => 
                           n16781, ZN => n8926);
   U3446 : OAI22_X1 port map( A1 => n17028, A2 => n12186, B1 => n17024, B2 => 
                           n16781, ZN => n8934);
   U3447 : OAI22_X1 port map( A1 => n17041, A2 => n15050, B1 => n17037, B2 => 
                           n16781, ZN => n8935);
   U3448 : OAI22_X1 port map( A1 => n17054, A2 => n14389, B1 => n17050, B2 => 
                           n16781, ZN => n8936);
   U3449 : OAI22_X1 port map( A1 => n17067, A2 => n15166, B1 => n17063, B2 => 
                           n16781, ZN => n8937);
   U3450 : OAI22_X1 port map( A1 => n17080, A2 => n15607, B1 => n17076, B2 => 
                           n16782, ZN => n8938);
   U3451 : OAI22_X1 port map( A1 => n17093, A2 => n15509, B1 => n17089, B2 => 
                           n16782, ZN => n8939);
   U3452 : OAI22_X1 port map( A1 => n17106, A2 => n11857, B1 => n17102, B2 => 
                           n16782, ZN => n8940);
   U3453 : OAI22_X1 port map( A1 => n17133, A2 => n15749, B1 => n17128, B2 => 
                           n16782, ZN => n8942);
   U3454 : OAI22_X1 port map( A1 => n17234, A2 => n15386, B1 => n17230, B2 => 
                           n16783, ZN => n8951);
   U3455 : OAI22_X1 port map( A1 => n17247, A2 => n12256, B1 => n17243, B2 => 
                           n16783, ZN => n8952);
   U3456 : OAI22_X1 port map( A1 => n17260, A2 => n14845, B1 => n17256, B2 => 
                           n16783, ZN => n8953);
   U3457 : OAI22_X1 port map( A1 => n17286, A2 => n14390, B1 => n17282, B2 => 
                           n16783, ZN => n8955);
   U3458 : OAI22_X1 port map( A1 => n17299, A2 => n14619, B1 => n17295, B2 => 
                           n16783, ZN => n8956);
   U3459 : OAI22_X1 port map( A1 => n17325, A2 => n15306, B1 => n17321, B2 => 
                           n16783, ZN => n8958);
   U3460 : OAI22_X1 port map( A1 => n17338, A2 => n11895, B1 => n17334, B2 => 
                           n16783, ZN => n8959);
   U3461 : OAI22_X1 port map( A1 => n17351, A2 => n15099, B1 => n17347, B2 => 
                           n16783, ZN => n8960);
   U3462 : OAI22_X1 port map( A1 => n17364, A2 => n15683, B1 => n17360, B2 => 
                           n16783, ZN => n8961);
   U3463 : OAI22_X1 port map( A1 => n17377, A2 => n14453, B1 => n17373, B2 => 
                           n16784, ZN => n8962);
   U3464 : OAI22_X1 port map( A1 => n17390, A2 => n14741, B1 => n17386, B2 => 
                           n16784, ZN => n8963);
   U3465 : OAI22_X1 port map( A1 => n17403, A2 => n14343, B1 => n17399, B2 => 
                           n16784, ZN => n8964);
   U3466 : OAI22_X1 port map( A1 => n17429, A2 => n15341, B1 => n17425, B2 => 
                           n16784, ZN => n8966);
   U3467 : OAI22_X1 port map( A1 => n17442, A2 => n14032, B1 => n17438, B2 => 
                           n16784, ZN => n8967);
   U3468 : OAI22_X1 port map( A1 => n17455, A2 => n14740, B1 => n17450, B2 => 
                           n16784, ZN => n8968);
   U3469 : OAI22_X1 port map( A1 => n17468, A2 => n15536, B1 => n17464, B2 => 
                           n16784, ZN => n8969);
   U3470 : OAI22_X1 port map( A1 => n17481, A2 => n15773, B1 => n17477, B2 => 
                           n16784, ZN => n8970);
   U3471 : OAI22_X1 port map( A1 => n17494, A2 => n14799, B1 => n17490, B2 => 
                           n16784, ZN => n8971);
   U3472 : OAI22_X1 port map( A1 => n17507, A2 => n15608, B1 => n17503, B2 => 
                           n16784, ZN => n8972);
   U3473 : OAI22_X1 port map( A1 => n17581, A2 => n14255, B1 => n17576, B2 => 
                           n16785, ZN => n8977);
   U3474 : OAI22_X1 port map( A1 => n18009, A2 => n12103, B1 => n18004, B2 => 
                           n16786, ZN => n8990);
   U3475 : OAI22_X1 port map( A1 => n18022, A2 => n14584, B1 => n18017, B2 => 
                           n16786, ZN => n8991);
   U3476 : OAI22_X1 port map( A1 => n16939, A2 => n14561, B1 => n16935, B2 => 
                           n16787, ZN => n8998);
   U3477 : OAI22_X1 port map( A1 => n17028, A2 => n12187, B1 => n17024, B2 => 
                           n16787, ZN => n9006);
   U3478 : OAI22_X1 port map( A1 => n17041, A2 => n15051, B1 => n17037, B2 => 
                           n16787, ZN => n9007);
   U3479 : OAI22_X1 port map( A1 => n17054, A2 => n14391, B1 => n17050, B2 => 
                           n16787, ZN => n9008);
   U3480 : OAI22_X1 port map( A1 => n17067, A2 => n15167, B1 => n17063, B2 => 
                           n16787, ZN => n9009);
   U3481 : OAI22_X1 port map( A1 => n17080, A2 => n15609, B1 => n17076, B2 => 
                           n16788, ZN => n9010);
   U3482 : OAI22_X1 port map( A1 => n17093, A2 => n15510, B1 => n17089, B2 => 
                           n16788, ZN => n9011);
   U3483 : OAI22_X1 port map( A1 => n17106, A2 => n11858, B1 => n17102, B2 => 
                           n16788, ZN => n9012);
   U3484 : OAI22_X1 port map( A1 => n17132, A2 => n15750, B1 => n17128, B2 => 
                           n16788, ZN => n9014);
   U3485 : OAI22_X1 port map( A1 => n17234, A2 => n15387, B1 => n17230, B2 => 
                           n16789, ZN => n9023);
   U3486 : OAI22_X1 port map( A1 => n17247, A2 => n12257, B1 => n17243, B2 => 
                           n16789, ZN => n9024);
   U3487 : OAI22_X1 port map( A1 => n17260, A2 => n14846, B1 => n17256, B2 => 
                           n16789, ZN => n9025);
   U3488 : OAI22_X1 port map( A1 => n17286, A2 => n14392, B1 => n17282, B2 => 
                           n16789, ZN => n9027);
   U3489 : OAI22_X1 port map( A1 => n17299, A2 => n14620, B1 => n17295, B2 => 
                           n16789, ZN => n9028);
   U3490 : OAI22_X1 port map( A1 => n17325, A2 => n15307, B1 => n17321, B2 => 
                           n16789, ZN => n9030);
   U3491 : OAI22_X1 port map( A1 => n17338, A2 => n11896, B1 => n17334, B2 => 
                           n16789, ZN => n9031);
   U3492 : OAI22_X1 port map( A1 => n17351, A2 => n15101, B1 => n17347, B2 => 
                           n16789, ZN => n9032);
   U3493 : OAI22_X1 port map( A1 => n17364, A2 => n15684, B1 => n17360, B2 => 
                           n16789, ZN => n9033);
   U3494 : OAI22_X1 port map( A1 => n17377, A2 => n14455, B1 => n17373, B2 => 
                           n16790, ZN => n9034);
   U3495 : OAI22_X1 port map( A1 => n17390, A2 => n14743, B1 => n17386, B2 => 
                           n16790, ZN => n9035);
   U3496 : OAI22_X1 port map( A1 => n17403, A2 => n14344, B1 => n17399, B2 => 
                           n16790, ZN => n9036);
   U3497 : OAI22_X1 port map( A1 => n17429, A2 => n15342, B1 => n17425, B2 => 
                           n16790, ZN => n9038);
   U3498 : OAI22_X1 port map( A1 => n17442, A2 => n14036, B1 => n17438, B2 => 
                           n16790, ZN => n9039);
   U3499 : OAI22_X1 port map( A1 => n17455, A2 => n14742, B1 => n17450, B2 => 
                           n16790, ZN => n9040);
   U3500 : OAI22_X1 port map( A1 => n17468, A2 => n15537, B1 => n17464, B2 => 
                           n16790, ZN => n9041);
   U3501 : OAI22_X1 port map( A1 => n17481, A2 => n15774, B1 => n17477, B2 => 
                           n16790, ZN => n9042);
   U3502 : OAI22_X1 port map( A1 => n17494, A2 => n14801, B1 => n17490, B2 => 
                           n16790, ZN => n9043);
   U3503 : OAI22_X1 port map( A1 => n17507, A2 => n15610, B1 => n17503, B2 => 
                           n16790, ZN => n9044);
   U3504 : OAI22_X1 port map( A1 => n17581, A2 => n14261, B1 => n17576, B2 => 
                           n16791, ZN => n9049);
   U3505 : OAI22_X1 port map( A1 => n18008, A2 => n12104, B1 => n18004, B2 => 
                           n16792, ZN => n9062);
   U3506 : OAI22_X1 port map( A1 => n18021, A2 => n14585, B1 => n18017, B2 => 
                           n16792, ZN => n9063);
   U3507 : OAI22_X1 port map( A1 => n16939, A2 => n14562, B1 => n16935, B2 => 
                           n16793, ZN => n9070);
   U3508 : OAI22_X1 port map( A1 => n17028, A2 => n12188, B1 => n17024, B2 => 
                           n16793, ZN => n9078);
   U3509 : OAI22_X1 port map( A1 => n17041, A2 => n15052, B1 => n17037, B2 => 
                           n16793, ZN => n9079);
   U3510 : OAI22_X1 port map( A1 => n17054, A2 => n14393, B1 => n17050, B2 => 
                           n16793, ZN => n9080);
   U3511 : OAI22_X1 port map( A1 => n17067, A2 => n15168, B1 => n17063, B2 => 
                           n16793, ZN => n9081);
   U3512 : OAI22_X1 port map( A1 => n17080, A2 => n15611, B1 => n17076, B2 => 
                           n16794, ZN => n9082);
   U3513 : OAI22_X1 port map( A1 => n17093, A2 => n15511, B1 => n17089, B2 => 
                           n16794, ZN => n9083);
   U3514 : OAI22_X1 port map( A1 => n17106, A2 => n11860, B1 => n17102, B2 => 
                           n16794, ZN => n9084);
   U3515 : OAI22_X1 port map( A1 => n17132, A2 => n15751, B1 => n17128, B2 => 
                           n16794, ZN => n9086);
   U3516 : OAI22_X1 port map( A1 => n17234, A2 => n15388, B1 => n17230, B2 => 
                           n16795, ZN => n9095);
   U3517 : OAI22_X1 port map( A1 => n17247, A2 => n12258, B1 => n17243, B2 => 
                           n16795, ZN => n9096);
   U3518 : OAI22_X1 port map( A1 => n17260, A2 => n14847, B1 => n17256, B2 => 
                           n16795, ZN => n9097);
   U3519 : OAI22_X1 port map( A1 => n17286, A2 => n14394, B1 => n17282, B2 => 
                           n16795, ZN => n9099);
   U3520 : OAI22_X1 port map( A1 => n17299, A2 => n14621, B1 => n17295, B2 => 
                           n16795, ZN => n9100);
   U3521 : OAI22_X1 port map( A1 => n17325, A2 => n15308, B1 => n17321, B2 => 
                           n16795, ZN => n9102);
   U3522 : OAI22_X1 port map( A1 => n17338, A2 => n11897, B1 => n17334, B2 => 
                           n16795, ZN => n9103);
   U3523 : OAI22_X1 port map( A1 => n17351, A2 => n15103, B1 => n17347, B2 => 
                           n16795, ZN => n9104);
   U3524 : OAI22_X1 port map( A1 => n17364, A2 => n15685, B1 => n17360, B2 => 
                           n16795, ZN => n9105);
   U3525 : OAI22_X1 port map( A1 => n17377, A2 => n14457, B1 => n17373, B2 => 
                           n16796, ZN => n9106);
   U3526 : OAI22_X1 port map( A1 => n17390, A2 => n14745, B1 => n17386, B2 => 
                           n16796, ZN => n9107);
   U3527 : OAI22_X1 port map( A1 => n17403, A2 => n14345, B1 => n17399, B2 => 
                           n16796, ZN => n9108);
   U3528 : OAI22_X1 port map( A1 => n17429, A2 => n15343, B1 => n17425, B2 => 
                           n16796, ZN => n9110);
   U3529 : OAI22_X1 port map( A1 => n17442, A2 => n14038, B1 => n17438, B2 => 
                           n16796, ZN => n9111);
   U3530 : OAI22_X1 port map( A1 => n17455, A2 => n14744, B1 => n17450, B2 => 
                           n16796, ZN => n9112);
   U3531 : OAI22_X1 port map( A1 => n17468, A2 => n15538, B1 => n17464, B2 => 
                           n16796, ZN => n9113);
   U3532 : OAI22_X1 port map( A1 => n17481, A2 => n15775, B1 => n17477, B2 => 
                           n16796, ZN => n9114);
   U3533 : OAI22_X1 port map( A1 => n17494, A2 => n14803, B1 => n17490, B2 => 
                           n16796, ZN => n9115);
   U3534 : OAI22_X1 port map( A1 => n17507, A2 => n15612, B1 => n17503, B2 => 
                           n16796, ZN => n9116);
   U3535 : OAI22_X1 port map( A1 => n17581, A2 => n14264, B1 => n17576, B2 => 
                           n16797, ZN => n9121);
   U3536 : OAI22_X1 port map( A1 => n18008, A2 => n12105, B1 => n18004, B2 => 
                           n16798, ZN => n9134);
   U3537 : OAI22_X1 port map( A1 => n18021, A2 => n14586, B1 => n18017, B2 => 
                           n16798, ZN => n9135);
   U3538 : OAI22_X1 port map( A1 => n16939, A2 => n14563, B1 => n16935, B2 => 
                           n16799, ZN => n9142);
   U3539 : OAI22_X1 port map( A1 => n17028, A2 => n12189, B1 => n17024, B2 => 
                           n16799, ZN => n9150);
   U3540 : OAI22_X1 port map( A1 => n17041, A2 => n15053, B1 => n17037, B2 => 
                           n16799, ZN => n9151);
   U3541 : OAI22_X1 port map( A1 => n17054, A2 => n14395, B1 => n17050, B2 => 
                           n16799, ZN => n9152);
   U3542 : OAI22_X1 port map( A1 => n17080, A2 => n15613, B1 => n17076, B2 => 
                           n16800, ZN => n9154);
   U3543 : OAI22_X1 port map( A1 => n17132, A2 => n15752, B1 => n17128, B2 => 
                           n16800, ZN => n9158);
   U3544 : OAI22_X1 port map( A1 => n17234, A2 => n15389, B1 => n17230, B2 => 
                           n16801, ZN => n9167);
   U3545 : OAI22_X1 port map( A1 => n17247, A2 => n12301, B1 => n17243, B2 => 
                           n16801, ZN => n9168);
   U3546 : OAI22_X1 port map( A1 => n17325, A2 => n15309, B1 => n17321, B2 => 
                           n16801, ZN => n9174);
   U3547 : OAI22_X1 port map( A1 => n17338, A2 => n11898, B1 => n17334, B2 => 
                           n16801, ZN => n9175);
   U3548 : OAI22_X1 port map( A1 => n17351, A2 => n15105, B1 => n17347, B2 => 
                           n16801, ZN => n9176);
   U3549 : OAI22_X1 port map( A1 => n17377, A2 => n14459, B1 => n17373, B2 => 
                           n16802, ZN => n9178);
   U3550 : OAI22_X1 port map( A1 => n17428, A2 => n15344, B1 => n17425, B2 => 
                           n16802, ZN => n9182);
   U3551 : OAI22_X1 port map( A1 => n17441, A2 => n14040, B1 => n17438, B2 => 
                           n16802, ZN => n9183);
   U3552 : OAI22_X1 port map( A1 => n17454, A2 => n14746, B1 => n17450, B2 => 
                           n16802, ZN => n9184);
   U3553 : OAI22_X1 port map( A1 => n17480, A2 => n15776, B1 => n17477, B2 => 
                           n16802, ZN => n9186);
   U3554 : OAI22_X1 port map( A1 => n18008, A2 => n12148, B1 => n18004, B2 => 
                           n16804, ZN => n9206);
   U3555 : OAI22_X1 port map( A1 => n16939, A2 => n14564, B1 => n16935, B2 => 
                           n16805, ZN => n9214);
   U3556 : OAI22_X1 port map( A1 => n17027, A2 => n12190, B1 => n17024, B2 => 
                           n16805, ZN => n9222);
   U3557 : OAI22_X1 port map( A1 => n17132, A2 => n15753, B1 => n17128, B2 => 
                           n16806, ZN => n9230);
   U3558 : OAI22_X1 port map( A1 => n17324, A2 => n15310, B1 => n17321, B2 => 
                           n16807, ZN => n9246);
   U3559 : OAI22_X1 port map( A1 => n17428, A2 => n15345, B1 => n17425, B2 => 
                           n16808, ZN => n9254);
   U3560 : OAI22_X1 port map( A1 => n17582, A2 => n14268, B1 => n17576, B2 => 
                           n16821, ZN => n9409);
   U3561 : OAI22_X1 port map( A1 => n18009, A2 => n12152, B1 => n18004, B2 => 
                           n16822, ZN => n9422);
   U3562 : OAI22_X1 port map( A1 => n18022, A2 => n14590, B1 => n18017, B2 => 
                           n16822, ZN => n9423);
   U3563 : OAI22_X1 port map( A1 => n16940, A2 => n14545, B1 => n16935, B2 => 
                           n17514, ZN => n9934);
   U3564 : OAI22_X1 port map( A1 => n17029, A2 => n12170, B1 => n17024, B2 => 
                           n17514, ZN => n9942);
   U3565 : OAI22_X1 port map( A1 => n17042, A2 => n15054, B1 => n17037, B2 => 
                           n17514, ZN => n9943);
   U3566 : OAI22_X1 port map( A1 => n17055, A2 => n14396, B1 => n17050, B2 => 
                           n17514, ZN => n9944);
   U3567 : OAI22_X1 port map( A1 => n17068, A2 => n15169, B1 => n17063, B2 => 
                           n17514, ZN => n9945);
   U3568 : OAI22_X1 port map( A1 => n17081, A2 => n15614, B1 => n17076, B2 => 
                           n17515, ZN => n9946);
   U3569 : OAI22_X1 port map( A1 => n17094, A2 => n15494, B1 => n17089, B2 => 
                           n17515, ZN => n9947);
   U3570 : OAI22_X1 port map( A1 => n17107, A2 => n11861, B1 => n17102, B2 => 
                           n17515, ZN => n9948);
   U3571 : OAI22_X1 port map( A1 => n17133, A2 => n15734, B1 => n17128, B2 => 
                           n17515, ZN => n9950);
   U3572 : OAI22_X1 port map( A1 => n17235, A2 => n15390, B1 => n17230, B2 => 
                           n17516, ZN => n9959);
   U3573 : OAI22_X1 port map( A1 => n17248, A2 => n12204, B1 => n17243, B2 => 
                           n17516, ZN => n9960);
   U3574 : OAI22_X1 port map( A1 => n17261, A2 => n14830, B1 => n17256, B2 => 
                           n17516, ZN => n9961);
   U3575 : OAI22_X1 port map( A1 => n17287, A2 => n14397, B1 => n17282, B2 => 
                           n17516, ZN => n9963);
   U3576 : OAI22_X1 port map( A1 => n17300, A2 => n14604, B1 => n17295, B2 => 
                           n17516, ZN => n9964);
   U3577 : OAI22_X1 port map( A1 => n17326, A2 => n15291, B1 => n17321, B2 => 
                           n17516, ZN => n9966);
   U3578 : OAI22_X1 port map( A1 => n17339, A2 => n11880, B1 => n17334, B2 => 
                           n17516, ZN => n9967);
   U3579 : OAI22_X1 port map( A1 => n17352, A2 => n15070, B1 => n17347, B2 => 
                           n17516, ZN => n9968);
   U3580 : OAI22_X1 port map( A1 => n17365, A2 => n15668, B1 => n17360, B2 => 
                           n17516, ZN => n9969);
   U3581 : OAI22_X1 port map( A1 => n17378, A2 => n14424, B1 => n17373, B2 => 
                           n17517, ZN => n9970);
   U3582 : OAI22_X1 port map( A1 => n17391, A2 => n14710, B1 => n17386, B2 => 
                           n17517, ZN => n9971);
   U3583 : OAI22_X1 port map( A1 => n17404, A2 => n14357, B1 => n17399, B2 => 
                           n17517, ZN => n9972);
   U3584 : OAI22_X1 port map( A1 => n17430, A2 => n15325, B1 => n17425, B2 => 
                           n17517, ZN => n9974);
   U3585 : OAI22_X1 port map( A1 => n17443, A2 => n12347, B1 => n17438, B2 => 
                           n17517, ZN => n9975);
   U3586 : OAI22_X1 port map( A1 => n17456, A2 => n14709, B1 => n17450, B2 => 
                           n17517, ZN => n9976);
   U3587 : OAI22_X1 port map( A1 => n17469, A2 => n15457, B1 => n17464, B2 => 
                           n17517, ZN => n9977);
   U3588 : OAI22_X1 port map( A1 => n17482, A2 => n15735, B1 => n17477, B2 => 
                           n17517, ZN => n9978);
   U3589 : OAI22_X1 port map( A1 => n17495, A2 => n14769, B1 => n17490, B2 => 
                           n17517, ZN => n9979);
   U3590 : OAI22_X1 port map( A1 => n17508, A2 => n15615, B1 => n17503, B2 => 
                           n17517, ZN => n9980);
   U3591 : BUF_X1 port map( A => n4223, Z => n17666);
   U3592 : BUF_X1 port map( A => n4202, Z => n17690);
   U3593 : NAND2_X1 port map( A1 => N273, A2 => n14262, ZN => n14064);
   U3594 : OAI22_X1 port map( A1 => n16700, A2 => n14980, B1 => n16692, B2 => 
                           n16456, ZN => n7981);
   U3595 : OAI22_X1 port map( A1 => n16695, A2 => n14981, B1 => n16691, B2 => 
                           n16815, ZN => n8089);
   U3596 : OAI22_X1 port map( A1 => n16695, A2 => n14982, B1 => n16692, B2 => 
                           n16821, ZN => n8091);
   U3597 : OAI22_X1 port map( A1 => n16694, A2 => n14983, B1 => n16692, B2 => 
                           n16833, ZN => n8095);
   U3598 : OAI22_X1 port map( A1 => n16694, A2 => n14984, B1 => n16691, B2 => 
                           n16839, ZN => n8097);
   U3599 : OAI22_X1 port map( A1 => n16694, A2 => n14985, B1 => n16692, B2 => 
                           n16845, ZN => n8099);
   U3600 : OAI22_X1 port map( A1 => n16693, A2 => n14986, B1 => n16692, B2 => 
                           n16851, ZN => n8101);
   U3601 : OAI22_X1 port map( A1 => n16695, A2 => n14987, B1 => n16691, B2 => 
                           n16857, ZN => n8103);
   U3602 : OAI22_X1 port map( A1 => n16694, A2 => n14988, B1 => n16692, B2 => 
                           n17512, ZN => n8105);
   U3603 : OAI22_X1 port map( A1 => n18008, A2 => n12150, B1 => n18003, B2 => 
                           n16810, ZN => n9278);
   U3604 : OAI22_X1 port map( A1 => n16938, A2 => n14565, B1 => n16934, B2 => 
                           n16811, ZN => n9286);
   U3605 : OAI22_X1 port map( A1 => n17027, A2 => n12191, B1 => n17023, B2 => 
                           n16811, ZN => n9294);
   U3606 : OAI22_X1 port map( A1 => n17131, A2 => n15754, B1 => n17127, B2 => 
                           n16812, ZN => n9302);
   U3607 : OAI22_X1 port map( A1 => n17324, A2 => n15311, B1 => n17320, B2 => 
                           n16813, ZN => n9318);
   U3608 : OAI22_X1 port map( A1 => n17428, A2 => n15346, B1 => n17424, B2 => 
                           n16814, ZN => n9326);
   U3609 : OAI22_X1 port map( A1 => n18007, A2 => n12151, B1 => n18003, B2 => 
                           n16816, ZN => n9350);
   U3610 : OAI22_X1 port map( A1 => n16938, A2 => n14566, B1 => n16934, B2 => 
                           n16817, ZN => n9358);
   U3611 : OAI22_X1 port map( A1 => n17027, A2 => n12192, B1 => n17023, B2 => 
                           n16817, ZN => n9366);
   U3612 : OAI22_X1 port map( A1 => n17131, A2 => n15755, B1 => n17127, B2 => 
                           n16818, ZN => n9374);
   U3613 : OAI22_X1 port map( A1 => n17324, A2 => n15312, B1 => n17320, B2 => 
                           n16819, ZN => n9390);
   U3614 : OAI22_X1 port map( A1 => n17428, A2 => n15347, B1 => n17424, B2 => 
                           n16820, ZN => n9398);
   U3615 : OAI22_X1 port map( A1 => n16938, A2 => n14567, B1 => n16934, B2 => 
                           n16823, ZN => n9430);
   U3616 : OAI22_X1 port map( A1 => n17027, A2 => n12193, B1 => n17023, B2 => 
                           n16823, ZN => n9438);
   U3617 : OAI22_X1 port map( A1 => n17131, A2 => n15756, B1 => n17127, B2 => 
                           n16824, ZN => n9446);
   U3618 : OAI22_X1 port map( A1 => n17323, A2 => n15313, B1 => n17320, B2 => 
                           n16825, ZN => n9462);
   U3619 : OAI22_X1 port map( A1 => n17427, A2 => n15348, B1 => n17424, B2 => 
                           n16826, ZN => n9470);
   U3620 : OAI22_X1 port map( A1 => n18007, A2 => n12153, B1 => n18003, B2 => 
                           n16828, ZN => n9494);
   U3621 : OAI22_X1 port map( A1 => n16937, A2 => n14568, B1 => n16934, B2 => 
                           n16829, ZN => n9502);
   U3622 : OAI22_X1 port map( A1 => n17026, A2 => n12164, B1 => n17023, B2 => 
                           n16829, ZN => n9510);
   U3623 : OAI22_X1 port map( A1 => n17130, A2 => n15722, B1 => n17127, B2 => 
                           n16830, ZN => n9518);
   U3624 : OAI22_X1 port map( A1 => n17323, A2 => n15285, B1 => n17320, B2 => 
                           n16831, ZN => n9534);
   U3625 : OAI22_X1 port map( A1 => n17427, A2 => n15319, B1 => n17424, B2 => 
                           n16832, ZN => n9542);
   U3626 : OAI22_X1 port map( A1 => n18007, A2 => n12154, B1 => n18003, B2 => 
                           n16834, ZN => n9566);
   U3627 : OAI22_X1 port map( A1 => n16938, A2 => n14540, B1 => n16934, B2 => 
                           n16835, ZN => n9574);
   U3628 : OAI22_X1 port map( A1 => n17026, A2 => n12165, B1 => n17023, B2 => 
                           n16835, ZN => n9582);
   U3629 : OAI22_X1 port map( A1 => n17131, A2 => n15724, B1 => n17127, B2 => 
                           n16836, ZN => n9590);
   U3630 : OAI22_X1 port map( A1 => n17324, A2 => n15286, B1 => n17320, B2 => 
                           n16837, ZN => n9606);
   U3631 : OAI22_X1 port map( A1 => n17427, A2 => n15320, B1 => n17424, B2 => 
                           n16838, ZN => n9614);
   U3632 : OAI22_X1 port map( A1 => n18007, A2 => n12155, B1 => n18003, B2 => 
                           n16840, ZN => n9638);
   U3633 : OAI22_X1 port map( A1 => n16937, A2 => n14541, B1 => n16934, B2 => 
                           n16841, ZN => n9646);
   U3634 : OAI22_X1 port map( A1 => n17026, A2 => n12166, B1 => n17023, B2 => 
                           n16841, ZN => n9654);
   U3635 : OAI22_X1 port map( A1 => n17130, A2 => n15726, B1 => n17127, B2 => 
                           n16842, ZN => n9662);
   U3636 : OAI22_X1 port map( A1 => n17323, A2 => n15287, B1 => n17320, B2 => 
                           n16843, ZN => n9678);
   U3637 : OAI22_X1 port map( A1 => n17427, A2 => n15321, B1 => n17424, B2 => 
                           n16844, ZN => n9686);
   U3638 : OAI22_X1 port map( A1 => n18006, A2 => n12156, B1 => n18003, B2 => 
                           n16846, ZN => n9710);
   U3639 : OAI22_X1 port map( A1 => n16937, A2 => n14542, B1 => n16934, B2 => 
                           n16847, ZN => n9718);
   U3640 : OAI22_X1 port map( A1 => n17026, A2 => n12167, B1 => n17023, B2 => 
                           n16847, ZN => n9726);
   U3641 : OAI22_X1 port map( A1 => n17130, A2 => n15728, B1 => n17127, B2 => 
                           n16848, ZN => n9734);
   U3642 : OAI22_X1 port map( A1 => n17323, A2 => n15288, B1 => n17320, B2 => 
                           n16849, ZN => n9750);
   U3643 : OAI22_X1 port map( A1 => n17426, A2 => n15322, B1 => n17424, B2 => 
                           n16850, ZN => n9758);
   U3644 : OAI22_X1 port map( A1 => n18006, A2 => n12157, B1 => n18003, B2 => 
                           n16852, ZN => n9782);
   U3645 : OAI22_X1 port map( A1 => n16937, A2 => n14543, B1 => n16934, B2 => 
                           n16853, ZN => n9790);
   U3646 : OAI22_X1 port map( A1 => n17025, A2 => n12168, B1 => n17023, B2 => 
                           n16853, ZN => n9798);
   U3647 : OAI22_X1 port map( A1 => n17130, A2 => n15730, B1 => n17127, B2 => 
                           n16854, ZN => n9806);
   U3648 : OAI22_X1 port map( A1 => n17322, A2 => n15289, B1 => n17320, B2 => 
                           n16855, ZN => n9822);
   U3649 : OAI22_X1 port map( A1 => n17426, A2 => n15323, B1 => n17424, B2 => 
                           n16856, ZN => n9830);
   U3650 : OAI22_X1 port map( A1 => n18006, A2 => n12158, B1 => n18003, B2 => 
                           n16858, ZN => n9854);
   U3651 : OAI22_X1 port map( A1 => n16936, A2 => n14544, B1 => n16934, B2 => 
                           n16859, ZN => n9862);
   U3652 : OAI22_X1 port map( A1 => n17025, A2 => n12169, B1 => n17023, B2 => 
                           n16859, ZN => n9870);
   U3653 : OAI22_X1 port map( A1 => n17129, A2 => n15732, B1 => n17127, B2 => 
                           n16860, ZN => n9878);
   U3654 : OAI22_X1 port map( A1 => n17322, A2 => n15290, B1 => n17320, B2 => 
                           n16861, ZN => n9894);
   U3655 : OAI22_X1 port map( A1 => n17426, A2 => n15324, B1 => n17424, B2 => 
                           n16862, ZN => n9902);
   U3656 : OAI22_X1 port map( A1 => n18006, A2 => n12159, B1 => n18003, B2 => 
                           n17513, ZN => n9926_port);
   U3657 : OAI22_X1 port map( A1 => n17581, A2 => n14269, B1 => n17576, B2 => 
                           n16803, ZN => n9193);
   U3658 : OAI22_X1 port map( A1 => n18021, A2 => n14587, B1 => n18016, B2 => 
                           n16804, ZN => n9207);
   U3659 : OAI22_X1 port map( A1 => n17040, A2 => n15055, B1 => n17036, B2 => 
                           n16805, ZN => n9223);
   U3660 : OAI22_X1 port map( A1 => n17053, A2 => n14398, B1 => n17049, B2 => 
                           n16805, ZN => n9224);
   U3661 : OAI22_X1 port map( A1 => n17079, A2 => n15616, B1 => n17075, B2 => 
                           n16806, ZN => n9226);
   U3662 : OAI22_X1 port map( A1 => n17233, A2 => n15391, B1 => n17229, B2 => 
                           n16807, ZN => n9239);
   U3663 : OAI22_X1 port map( A1 => n17246, A2 => n12303, B1 => n17242, B2 => 
                           n16807, ZN => n9240);
   U3664 : OAI22_X1 port map( A1 => n17337, A2 => n11899, B1 => n17333, B2 => 
                           n16807, ZN => n9247);
   U3665 : OAI22_X1 port map( A1 => n17350, A2 => n15107, B1 => n17346, B2 => 
                           n16807, ZN => n9248);
   U3666 : OAI22_X1 port map( A1 => n17376, A2 => n14461, B1 => n17372, B2 => 
                           n16808, ZN => n9250);
   U3667 : OAI22_X1 port map( A1 => n17441, A2 => n14042, B1 => n17437, B2 => 
                           n16808, ZN => n9255);
   U3668 : OAI22_X1 port map( A1 => n17454, A2 => n14748, B1 => n17450, B2 => 
                           n16808, ZN => n9256);
   U3669 : OAI22_X1 port map( A1 => n17480, A2 => n15777, B1 => n17476, B2 => 
                           n16808, ZN => n9258);
   U3670 : OAI22_X1 port map( A1 => n17580, A2 => n14270, B1 => n17576, B2 => 
                           n16809, ZN => n9265);
   U3671 : OAI22_X1 port map( A1 => n18021, A2 => n14588, B1 => n18016, B2 => 
                           n16810, ZN => n9279);
   U3672 : OAI22_X1 port map( A1 => n17040, A2 => n15056, B1 => n17036, B2 => 
                           n16811, ZN => n9295);
   U3673 : OAI22_X1 port map( A1 => n17053, A2 => n14399, B1 => n17049, B2 => 
                           n16811, ZN => n9296);
   U3674 : OAI22_X1 port map( A1 => n17079, A2 => n15617, B1 => n17075, B2 => 
                           n16812, ZN => n9298);
   U3675 : OAI22_X1 port map( A1 => n17233, A2 => n15392, B1 => n17229, B2 => 
                           n16813, ZN => n9311);
   U3676 : OAI22_X1 port map( A1 => n17246, A2 => n12304, B1 => n17242, B2 => 
                           n16813, ZN => n9312);
   U3677 : OAI22_X1 port map( A1 => n17337, A2 => n11900, B1 => n17333, B2 => 
                           n16813, ZN => n9319);
   U3678 : OAI22_X1 port map( A1 => n17350, A2 => n15109, B1 => n17346, B2 => 
                           n16813, ZN => n9320);
   U3679 : OAI22_X1 port map( A1 => n17376, A2 => n14463, B1 => n17372, B2 => 
                           n16814, ZN => n9322);
   U3680 : OAI22_X1 port map( A1 => n17441, A2 => n14044, B1 => n17437, B2 => 
                           n16814, ZN => n9327);
   U3681 : OAI22_X1 port map( A1 => n17454, A2 => n14750, B1 => n17450, B2 => 
                           n16814, ZN => n9328);
   U3682 : OAI22_X1 port map( A1 => n17480, A2 => n15778, B1 => n17476, B2 => 
                           n16814, ZN => n9330);
   U3683 : OAI22_X1 port map( A1 => n17580, A2 => n14271, B1 => n17577, B2 => 
                           n16815, ZN => n9337);
   U3684 : OAI22_X1 port map( A1 => n18020, A2 => n14589, B1 => n18016, B2 => 
                           n16816, ZN => n9351);
   U3685 : OAI22_X1 port map( A1 => n17040, A2 => n15057, B1 => n17036, B2 => 
                           n16817, ZN => n9367);
   U3686 : OAI22_X1 port map( A1 => n17053, A2 => n14400, B1 => n17049, B2 => 
                           n16817, ZN => n9368);
   U3687 : OAI22_X1 port map( A1 => n17079, A2 => n15618, B1 => n17075, B2 => 
                           n16818, ZN => n9370);
   U3688 : OAI22_X1 port map( A1 => n17233, A2 => n15393, B1 => n17229, B2 => 
                           n16819, ZN => n9383);
   U3689 : OAI22_X1 port map( A1 => n17246, A2 => n12305, B1 => n17242, B2 => 
                           n16819, ZN => n9384);
   U3690 : OAI22_X1 port map( A1 => n17337, A2 => n11901, B1 => n17333, B2 => 
                           n16819, ZN => n9391);
   U3691 : OAI22_X1 port map( A1 => n17350, A2 => n15111, B1 => n17346, B2 => 
                           n16819, ZN => n9392);
   U3692 : OAI22_X1 port map( A1 => n17376, A2 => n14465, B1 => n17372, B2 => 
                           n16820, ZN => n9394);
   U3693 : OAI22_X1 port map( A1 => n17441, A2 => n14046, B1 => n17437, B2 => 
                           n16820, ZN => n9399);
   U3694 : OAI22_X1 port map( A1 => n17454, A2 => n14752, B1 => n17451, B2 => 
                           n16820, ZN => n9400);
   U3695 : OAI22_X1 port map( A1 => n17480, A2 => n15779, B1 => n17476, B2 => 
                           n16820, ZN => n9402);
   U3696 : OAI22_X1 port map( A1 => n17040, A2 => n15058, B1 => n17036, B2 => 
                           n16823, ZN => n9439);
   U3697 : OAI22_X1 port map( A1 => n17053, A2 => n14401, B1 => n17049, B2 => 
                           n16823, ZN => n9440);
   U3698 : OAI22_X1 port map( A1 => n17079, A2 => n15619, B1 => n17075, B2 => 
                           n16824, ZN => n9442);
   U3699 : OAI22_X1 port map( A1 => n17233, A2 => n15394, B1 => n17229, B2 => 
                           n16825, ZN => n9455);
   U3700 : OAI22_X1 port map( A1 => n17246, A2 => n12306, B1 => n17242, B2 => 
                           n16825, ZN => n9456);
   U3701 : OAI22_X1 port map( A1 => n17336, A2 => n11902, B1 => n17333, B2 => 
                           n16825, ZN => n9463);
   U3702 : OAI22_X1 port map( A1 => n17349, A2 => n15113, B1 => n17346, B2 => 
                           n16825, ZN => n9464);
   U3703 : OAI22_X1 port map( A1 => n17375, A2 => n14467, B1 => n17372, B2 => 
                           n16826, ZN => n9466);
   U3704 : OAI22_X1 port map( A1 => n17440, A2 => n14048, B1 => n17437, B2 => 
                           n16826, ZN => n9471);
   U3705 : OAI22_X1 port map( A1 => n17453, A2 => n14754, B1 => n17451, B2 => 
                           n16826, ZN => n9472);
   U3706 : OAI22_X1 port map( A1 => n17479, A2 => n15780, B1 => n17476, B2 => 
                           n16826, ZN => n9474);
   U3707 : OAI22_X1 port map( A1 => n17580, A2 => n14272, B1 => n17577, B2 => 
                           n16827, ZN => n9481);
   U3708 : OAI22_X1 port map( A1 => n18020, A2 => n14591, B1 => n18016, B2 => 
                           n16828, ZN => n9495);
   U3709 : OAI22_X1 port map( A1 => n17039, A2 => n15059, B1 => n17036, B2 => 
                           n16829, ZN => n9511);
   U3710 : OAI22_X1 port map( A1 => n17052, A2 => n14402, B1 => n17049, B2 => 
                           n16829, ZN => n9512);
   U3711 : OAI22_X1 port map( A1 => n17078, A2 => n15620, B1 => n17075, B2 => 
                           n16830, ZN => n9514);
   U3712 : OAI22_X1 port map( A1 => n17232, A2 => n15395, B1 => n17229, B2 => 
                           n16831, ZN => n9527);
   U3713 : OAI22_X1 port map( A1 => n17245, A2 => n12198, B1 => n17242, B2 => 
                           n16831, ZN => n9528);
   U3714 : OAI22_X1 port map( A1 => n17336, A2 => n11874, B1 => n17333, B2 => 
                           n16831, ZN => n9535);
   U3715 : OAI22_X1 port map( A1 => n17349, A2 => n15115, B1 => n17346, B2 => 
                           n16831, ZN => n9536);
   U3716 : OAI22_X1 port map( A1 => n17375, A2 => n14469, B1 => n17372, B2 => 
                           n16832, ZN => n9538);
   U3717 : OAI22_X1 port map( A1 => n17440, A2 => n14050, B1 => n17437, B2 => 
                           n16832, ZN => n9543);
   U3718 : OAI22_X1 port map( A1 => n17453, A2 => n14817, B1 => n17451, B2 => 
                           n16832, ZN => n9544);
   U3719 : OAI22_X1 port map( A1 => n17479, A2 => n15723, B1 => n17476, B2 => 
                           n16832, ZN => n9546);
   U3720 : OAI22_X1 port map( A1 => n17579, A2 => n14273, B1 => n17577, B2 => 
                           n16833, ZN => n9553);
   U3721 : OAI22_X1 port map( A1 => n18020, A2 => n14592, B1 => n18016, B2 => 
                           n16834, ZN => n9567);
   U3722 : OAI22_X1 port map( A1 => n17039, A2 => n15060, B1 => n17036, B2 => 
                           n16835, ZN => n9583);
   U3723 : OAI22_X1 port map( A1 => n17052, A2 => n14403, B1 => n17049, B2 => 
                           n16835, ZN => n9584);
   U3724 : OAI22_X1 port map( A1 => n17078, A2 => n15621, B1 => n17075, B2 => 
                           n16836, ZN => n9586);
   U3725 : OAI22_X1 port map( A1 => n17232, A2 => n15396, B1 => n17229, B2 => 
                           n16837, ZN => n9599);
   U3726 : OAI22_X1 port map( A1 => n17245, A2 => n12199, B1 => n17242, B2 => 
                           n16837, ZN => n9600);
   U3727 : OAI22_X1 port map( A1 => n17337, A2 => n11875, B1 => n17333, B2 => 
                           n16837, ZN => n9607);
   U3728 : OAI22_X1 port map( A1 => n17350, A2 => n15065, B1 => n17346, B2 => 
                           n16837, ZN => n9608);
   U3729 : OAI22_X1 port map( A1 => n17376, A2 => n14419, B1 => n17372, B2 => 
                           n16838, ZN => n9610);
   U3730 : OAI22_X1 port map( A1 => n17440, A2 => n12342, B1 => n17437, B2 => 
                           n16838, ZN => n9615);
   U3731 : OAI22_X1 port map( A1 => n17453, A2 => n14818, B1 => n17451, B2 => 
                           n16838, ZN => n9616);
   U3732 : OAI22_X1 port map( A1 => n17479, A2 => n15725, B1 => n17476, B2 => 
                           n16838, ZN => n9618);
   U3733 : OAI22_X1 port map( A1 => n17580, A2 => n14274, B1 => n17577, B2 => 
                           n16839, ZN => n9625);
   U3734 : OAI22_X1 port map( A1 => n18020, A2 => n14593, B1 => n18016, B2 => 
                           n16840, ZN => n9639);
   U3735 : OAI22_X1 port map( A1 => n17039, A2 => n15061, B1 => n17036, B2 => 
                           n16841, ZN => n9655);
   U3736 : OAI22_X1 port map( A1 => n17052, A2 => n14404, B1 => n17049, B2 => 
                           n16841, ZN => n9656);
   U3737 : OAI22_X1 port map( A1 => n17078, A2 => n15622, B1 => n17075, B2 => 
                           n16842, ZN => n9658);
   U3738 : OAI22_X1 port map( A1 => n17232, A2 => n15397, B1 => n17229, B2 => 
                           n16843, ZN => n9671);
   U3739 : OAI22_X1 port map( A1 => n17245, A2 => n12200, B1 => n17242, B2 => 
                           n16843, ZN => n9672);
   U3740 : OAI22_X1 port map( A1 => n17336, A2 => n11876, B1 => n17333, B2 => 
                           n16843, ZN => n9679);
   U3741 : OAI22_X1 port map( A1 => n17349, A2 => n15066, B1 => n17346, B2 => 
                           n16843, ZN => n9680);
   U3742 : OAI22_X1 port map( A1 => n17375, A2 => n14420, B1 => n17372, B2 => 
                           n16844, ZN => n9682);
   U3743 : OAI22_X1 port map( A1 => n17440, A2 => n12343, B1 => n17437, B2 => 
                           n16844, ZN => n9687);
   U3744 : OAI22_X1 port map( A1 => n17453, A2 => n14819, B1 => n17451, B2 => 
                           n16844, ZN => n9688);
   U3745 : OAI22_X1 port map( A1 => n17479, A2 => n15727, B1 => n17476, B2 => 
                           n16844, ZN => n9690);
   U3746 : OAI22_X1 port map( A1 => n17579, A2 => n14275, B1 => n17577, B2 => 
                           n16845, ZN => n9697);
   U3747 : OAI22_X1 port map( A1 => n18019, A2 => n14594, B1 => n18016, B2 => 
                           n16846, ZN => n9711);
   U3748 : OAI22_X1 port map( A1 => n17039, A2 => n15062, B1 => n17036, B2 => 
                           n16847, ZN => n9727);
   U3749 : OAI22_X1 port map( A1 => n17052, A2 => n14405, B1 => n17049, B2 => 
                           n16847, ZN => n9728);
   U3750 : OAI22_X1 port map( A1 => n17078, A2 => n15623, B1 => n17075, B2 => 
                           n16848, ZN => n9730);
   U3751 : OAI22_X1 port map( A1 => n17232, A2 => n15398, B1 => n17229, B2 => 
                           n16849, ZN => n9743);
   U3752 : OAI22_X1 port map( A1 => n17245, A2 => n12201, B1 => n17242, B2 => 
                           n16849, ZN => n9744);
   U3753 : OAI22_X1 port map( A1 => n17336, A2 => n11877, B1 => n17333, B2 => 
                           n16849, ZN => n9751);
   U3754 : OAI22_X1 port map( A1 => n17349, A2 => n15067, B1 => n17346, B2 => 
                           n16849, ZN => n9752);
   U3755 : OAI22_X1 port map( A1 => n17375, A2 => n14421, B1 => n17372, B2 => 
                           n16850, ZN => n9754);
   U3756 : OAI22_X1 port map( A1 => n17439, A2 => n12344, B1 => n17437, B2 => 
                           n16850, ZN => n9759);
   U3757 : OAI22_X1 port map( A1 => n17452, A2 => n14703, B1 => n17451, B2 => 
                           n16850, ZN => n9760);
   U3758 : OAI22_X1 port map( A1 => n17478, A2 => n15729, B1 => n17476, B2 => 
                           n16850, ZN => n9762);
   U3759 : OAI22_X1 port map( A1 => n17579, A2 => n14276, B1 => n17577, B2 => 
                           n16851, ZN => n9769);
   U3760 : OAI22_X1 port map( A1 => n18019, A2 => n14595, B1 => n18016, B2 => 
                           n16852, ZN => n9783);
   U3761 : OAI22_X1 port map( A1 => n17038, A2 => n15063, B1 => n17036, B2 => 
                           n16853, ZN => n9799);
   U3762 : OAI22_X1 port map( A1 => n17051, A2 => n14406, B1 => n17049, B2 => 
                           n16853, ZN => n9800);
   U3763 : OAI22_X1 port map( A1 => n17077, A2 => n15624, B1 => n17075, B2 => 
                           n16854, ZN => n9802);
   U3764 : OAI22_X1 port map( A1 => n17231, A2 => n15399, B1 => n17229, B2 => 
                           n16855, ZN => n9815);
   U3765 : OAI22_X1 port map( A1 => n17244, A2 => n12202, B1 => n17242, B2 => 
                           n16855, ZN => n9816);
   U3766 : OAI22_X1 port map( A1 => n17335, A2 => n11878, B1 => n17333, B2 => 
                           n16855, ZN => n9823);
   U3767 : OAI22_X1 port map( A1 => n17348, A2 => n15068, B1 => n17346, B2 => 
                           n16855, ZN => n9824);
   U3768 : OAI22_X1 port map( A1 => n17374, A2 => n14422, B1 => n17372, B2 => 
                           n16856, ZN => n9826);
   U3769 : OAI22_X1 port map( A1 => n17439, A2 => n12345, B1 => n17437, B2 => 
                           n16856, ZN => n9831);
   U3770 : OAI22_X1 port map( A1 => n17452, A2 => n14705, B1 => n17450, B2 => 
                           n16856, ZN => n9832);
   U3771 : OAI22_X1 port map( A1 => n17478, A2 => n15731, B1 => n17476, B2 => 
                           n16856, ZN => n9834);
   U3772 : OAI22_X1 port map( A1 => n17579, A2 => n14277, B1 => n17576, B2 => 
                           n16857, ZN => n9841);
   U3773 : OAI22_X1 port map( A1 => n18019, A2 => n14596, B1 => n18016, B2 => 
                           n16858, ZN => n9855);
   U3774 : OAI22_X1 port map( A1 => n17038, A2 => n15064, B1 => n17036, B2 => 
                           n16859, ZN => n9871);
   U3775 : OAI22_X1 port map( A1 => n17051, A2 => n14407, B1 => n17049, B2 => 
                           n16859, ZN => n9872);
   U3776 : OAI22_X1 port map( A1 => n17077, A2 => n15625, B1 => n17075, B2 => 
                           n16860, ZN => n9874);
   U3777 : OAI22_X1 port map( A1 => n17231, A2 => n15400, B1 => n17229, B2 => 
                           n16861, ZN => n9887);
   U3778 : OAI22_X1 port map( A1 => n17244, A2 => n12203, B1 => n17242, B2 => 
                           n16861, ZN => n9888);
   U3779 : OAI22_X1 port map( A1 => n17335, A2 => n11879, B1 => n17333, B2 => 
                           n16861, ZN => n9895);
   U3780 : OAI22_X1 port map( A1 => n17348, A2 => n15069, B1 => n17346, B2 => 
                           n16861, ZN => n9896);
   U3781 : OAI22_X1 port map( A1 => n17374, A2 => n14423, B1 => n17372, B2 => 
                           n16862, ZN => n9898);
   U3782 : OAI22_X1 port map( A1 => n17439, A2 => n12346, B1 => n17437, B2 => 
                           n16862, ZN => n9903);
   U3783 : OAI22_X1 port map( A1 => n17452, A2 => n14707, B1 => n17451, B2 => 
                           n16862, ZN => n9904);
   U3784 : OAI22_X1 port map( A1 => n17478, A2 => n15733, B1 => n17476, B2 => 
                           n16862, ZN => n9906);
   U3785 : OAI22_X1 port map( A1 => n17578, A2 => n14278, B1 => n17577, B2 => 
                           n17512, ZN => n9913);
   U3786 : OAI22_X1 port map( A1 => n18019, A2 => n14597, B1 => n18016, B2 => 
                           n17513, ZN => n9927);
   U3787 : OAI22_X1 port map( A1 => n17067, A2 => n15170, B1 => n17062, B2 => 
                           n16799, ZN => n9153);
   U3788 : OAI22_X1 port map( A1 => n17093, A2 => n15512, B1 => n17088, B2 => 
                           n16800, ZN => n9155);
   U3789 : OAI22_X1 port map( A1 => n17106, A2 => n11862, B1 => n17101, B2 => 
                           n16800, ZN => n9156);
   U3790 : OAI22_X1 port map( A1 => n17260, A2 => n14848, B1 => n17255, B2 => 
                           n16801, ZN => n9169);
   U3791 : OAI22_X1 port map( A1 => n17286, A2 => n14408, B1 => n17281, B2 => 
                           n16801, ZN => n9171);
   U3792 : OAI22_X1 port map( A1 => n17299, A2 => n14622, B1 => n17294, B2 => 
                           n16801, ZN => n9172);
   U3793 : OAI22_X1 port map( A1 => n17364, A2 => n15686, B1 => n17359, B2 => 
                           n16801, ZN => n9177);
   U3794 : OAI22_X1 port map( A1 => n17390, A2 => n14747, B1 => n17385, B2 => 
                           n16802, ZN => n9179);
   U3795 : OAI22_X1 port map( A1 => n17403, A2 => n14346, B1 => n17398, B2 => 
                           n16802, ZN => n9180);
   U3796 : OAI22_X1 port map( A1 => n17467, A2 => n15539, B1 => n17463, B2 => 
                           n16802, ZN => n9185);
   U3797 : OAI22_X1 port map( A1 => n17493, A2 => n14805, B1 => n17489, B2 => 
                           n16802, ZN => n9187);
   U3798 : OAI22_X1 port map( A1 => n17506, A2 => n15626, B1 => n17502, B2 => 
                           n16802, ZN => n9188);
   U3799 : OAI22_X1 port map( A1 => n17066, A2 => n15171, B1 => n17062, B2 => 
                           n16805, ZN => n9225);
   U3800 : OAI22_X1 port map( A1 => n17092, A2 => n15513, B1 => n17088, B2 => 
                           n16806, ZN => n9227);
   U3801 : OAI22_X1 port map( A1 => n17105, A2 => n11863, B1 => n17101, B2 => 
                           n16806, ZN => n9228);
   U3802 : OAI22_X1 port map( A1 => n17259, A2 => n14849, B1 => n17255, B2 => 
                           n16807, ZN => n9241);
   U3803 : OAI22_X1 port map( A1 => n17285, A2 => n14409, B1 => n17281, B2 => 
                           n16807, ZN => n9243);
   U3804 : OAI22_X1 port map( A1 => n17298, A2 => n14623, B1 => n17294, B2 => 
                           n16807, ZN => n9244);
   U3805 : OAI22_X1 port map( A1 => n17363, A2 => n15687, B1 => n17359, B2 => 
                           n16807, ZN => n9249);
   U3806 : OAI22_X1 port map( A1 => n17389, A2 => n14749, B1 => n17385, B2 => 
                           n16808, ZN => n9251);
   U3807 : OAI22_X1 port map( A1 => n17402, A2 => n14347, B1 => n17398, B2 => 
                           n16808, ZN => n9252);
   U3808 : OAI22_X1 port map( A1 => n17467, A2 => n15540, B1 => n17463, B2 => 
                           n16808, ZN => n9257);
   U3809 : OAI22_X1 port map( A1 => n17493, A2 => n14807, B1 => n17489, B2 => 
                           n16808, ZN => n9259);
   U3810 : OAI22_X1 port map( A1 => n17506, A2 => n15627, B1 => n17502, B2 => 
                           n16808, ZN => n9260);
   U3811 : OAI22_X1 port map( A1 => n17066, A2 => n15172, B1 => n17062, B2 => 
                           n16811, ZN => n9297);
   U3812 : OAI22_X1 port map( A1 => n17092, A2 => n15514, B1 => n17088, B2 => 
                           n16812, ZN => n9299);
   U3813 : OAI22_X1 port map( A1 => n17105, A2 => n11864, B1 => n17101, B2 => 
                           n16812, ZN => n9300);
   U3814 : OAI22_X1 port map( A1 => n17259, A2 => n14850, B1 => n17255, B2 => 
                           n16813, ZN => n9313);
   U3815 : OAI22_X1 port map( A1 => n17285, A2 => n14410, B1 => n17281, B2 => 
                           n16813, ZN => n9315);
   U3816 : OAI22_X1 port map( A1 => n17298, A2 => n14624, B1 => n17294, B2 => 
                           n16813, ZN => n9316);
   U3817 : OAI22_X1 port map( A1 => n17363, A2 => n15688, B1 => n17359, B2 => 
                           n16813, ZN => n9321);
   U3818 : OAI22_X1 port map( A1 => n17389, A2 => n14751, B1 => n17385, B2 => 
                           n16814, ZN => n9323);
   U3819 : OAI22_X1 port map( A1 => n17402, A2 => n14348, B1 => n17398, B2 => 
                           n16814, ZN => n9324);
   U3820 : OAI22_X1 port map( A1 => n17467, A2 => n15541, B1 => n17463, B2 => 
                           n16814, ZN => n9329);
   U3821 : OAI22_X1 port map( A1 => n17493, A2 => n14809, B1 => n17489, B2 => 
                           n16814, ZN => n9331);
   U3822 : OAI22_X1 port map( A1 => n17506, A2 => n15628, B1 => n17502, B2 => 
                           n16814, ZN => n9332);
   U3823 : OAI22_X1 port map( A1 => n17066, A2 => n15173, B1 => n17062, B2 => 
                           n16817, ZN => n9369);
   U3824 : OAI22_X1 port map( A1 => n17092, A2 => n15515, B1 => n17088, B2 => 
                           n16818, ZN => n9371);
   U3825 : OAI22_X1 port map( A1 => n17105, A2 => n11865, B1 => n17101, B2 => 
                           n16818, ZN => n9372);
   U3826 : OAI22_X1 port map( A1 => n17259, A2 => n14851, B1 => n17255, B2 => 
                           n16819, ZN => n9385);
   U3827 : OAI22_X1 port map( A1 => n17285, A2 => n14411, B1 => n17281, B2 => 
                           n16819, ZN => n9387);
   U3828 : OAI22_X1 port map( A1 => n17298, A2 => n14625, B1 => n17294, B2 => 
                           n16819, ZN => n9388);
   U3829 : OAI22_X1 port map( A1 => n17363, A2 => n15689, B1 => n17359, B2 => 
                           n16819, ZN => n9393);
   U3830 : OAI22_X1 port map( A1 => n17389, A2 => n14753, B1 => n17385, B2 => 
                           n16820, ZN => n9395);
   U3831 : OAI22_X1 port map( A1 => n17402, A2 => n14349, B1 => n17398, B2 => 
                           n16820, ZN => n9396);
   U3832 : OAI22_X1 port map( A1 => n17467, A2 => n15542, B1 => n17463, B2 => 
                           n16820, ZN => n9401);
   U3833 : OAI22_X1 port map( A1 => n17493, A2 => n14811, B1 => n17489, B2 => 
                           n16820, ZN => n9403);
   U3834 : OAI22_X1 port map( A1 => n17506, A2 => n15629, B1 => n17502, B2 => 
                           n16820, ZN => n9404);
   U3835 : OAI22_X1 port map( A1 => n17066, A2 => n15174, B1 => n17062, B2 => 
                           n16823, ZN => n9441);
   U3836 : OAI22_X1 port map( A1 => n17092, A2 => n15516, B1 => n17088, B2 => 
                           n16824, ZN => n9443);
   U3837 : OAI22_X1 port map( A1 => n17105, A2 => n11866, B1 => n17101, B2 => 
                           n16824, ZN => n9444);
   U3838 : OAI22_X1 port map( A1 => n17259, A2 => n14852, B1 => n17255, B2 => 
                           n16825, ZN => n9457);
   U3839 : OAI22_X1 port map( A1 => n17285, A2 => n14412, B1 => n17281, B2 => 
                           n16825, ZN => n9459);
   U3840 : OAI22_X1 port map( A1 => n17298, A2 => n14626, B1 => n17294, B2 => 
                           n16825, ZN => n9460);
   U3841 : OAI22_X1 port map( A1 => n17362, A2 => n15690, B1 => n17359, B2 => 
                           n16825, ZN => n9465);
   U3842 : OAI22_X1 port map( A1 => n17388, A2 => n14755, B1 => n17385, B2 => 
                           n16826, ZN => n9467);
   U3843 : OAI22_X1 port map( A1 => n17401, A2 => n14350, B1 => n17398, B2 => 
                           n16826, ZN => n9468);
   U3844 : OAI22_X1 port map( A1 => n17466, A2 => n15543, B1 => n17463, B2 => 
                           n16826, ZN => n9473);
   U3845 : OAI22_X1 port map( A1 => n17492, A2 => n14813, B1 => n17489, B2 => 
                           n16826, ZN => n9475);
   U3846 : OAI22_X1 port map( A1 => n17505, A2 => n15630, B1 => n17502, B2 => 
                           n16826, ZN => n9476);
   U3847 : OAI22_X1 port map( A1 => n17065, A2 => n15175, B1 => n17062, B2 => 
                           n16829, ZN => n9513);
   U3848 : OAI22_X1 port map( A1 => n17091, A2 => n15488, B1 => n17088, B2 => 
                           n16830, ZN => n9515);
   U3849 : OAI22_X1 port map( A1 => n17104, A2 => n11867, B1 => n17101, B2 => 
                           n16830, ZN => n9516);
   U3850 : OAI22_X1 port map( A1 => n17258, A2 => n14824, B1 => n17255, B2 => 
                           n16831, ZN => n9529);
   U3851 : OAI22_X1 port map( A1 => n17284, A2 => n14413, B1 => n17281, B2 => 
                           n16831, ZN => n9531);
   U3852 : OAI22_X1 port map( A1 => n17297, A2 => n14598, B1 => n17294, B2 => 
                           n16831, ZN => n9532);
   U3853 : OAI22_X1 port map( A1 => n17362, A2 => n15662, B1 => n17359, B2 => 
                           n16831, ZN => n9537);
   U3854 : OAI22_X1 port map( A1 => n17388, A2 => n14700, B1 => n17385, B2 => 
                           n16832, ZN => n9539);
   U3855 : OAI22_X1 port map( A1 => n17401, A2 => n14351, B1 => n17398, B2 => 
                           n16832, ZN => n9540);
   U3856 : OAI22_X1 port map( A1 => n17466, A2 => n15544, B1 => n17463, B2 => 
                           n16832, ZN => n9545);
   U3857 : OAI22_X1 port map( A1 => n17492, A2 => n14757, B1 => n17489, B2 => 
                           n16832, ZN => n9547);
   U3858 : OAI22_X1 port map( A1 => n17505, A2 => n15631, B1 => n17502, B2 => 
                           n16832, ZN => n9548);
   U3859 : OAI22_X1 port map( A1 => n17065, A2 => n15176, B1 => n17062, B2 => 
                           n16835, ZN => n9585);
   U3860 : OAI22_X1 port map( A1 => n17091, A2 => n15489, B1 => n17088, B2 => 
                           n16836, ZN => n9587);
   U3861 : OAI22_X1 port map( A1 => n17104, A2 => n11869, B1 => n17101, B2 => 
                           n16836, ZN => n9588);
   U3862 : OAI22_X1 port map( A1 => n17258, A2 => n14825, B1 => n17255, B2 => 
                           n16837, ZN => n9601);
   U3863 : OAI22_X1 port map( A1 => n17284, A2 => n14414, B1 => n17281, B2 => 
                           n16837, ZN => n9603);
   U3864 : OAI22_X1 port map( A1 => n17297, A2 => n14599, B1 => n17294, B2 => 
                           n16837, ZN => n9604);
   U3865 : OAI22_X1 port map( A1 => n17363, A2 => n15663, B1 => n17359, B2 => 
                           n16837, ZN => n9609);
   U3866 : OAI22_X1 port map( A1 => n17389, A2 => n14701, B1 => n17385, B2 => 
                           n16838, ZN => n9611);
   U3867 : OAI22_X1 port map( A1 => n17402, A2 => n14352, B1 => n17398, B2 => 
                           n16838, ZN => n9612);
   U3868 : OAI22_X1 port map( A1 => n17466, A2 => n15452, B1 => n17463, B2 => 
                           n16838, ZN => n9617);
   U3869 : OAI22_X1 port map( A1 => n17492, A2 => n14759, B1 => n17489, B2 => 
                           n16838, ZN => n9619);
   U3870 : OAI22_X1 port map( A1 => n17505, A2 => n15632, B1 => n17502, B2 => 
                           n16838, ZN => n9620);
   U3871 : OAI22_X1 port map( A1 => n17065, A2 => n15177, B1 => n17062, B2 => 
                           n16841, ZN => n9657);
   U3872 : OAI22_X1 port map( A1 => n17091, A2 => n15490, B1 => n17088, B2 => 
                           n16842, ZN => n9659);
   U3873 : OAI22_X1 port map( A1 => n17104, A2 => n11870, B1 => n17101, B2 => 
                           n16842, ZN => n9660);
   U3874 : OAI22_X1 port map( A1 => n17258, A2 => n14826, B1 => n17255, B2 => 
                           n16843, ZN => n9673);
   U3875 : OAI22_X1 port map( A1 => n17284, A2 => n14415, B1 => n17281, B2 => 
                           n16843, ZN => n9675);
   U3876 : OAI22_X1 port map( A1 => n17297, A2 => n14600, B1 => n17294, B2 => 
                           n16843, ZN => n9676);
   U3877 : OAI22_X1 port map( A1 => n17362, A2 => n15664, B1 => n17359, B2 => 
                           n16843, ZN => n9681);
   U3878 : OAI22_X1 port map( A1 => n17388, A2 => n14702, B1 => n17385, B2 => 
                           n16844, ZN => n9683);
   U3879 : OAI22_X1 port map( A1 => n17401, A2 => n14353, B1 => n17398, B2 => 
                           n16844, ZN => n9684);
   U3880 : OAI22_X1 port map( A1 => n17466, A2 => n15453, B1 => n17463, B2 => 
                           n16844, ZN => n9689);
   U3881 : OAI22_X1 port map( A1 => n17492, A2 => n14761, B1 => n17489, B2 => 
                           n16844, ZN => n9691);
   U3882 : OAI22_X1 port map( A1 => n17505, A2 => n15633, B1 => n17502, B2 => 
                           n16844, ZN => n9692);
   U3883 : OAI22_X1 port map( A1 => n17065, A2 => n15178, B1 => n17062, B2 => 
                           n16847, ZN => n9729);
   U3884 : OAI22_X1 port map( A1 => n17091, A2 => n15491, B1 => n17088, B2 => 
                           n16848, ZN => n9731);
   U3885 : OAI22_X1 port map( A1 => n17104, A2 => n11871, B1 => n17101, B2 => 
                           n16848, ZN => n9732);
   U3886 : OAI22_X1 port map( A1 => n17258, A2 => n14827, B1 => n17255, B2 => 
                           n16849, ZN => n9745);
   U3887 : OAI22_X1 port map( A1 => n17284, A2 => n14416, B1 => n17281, B2 => 
                           n16849, ZN => n9747);
   U3888 : OAI22_X1 port map( A1 => n17297, A2 => n14601, B1 => n17294, B2 => 
                           n16849, ZN => n9748);
   U3889 : OAI22_X1 port map( A1 => n17362, A2 => n15665, B1 => n17359, B2 => 
                           n16849, ZN => n9753);
   U3890 : OAI22_X1 port map( A1 => n17388, A2 => n14704, B1 => n17385, B2 => 
                           n16850, ZN => n9755);
   U3891 : OAI22_X1 port map( A1 => n17401, A2 => n14354, B1 => n17398, B2 => 
                           n16850, ZN => n9756);
   U3892 : OAI22_X1 port map( A1 => n17465, A2 => n15454, B1 => n17463, B2 => 
                           n16850, ZN => n9761);
   U3893 : OAI22_X1 port map( A1 => n17491, A2 => n14763, B1 => n17489, B2 => 
                           n16850, ZN => n9763);
   U3894 : OAI22_X1 port map( A1 => n17504, A2 => n15634, B1 => n17502, B2 => 
                           n16850, ZN => n9764);
   U3895 : OAI22_X1 port map( A1 => n17064, A2 => n15179, B1 => n17062, B2 => 
                           n16853, ZN => n9801);
   U3896 : OAI22_X1 port map( A1 => n17090, A2 => n15492, B1 => n17088, B2 => 
                           n16854, ZN => n9803);
   U3897 : OAI22_X1 port map( A1 => n17103, A2 => n11872, B1 => n17101, B2 => 
                           n16854, ZN => n9804);
   U3898 : OAI22_X1 port map( A1 => n17257, A2 => n14828, B1 => n17255, B2 => 
                           n16855, ZN => n9817);
   U3899 : OAI22_X1 port map( A1 => n17283, A2 => n14417, B1 => n17281, B2 => 
                           n16855, ZN => n9819);
   U3900 : OAI22_X1 port map( A1 => n17296, A2 => n14602, B1 => n17294, B2 => 
                           n16855, ZN => n9820);
   U3901 : OAI22_X1 port map( A1 => n17361, A2 => n15666, B1 => n17359, B2 => 
                           n16855, ZN => n9825);
   U3902 : OAI22_X1 port map( A1 => n17387, A2 => n14706, B1 => n17385, B2 => 
                           n16856, ZN => n9827);
   U3903 : OAI22_X1 port map( A1 => n17400, A2 => n14355, B1 => n17398, B2 => 
                           n16856, ZN => n9828);
   U3904 : OAI22_X1 port map( A1 => n17465, A2 => n15455, B1 => n17463, B2 => 
                           n16856, ZN => n9833);
   U3905 : OAI22_X1 port map( A1 => n17491, A2 => n14765, B1 => n17489, B2 => 
                           n16856, ZN => n9835);
   U3906 : OAI22_X1 port map( A1 => n17504, A2 => n15635, B1 => n17502, B2 => 
                           n16856, ZN => n9836);
   U3907 : OAI22_X1 port map( A1 => n17064, A2 => n15180, B1 => n17062, B2 => 
                           n16859, ZN => n9873);
   U3908 : OAI22_X1 port map( A1 => n17090, A2 => n15493, B1 => n17088, B2 => 
                           n16860, ZN => n9875);
   U3909 : OAI22_X1 port map( A1 => n17103, A2 => n11873, B1 => n17101, B2 => 
                           n16860, ZN => n9876);
   U3910 : OAI22_X1 port map( A1 => n17257, A2 => n14829, B1 => n17255, B2 => 
                           n16861, ZN => n9889);
   U3911 : OAI22_X1 port map( A1 => n17283, A2 => n14418, B1 => n17281, B2 => 
                           n16861, ZN => n9891);
   U3912 : OAI22_X1 port map( A1 => n17296, A2 => n14603, B1 => n17294, B2 => 
                           n16861, ZN => n9892);
   U3913 : OAI22_X1 port map( A1 => n17361, A2 => n15667, B1 => n17359, B2 => 
                           n16861, ZN => n9897);
   U3914 : OAI22_X1 port map( A1 => n17387, A2 => n14708, B1 => n17385, B2 => 
                           n16862, ZN => n9899);
   U3915 : OAI22_X1 port map( A1 => n17400, A2 => n14356, B1 => n17398, B2 => 
                           n16862, ZN => n9900);
   U3916 : OAI22_X1 port map( A1 => n17465, A2 => n15456, B1 => n17463, B2 => 
                           n16862, ZN => n9905);
   U3917 : OAI22_X1 port map( A1 => n17491, A2 => n14767, B1 => n17489, B2 => 
                           n16862, ZN => n9907);
   U3918 : OAI22_X1 port map( A1 => n17504, A2 => n15636, B1 => n17502, B2 => 
                           n16862, ZN => n9908_port);
   U3919 : OAI22_X1 port map( A1 => n17122, A2 => n12315, B1 => n17115, B2 => 
                           n16727, ZN => n8293);
   U3920 : OAI22_X1 port map( A1 => n17315, A2 => n15704, B1 => n17308, B2 => 
                           n16728, ZN => n8309);
   U3921 : OAI22_X1 port map( A1 => n17419, A2 => n15215, B1 => n17412, B2 => 
                           n16729, ZN => n8317);
   U3922 : OAI22_X1 port map( A1 => n17122, A2 => n12316, B1 => n17115, B2 => 
                           n16734, ZN => n8365);
   U3923 : OAI22_X1 port map( A1 => n17315, A2 => n15705, B1 => n17308, B2 => 
                           n16735, ZN => n8381);
   U3924 : OAI22_X1 port map( A1 => n17419, A2 => n15216, B1 => n17412, B2 => 
                           n16736, ZN => n8389);
   U3925 : OAI22_X1 port map( A1 => n17121, A2 => n12317, B1 => n17115, B2 => 
                           n16740, ZN => n8437);
   U3926 : OAI22_X1 port map( A1 => n17314, A2 => n15706, B1 => n17308, B2 => 
                           n16741, ZN => n8453);
   U3927 : OAI22_X1 port map( A1 => n17418, A2 => n15217, B1 => n17412, B2 => 
                           n16742, ZN => n8461);
   U3928 : OAI22_X1 port map( A1 => n17121, A2 => n12318, B1 => n17115, B2 => 
                           n16746, ZN => n8509);
   U3929 : OAI22_X1 port map( A1 => n17314, A2 => n15707, B1 => n17308, B2 => 
                           n16747, ZN => n8525);
   U3930 : OAI22_X1 port map( A1 => n17418, A2 => n15218, B1 => n17412, B2 => 
                           n16748, ZN => n8533);
   U3931 : OAI22_X1 port map( A1 => n17121, A2 => n12319, B1 => n17115, B2 => 
                           n16752, ZN => n8581);
   U3932 : OAI22_X1 port map( A1 => n17314, A2 => n15708, B1 => n17308, B2 => 
                           n16753, ZN => n8597);
   U3933 : OAI22_X1 port map( A1 => n17418, A2 => n15219, B1 => n17412, B2 => 
                           n16754, ZN => n8605);
   U3934 : OAI22_X1 port map( A1 => n17121, A2 => n12320, B1 => n17115, B2 => 
                           n16758, ZN => n8653);
   U3935 : OAI22_X1 port map( A1 => n17314, A2 => n15709, B1 => n17308, B2 => 
                           n16759, ZN => n8669);
   U3936 : OAI22_X1 port map( A1 => n17418, A2 => n15220, B1 => n17412, B2 => 
                           n16760, ZN => n8677);
   U3937 : OAI22_X1 port map( A1 => n17120, A2 => n12321, B1 => n17115, B2 => 
                           n16764, ZN => n8725);
   U3938 : OAI22_X1 port map( A1 => n17313, A2 => n15710, B1 => n17308, B2 => 
                           n16765, ZN => n8741);
   U3939 : OAI22_X1 port map( A1 => n17417, A2 => n15221, B1 => n17412, B2 => 
                           n16766, ZN => n8749);
   U3940 : OAI22_X1 port map( A1 => n17120, A2 => n12322, B1 => n17115, B2 => 
                           n16770, ZN => n8797);
   U3941 : OAI22_X1 port map( A1 => n17313, A2 => n15711, B1 => n17308, B2 => 
                           n16771, ZN => n8813);
   U3942 : OAI22_X1 port map( A1 => n17417, A2 => n15222, B1 => n17412, B2 => 
                           n16772, ZN => n8821);
   U3943 : OAI22_X1 port map( A1 => n17120, A2 => n12323, B1 => n17115, B2 => 
                           n16776, ZN => n8869);
   U3944 : OAI22_X1 port map( A1 => n17313, A2 => n15712, B1 => n17308, B2 => 
                           n16777, ZN => n8885);
   U3945 : OAI22_X1 port map( A1 => n17417, A2 => n15223, B1 => n17412, B2 => 
                           n16778, ZN => n8893);
   U3946 : OAI22_X1 port map( A1 => n17119, A2 => n12324, B1 => n17115, B2 => 
                           n16782, ZN => n8941);
   U3947 : OAI22_X1 port map( A1 => n17312, A2 => n15713, B1 => n17308, B2 => 
                           n16783, ZN => n8957);
   U3948 : OAI22_X1 port map( A1 => n17416, A2 => n15224, B1 => n17412, B2 => 
                           n16784, ZN => n8965);
   U3949 : OAI22_X1 port map( A1 => n17119, A2 => n12325, B1 => n17115, B2 => 
                           n16788, ZN => n9013);
   U3950 : OAI22_X1 port map( A1 => n17312, A2 => n15714, B1 => n17308, B2 => 
                           n16789, ZN => n9029);
   U3951 : OAI22_X1 port map( A1 => n17416, A2 => n15225, B1 => n17412, B2 => 
                           n16790, ZN => n9037);
   U3952 : OAI22_X1 port map( A1 => n17119, A2 => n12326, B1 => n17114, B2 => 
                           n16794, ZN => n9085);
   U3953 : OAI22_X1 port map( A1 => n17312, A2 => n15715, B1 => n17307, B2 => 
                           n16795, ZN => n9101);
   U3954 : OAI22_X1 port map( A1 => n17416, A2 => n15226, B1 => n17411, B2 => 
                           n16796, ZN => n9109);
   U3955 : OAI22_X1 port map( A1 => n17119, A2 => n12327, B1 => n17114, B2 => 
                           n16800, ZN => n9157);
   U3956 : OAI22_X1 port map( A1 => n17312, A2 => n15716, B1 => n17307, B2 => 
                           n16801, ZN => n9173);
   U3957 : OAI22_X1 port map( A1 => n17416, A2 => n15227, B1 => n17411, B2 => 
                           n16802, ZN => n9181);
   U3958 : OAI22_X1 port map( A1 => n17118, A2 => n12328, B1 => n17114, B2 => 
                           n16806, ZN => n9229);
   U3959 : OAI22_X1 port map( A1 => n17311, A2 => n15717, B1 => n17307, B2 => 
                           n16807, ZN => n9245);
   U3960 : OAI22_X1 port map( A1 => n17415, A2 => n15228, B1 => n17411, B2 => 
                           n16808, ZN => n9253);
   U3961 : OAI22_X1 port map( A1 => n17118, A2 => n12329, B1 => n17114, B2 => 
                           n16812, ZN => n9301);
   U3962 : OAI22_X1 port map( A1 => n17311, A2 => n15718, B1 => n17307, B2 => 
                           n16813, ZN => n9317);
   U3963 : OAI22_X1 port map( A1 => n17415, A2 => n15229, B1 => n17411, B2 => 
                           n16814, ZN => n9325);
   U3964 : OAI22_X1 port map( A1 => n17118, A2 => n12330, B1 => n17114, B2 => 
                           n16818, ZN => n9373);
   U3965 : OAI22_X1 port map( A1 => n17311, A2 => n15719, B1 => n17307, B2 => 
                           n16819, ZN => n9389);
   U3966 : OAI22_X1 port map( A1 => n17415, A2 => n15230, B1 => n17411, B2 => 
                           n16820, ZN => n9397);
   U3967 : OAI22_X1 port map( A1 => n17118, A2 => n12331, B1 => n17114, B2 => 
                           n16824, ZN => n9445);
   U3968 : OAI22_X1 port map( A1 => n17311, A2 => n15720, B1 => n17307, B2 => 
                           n16825, ZN => n9461);
   U3969 : OAI22_X1 port map( A1 => n17414, A2 => n15231, B1 => n17411, B2 => 
                           n16826, ZN => n9469);
   U3970 : OAI22_X1 port map( A1 => n17117, A2 => n12332, B1 => n17114, B2 => 
                           n16830, ZN => n9517);
   U3971 : OAI22_X1 port map( A1 => n17310, A2 => n15692, B1 => n17307, B2 => 
                           n16831, ZN => n9533);
   U3972 : OAI22_X1 port map( A1 => n17414, A2 => n15232, B1 => n17411, B2 => 
                           n16832, ZN => n9541);
   U3973 : OAI22_X1 port map( A1 => n17117, A2 => n12333, B1 => n17114, B2 => 
                           n16836, ZN => n9589);
   U3974 : OAI22_X1 port map( A1 => n17310, A2 => n15693, B1 => n17307, B2 => 
                           n16837, ZN => n9605);
   U3975 : OAI22_X1 port map( A1 => n17415, A2 => n15233, B1 => n17411, B2 => 
                           n16838, ZN => n9613);
   U3976 : OAI22_X1 port map( A1 => n17117, A2 => n12334, B1 => n17114, B2 => 
                           n16842, ZN => n9661);
   U3977 : OAI22_X1 port map( A1 => n17310, A2 => n15694, B1 => n17307, B2 => 
                           n16843, ZN => n9677);
   U3978 : OAI22_X1 port map( A1 => n17414, A2 => n15234, B1 => n17411, B2 => 
                           n16844, ZN => n9685);
   U3979 : OAI22_X1 port map( A1 => n17117, A2 => n12335, B1 => n17114, B2 => 
                           n16848, ZN => n9733);
   U3980 : OAI22_X1 port map( A1 => n17310, A2 => n15695, B1 => n17307, B2 => 
                           n16849, ZN => n9749);
   U3981 : OAI22_X1 port map( A1 => n17414, A2 => n15235, B1 => n17411, B2 => 
                           n16850, ZN => n9757);
   U3982 : OAI22_X1 port map( A1 => n17116, A2 => n12336, B1 => n17114, B2 => 
                           n16854, ZN => n9805);
   U3983 : OAI22_X1 port map( A1 => n17309, A2 => n15696, B1 => n17307, B2 => 
                           n16855, ZN => n9821);
   U3984 : OAI22_X1 port map( A1 => n17413, A2 => n15236, B1 => n17411, B2 => 
                           n16856, ZN => n9829);
   U3985 : OAI22_X1 port map( A1 => n17116, A2 => n12337, B1 => n17114, B2 => 
                           n16860, ZN => n9877);
   U3986 : OAI22_X1 port map( A1 => n17309, A2 => n15697, B1 => n17307, B2 => 
                           n16861, ZN => n9893);
   U3987 : OAI22_X1 port map( A1 => n17413, A2 => n15237, B1 => n17411, B2 => 
                           n16862, ZN => n9901);
   U3988 : OAI22_X1 port map( A1 => n17120, A2 => n12339, B1 => n17115, B2 => 
                           n17515, ZN => n9949);
   U3989 : OAI22_X1 port map( A1 => n17313, A2 => n15698, B1 => n17308, B2 => 
                           n17516, ZN => n9965);
   U3990 : OAI22_X1 port map( A1 => n17417, A2 => n15238, B1 => n17412, B2 => 
                           n17517, ZN => n9973);
   U3991 : INV_X1 port map( A => N9926, ZN => n14174);
   U3992 : OAI22_X1 port map( A1 => n16885, A2 => n18031, B1 => n14855, B2 => 
                           n4462, ZN => n10001);
   U3993 : OAI22_X1 port map( A1 => n16895, A2 => n18031, B1 => n15272, B2 => 
                           n4459, ZN => n10002);
   U3994 : OAI22_X1 port map( A1 => n16918, A2 => n18031, B1 => n14065, B2 => 
                           n4451, ZN => n10004);
   U3995 : OAI22_X1 port map( A1 => n16953, A2 => n18031, B1 => n11670, B2 => 
                           n4438, ZN => n10007);
   U3996 : OAI22_X1 port map( A1 => n16964, A2 => n18031, B1 => n14631, B2 => 
                           n4435, ZN => n10008);
   U3997 : OAI22_X1 port map( A1 => n16974, A2 => n18031, B1 => n15275, B2 => 
                           n16966, ZN => n10009);
   U3998 : OAI22_X1 port map( A1 => n16984, A2 => n18031, B1 => n14854, B2 => 
                           n4429, ZN => n10010);
   U3999 : OAI22_X1 port map( A1 => n17007, A2 => n18030, B1 => n14069, B2 => 
                           n16999, ZN => n10012);
   U4000 : OAI22_X1 port map( A1 => n17145, A2 => n18030, B1 => n14628, B2 => 
                           n4382, ZN => n10023);
   U4001 : OAI22_X1 port map( A1 => n17168, A2 => n18029, B1 => n14857, B2 => 
                           n4376, ZN => n10025);
   U4002 : OAI22_X1 port map( A1 => n17179, A2 => n18029, B1 => n11904, B2 => 
                           n4373, ZN => n10026);
   U4003 : OAI22_X1 port map( A1 => n17190, A2 => n18029, B1 => n12197, B2 => 
                           n4370, ZN => n10027);
   U4004 : OAI22_X1 port map( A1 => n17200, A2 => n18029, B1 => n14054, B2 => 
                           n4367, ZN => n10028);
   U4005 : INV_X1 port map( A => N9922, ZN => n14173);
   U4006 : INV_X1 port map( A => n14178, ZN => n14003);
   U4007 : OAI22_X1 port map( A1 => n17944, A2 => n14886, B1 => n17947, B2 => 
                           n17513, ZN => n9923_port);
   U4008 : OAI22_X1 port map( A1 => n17965, A2 => n15269, B1 => n17968, B2 => 
                           n17513, ZN => n9924_port);
   U4009 : OAI22_X1 port map( A1 => n17836, A2 => n14483, B1 => n17840, B2 => 
                           n17512, ZN => n9918);
   U4010 : OAI22_X1 port map( A1 => n17902, A2 => n14644, B1 => n17905, B2 => 
                           n17512, ZN => n9921_port);
   U4011 : OAI22_X1 port map( A1 => n17946, A2 => n14912, B1 => n17959, B2 => 
                           n16448, ZN => n7917);
   U4012 : OAI22_X1 port map( A1 => n17967, A2 => n15244, B1 => n17980, B2 => 
                           n16448, ZN => n7918);
   U4013 : OAI22_X1 port map( A1 => n17925, A2 => n15435, B1 => n17938, B2 => 
                           n16725, ZN => n8266);
   U4014 : OAI22_X1 port map( A1 => n17946, A2 => n14913, B1 => n17958, B2 => 
                           n16725, ZN => n8267);
   U4015 : OAI22_X1 port map( A1 => n17967, A2 => n15246, B1 => n17979, B2 => 
                           n16725, ZN => n8268);
   U4016 : OAI22_X1 port map( A1 => n17925, A2 => n15436, B1 => n17938, B2 => 
                           n16732, ZN => n8338);
   U4017 : OAI22_X1 port map( A1 => n17946, A2 => n14914, B1 => n17959, B2 => 
                           n16732, ZN => n8339);
   U4018 : OAI22_X1 port map( A1 => n17967, A2 => n15247, B1 => n17980, B2 => 
                           n16732, ZN => n8340);
   U4019 : OAI22_X1 port map( A1 => n17925, A2 => n15437, B1 => n17937, B2 => 
                           n16738, ZN => n8410);
   U4020 : OAI22_X1 port map( A1 => n17946, A2 => n14915, B1 => n17957, B2 => 
                           n16738, ZN => n8411);
   U4021 : OAI22_X1 port map( A1 => n17967, A2 => n15248, B1 => n17978, B2 => 
                           n16738, ZN => n8412);
   U4022 : OAI22_X1 port map( A1 => n17925, A2 => n15438, B1 => n17937, B2 => 
                           n16744, ZN => n8482);
   U4023 : OAI22_X1 port map( A1 => n17946, A2 => n14916, B1 => n17958, B2 => 
                           n16744, ZN => n8483);
   U4024 : OAI22_X1 port map( A1 => n17967, A2 => n15249, B1 => n17979, B2 => 
                           n16744, ZN => n8484);
   U4025 : OAI22_X1 port map( A1 => n17924, A2 => n15439, B1 => n17936, B2 => 
                           n16750, ZN => n8554);
   U4026 : OAI22_X1 port map( A1 => n17945, A2 => n14917, B1 => n17956, B2 => 
                           n16750, ZN => n8555);
   U4027 : OAI22_X1 port map( A1 => n17966, A2 => n15250, B1 => n17977, B2 => 
                           n16750, ZN => n8556);
   U4028 : OAI22_X1 port map( A1 => n17924, A2 => n15440, B1 => n17936, B2 => 
                           n16756, ZN => n8626);
   U4029 : OAI22_X1 port map( A1 => n17945, A2 => n14918, B1 => n17957, B2 => 
                           n16756, ZN => n8627);
   U4030 : OAI22_X1 port map( A1 => n17966, A2 => n15251, B1 => n17978, B2 => 
                           n16756, ZN => n8628);
   U4031 : OAI22_X1 port map( A1 => n17924, A2 => n15441, B1 => n17935, B2 => 
                           n16762, ZN => n8698);
   U4032 : OAI22_X1 port map( A1 => n17945, A2 => n14919, B1 => n17955, B2 => 
                           n16762, ZN => n8699);
   U4033 : OAI22_X1 port map( A1 => n17966, A2 => n15252, B1 => n17976, B2 => 
                           n16762, ZN => n8700);
   U4034 : OAI22_X1 port map( A1 => n17924, A2 => n15442, B1 => n17935, B2 => 
                           n16768, ZN => n8770);
   U4035 : OAI22_X1 port map( A1 => n17945, A2 => n14920, B1 => n17956, B2 => 
                           n16768, ZN => n8771);
   U4036 : OAI22_X1 port map( A1 => n17966, A2 => n15253, B1 => n17977, B2 => 
                           n16768, ZN => n8772);
   U4037 : OAI22_X1 port map( A1 => n17924, A2 => n15443, B1 => n17934, B2 => 
                           n16774, ZN => n8842);
   U4038 : OAI22_X1 port map( A1 => n17945, A2 => n14921, B1 => n17955, B2 => 
                           n16774, ZN => n8843);
   U4039 : OAI22_X1 port map( A1 => n17966, A2 => n15254, B1 => n17976, B2 => 
                           n16774, ZN => n8844);
   U4040 : OAI22_X1 port map( A1 => n17924, A2 => n15444, B1 => n17934, B2 => 
                           n16780, ZN => n8914);
   U4041 : OAI22_X1 port map( A1 => n17945, A2 => n14922, B1 => n17954, B2 => 
                           n16780, ZN => n8915);
   U4042 : OAI22_X1 port map( A1 => n17966, A2 => n15255, B1 => n17975, B2 => 
                           n16780, ZN => n8916);
   U4043 : OAI22_X1 port map( A1 => n17924, A2 => n15445, B1 => n17933, B2 => 
                           n16786, ZN => n8986);
   U4044 : OAI22_X1 port map( A1 => n17945, A2 => n14923, B1 => n17954, B2 => 
                           n16786, ZN => n8987);
   U4045 : OAI22_X1 port map( A1 => n17966, A2 => n15256, B1 => n17975, B2 => 
                           n16786, ZN => n8988);
   U4046 : OAI22_X1 port map( A1 => n17924, A2 => n15446, B1 => n17933, B2 => 
                           n16792, ZN => n9058);
   U4047 : OAI22_X1 port map( A1 => n17945, A2 => n14924, B1 => n17953, B2 => 
                           n16792, ZN => n9059);
   U4048 : OAI22_X1 port map( A1 => n17966, A2 => n15257, B1 => n17974, B2 => 
                           n16792, ZN => n9060);
   U4049 : OAI22_X1 port map( A1 => n17924, A2 => n15447, B1 => n17932, B2 => 
                           n16798, ZN => n9130);
   U4050 : OAI22_X1 port map( A1 => n17945, A2 => n14925, B1 => n17953, B2 => 
                           n16798, ZN => n9131);
   U4051 : OAI22_X1 port map( A1 => n17966, A2 => n15258, B1 => n17974, B2 => 
                           n16798, ZN => n9132);
   U4052 : OAI22_X1 port map( A1 => n17924, A2 => n15448, B1 => n17932, B2 => 
                           n16804, ZN => n9202);
   U4053 : OAI22_X1 port map( A1 => n17945, A2 => n14926, B1 => n17952, B2 => 
                           n16804, ZN => n9203);
   U4054 : OAI22_X1 port map( A1 => n17966, A2 => n15259, B1 => n17973, B2 => 
                           n16804, ZN => n9204);
   U4055 : OAI22_X1 port map( A1 => n17924, A2 => n15449, B1 => n17931, B2 => 
                           n16810, ZN => n9274);
   U4056 : OAI22_X1 port map( A1 => n17945, A2 => n14927, B1 => n17952, B2 => 
                           n16810, ZN => n9275);
   U4057 : OAI22_X1 port map( A1 => n17966, A2 => n15260, B1 => n17973, B2 => 
                           n16810, ZN => n9276);
   U4058 : OAI22_X1 port map( A1 => n17924, A2 => n15450, B1 => n17931, B2 => 
                           n16816, ZN => n9346);
   U4059 : OAI22_X1 port map( A1 => n17945, A2 => n14928, B1 => n17951, B2 => 
                           n16816, ZN => n9347);
   U4060 : OAI22_X1 port map( A1 => n17966, A2 => n15261, B1 => n17972, B2 => 
                           n16816, ZN => n9348);
   U4061 : OAI22_X1 port map( A1 => n17924, A2 => n15451, B1 => n17930, B2 => 
                           n16822, ZN => n9418);
   U4062 : OAI22_X1 port map( A1 => n17945, A2 => n14929, B1 => n17951, B2 => 
                           n16822, ZN => n9419);
   U4063 : OAI22_X1 port map( A1 => n17966, A2 => n15262, B1 => n17972, B2 => 
                           n16822, ZN => n9420);
   U4064 : OAI22_X1 port map( A1 => n17923, A2 => n15518, B1 => n17930, B2 => 
                           n16828, ZN => n9490);
   U4065 : OAI22_X1 port map( A1 => n17944, A2 => n14930, B1 => n17950, B2 => 
                           n16828, ZN => n9491);
   U4066 : OAI22_X1 port map( A1 => n17965, A2 => n15263, B1 => n17971, B2 => 
                           n16828, ZN => n9492);
   U4067 : OAI22_X1 port map( A1 => n17923, A2 => n15519, B1 => n17929, B2 => 
                           n16834, ZN => n9562);
   U4068 : OAI22_X1 port map( A1 => n17944, A2 => n14876, B1 => n17950, B2 => 
                           n16834, ZN => n9563);
   U4069 : OAI22_X1 port map( A1 => n17965, A2 => n15264, B1 => n17971, B2 => 
                           n16834, ZN => n9564);
   U4070 : OAI22_X1 port map( A1 => n17923, A2 => n15520, B1 => n17929, B2 => 
                           n16840, ZN => n9634);
   U4071 : OAI22_X1 port map( A1 => n17944, A2 => n14878, B1 => n17949, B2 => 
                           n16840, ZN => n9635);
   U4072 : OAI22_X1 port map( A1 => n17965, A2 => n15265, B1 => n17970, B2 => 
                           n16840, ZN => n9636);
   U4073 : OAI22_X1 port map( A1 => n17923, A2 => n15428, B1 => n17928, B2 => 
                           n16846, ZN => n9706);
   U4074 : OAI22_X1 port map( A1 => n17944, A2 => n14880, B1 => n17949, B2 => 
                           n16846, ZN => n9707);
   U4075 : OAI22_X1 port map( A1 => n17965, A2 => n15266, B1 => n17970, B2 => 
                           n16846, ZN => n9708);
   U4076 : OAI22_X1 port map( A1 => n17923, A2 => n15429, B1 => n17928, B2 => 
                           n16852, ZN => n9778);
   U4077 : OAI22_X1 port map( A1 => n17944, A2 => n14882, B1 => n17948, B2 => 
                           n16852, ZN => n9779);
   U4078 : OAI22_X1 port map( A1 => n17965, A2 => n15267, B1 => n17969, B2 => 
                           n16852, ZN => n9780);
   U4079 : OAI22_X1 port map( A1 => n17923, A2 => n15430, B1 => n17927, B2 => 
                           n16858, ZN => n9850);
   U4080 : OAI22_X1 port map( A1 => n17944, A2 => n14884, B1 => n17948, B2 => 
                           n16858, ZN => n9851);
   U4081 : OAI22_X1 port map( A1 => n17965, A2 => n15268, B1 => n17969, B2 => 
                           n16858, ZN => n9852);
   U4082 : OAI22_X1 port map( A1 => n17923, A2 => n15431, B1 => n17927, B2 => 
                           n17513, ZN => n9922_port);
   U4083 : OAI22_X1 port map( A1 => n17904, A2 => n14645, B1 => n17917, B2 => 
                           n16442, ZN => n7841);
   U4084 : OAI22_X1 port map( A1 => n17838, A2 => n14509, B1 => n17851, B2 => 
                           n16725, ZN => n8262);
   U4085 : OAI22_X1 port map( A1 => n17860, A2 => n15126, B1 => n17873, B2 => 
                           n16725, ZN => n8263);
   U4086 : OAI22_X1 port map( A1 => n17882, A2 => n15637, B1 => n17895, B2 => 
                           n16725, ZN => n8264);
   U4087 : OAI22_X1 port map( A1 => n17904, A2 => n14646, B1 => n17916, B2 => 
                           n16725, ZN => n8265);
   U4088 : OAI22_X1 port map( A1 => n17860, A2 => n15127, B1 => n17873, B2 => 
                           n16731, ZN => n8335);
   U4089 : OAI22_X1 port map( A1 => n17882, A2 => n15638, B1 => n17895, B2 => 
                           n16731, ZN => n8336);
   U4090 : OAI22_X1 port map( A1 => n17904, A2 => n14647, B1 => n17917, B2 => 
                           n16731, ZN => n8337);
   U4091 : OAI22_X1 port map( A1 => n17838, A2 => n14511, B1 => n17848, B2 => 
                           n16737, ZN => n8406);
   U4092 : OAI22_X1 port map( A1 => n17860, A2 => n15128, B1 => n17872, B2 => 
                           n16737, ZN => n8407);
   U4093 : OAI22_X1 port map( A1 => n17882, A2 => n15639, B1 => n17894, B2 => 
                           n16737, ZN => n8408);
   U4094 : OAI22_X1 port map( A1 => n17904, A2 => n14648, B1 => n17915, B2 => 
                           n16737, ZN => n8409);
   U4095 : OAI22_X1 port map( A1 => n17838, A2 => n14512, B1 => n17851, B2 => 
                           n16743, ZN => n8478);
   U4096 : OAI22_X1 port map( A1 => n17860, A2 => n15129, B1 => n17872, B2 => 
                           n16743, ZN => n8479);
   U4097 : OAI22_X1 port map( A1 => n17882, A2 => n15640, B1 => n17894, B2 => 
                           n16743, ZN => n8480);
   U4098 : OAI22_X1 port map( A1 => n17904, A2 => n14649, B1 => n17916, B2 => 
                           n16743, ZN => n8481);
   U4099 : OAI22_X1 port map( A1 => n17837, A2 => n14513, B1 => n17850, B2 => 
                           n16749, ZN => n8550);
   U4100 : OAI22_X1 port map( A1 => n17859, A2 => n15130, B1 => n17871, B2 => 
                           n16749, ZN => n8551);
   U4101 : OAI22_X1 port map( A1 => n17881, A2 => n15641, B1 => n17893, B2 => 
                           n16749, ZN => n8552);
   U4102 : OAI22_X1 port map( A1 => n17903, A2 => n14650, B1 => n17914, B2 => 
                           n16749, ZN => n8553);
   U4103 : OAI22_X1 port map( A1 => n17837, A2 => n14514, B1 => n17850, B2 => 
                           n16755, ZN => n8622);
   U4104 : OAI22_X1 port map( A1 => n17859, A2 => n15131, B1 => n17871, B2 => 
                           n16755, ZN => n8623);
   U4105 : OAI22_X1 port map( A1 => n17881, A2 => n15642, B1 => n17893, B2 => 
                           n16755, ZN => n8624);
   U4106 : OAI22_X1 port map( A1 => n17903, A2 => n14651, B1 => n17915, B2 => 
                           n16755, ZN => n8625);
   U4107 : OAI22_X1 port map( A1 => n17837, A2 => n14515, B1 => n17849, B2 => 
                           n16761, ZN => n8694);
   U4108 : OAI22_X1 port map( A1 => n17859, A2 => n15132, B1 => n17870, B2 => 
                           n16761, ZN => n8695);
   U4109 : OAI22_X1 port map( A1 => n17881, A2 => n15643, B1 => n17892, B2 => 
                           n16761, ZN => n8696);
   U4110 : OAI22_X1 port map( A1 => n17903, A2 => n14652, B1 => n17913, B2 => 
                           n16761, ZN => n8697);
   U4111 : OAI22_X1 port map( A1 => n17837, A2 => n14516, B1 => n17849, B2 => 
                           n16767, ZN => n8766);
   U4112 : OAI22_X1 port map( A1 => n17859, A2 => n15133, B1 => n17870, B2 => 
                           n16767, ZN => n8767);
   U4113 : OAI22_X1 port map( A1 => n17881, A2 => n15644, B1 => n17892, B2 => 
                           n16767, ZN => n8768);
   U4114 : OAI22_X1 port map( A1 => n17903, A2 => n14653, B1 => n17914, B2 => 
                           n16767, ZN => n8769);
   U4115 : OAI22_X1 port map( A1 => n17837, A2 => n14517, B1 => n17847, B2 => 
                           n16773, ZN => n8838);
   U4116 : OAI22_X1 port map( A1 => n17859, A2 => n15134, B1 => n17869, B2 => 
                           n16773, ZN => n8839);
   U4117 : OAI22_X1 port map( A1 => n17881, A2 => n15645, B1 => n17891, B2 => 
                           n16773, ZN => n8840);
   U4118 : OAI22_X1 port map( A1 => n17903, A2 => n14654, B1 => n17913, B2 => 
                           n16773, ZN => n8841);
   U4119 : OAI22_X1 port map( A1 => n17837, A2 => n14518, B1 => n17848, B2 => 
                           n16779, ZN => n8910);
   U4120 : OAI22_X1 port map( A1 => n17859, A2 => n15135, B1 => n17869, B2 => 
                           n16779, ZN => n8911);
   U4121 : OAI22_X1 port map( A1 => n17881, A2 => n15646, B1 => n17891, B2 => 
                           n16779, ZN => n8912);
   U4122 : OAI22_X1 port map( A1 => n17903, A2 => n14655, B1 => n17912, B2 => 
                           n16779, ZN => n8913);
   U4123 : OAI22_X1 port map( A1 => n17837, A2 => n14519, B1 => n17847, B2 => 
                           n16785, ZN => n8982);
   U4124 : OAI22_X1 port map( A1 => n17859, A2 => n15136, B1 => n17868, B2 => 
                           n16785, ZN => n8983);
   U4125 : OAI22_X1 port map( A1 => n17881, A2 => n15647, B1 => n17890, B2 => 
                           n16785, ZN => n8984);
   U4126 : OAI22_X1 port map( A1 => n17903, A2 => n14656, B1 => n17912, B2 => 
                           n16785, ZN => n8985);
   U4127 : OAI22_X1 port map( A1 => n17837, A2 => n14520, B1 => n17846, B2 => 
                           n16791, ZN => n9054);
   U4128 : OAI22_X1 port map( A1 => n17859, A2 => n15137, B1 => n17868, B2 => 
                           n16791, ZN => n9055);
   U4129 : OAI22_X1 port map( A1 => n17881, A2 => n15648, B1 => n17890, B2 => 
                           n16791, ZN => n9056);
   U4130 : OAI22_X1 port map( A1 => n17903, A2 => n14657, B1 => n17911, B2 => 
                           n16791, ZN => n9057);
   U4131 : OAI22_X1 port map( A1 => n17837, A2 => n14521, B1 => n17846, B2 => 
                           n16797, ZN => n9126);
   U4132 : OAI22_X1 port map( A1 => n17859, A2 => n15138, B1 => n17867, B2 => 
                           n16797, ZN => n9127);
   U4133 : OAI22_X1 port map( A1 => n17881, A2 => n15649, B1 => n17889, B2 => 
                           n16797, ZN => n9128);
   U4134 : OAI22_X1 port map( A1 => n17903, A2 => n14658, B1 => n17911, B2 => 
                           n16797, ZN => n9129);
   U4135 : OAI22_X1 port map( A1 => n17837, A2 => n14522, B1 => n17845, B2 => 
                           n16803, ZN => n9198);
   U4136 : OAI22_X1 port map( A1 => n17859, A2 => n15139, B1 => n17867, B2 => 
                           n16803, ZN => n9199);
   U4137 : OAI22_X1 port map( A1 => n17881, A2 => n15650, B1 => n17889, B2 => 
                           n16803, ZN => n9200);
   U4138 : OAI22_X1 port map( A1 => n17903, A2 => n14659, B1 => n17910, B2 => 
                           n16803, ZN => n9201);
   U4139 : OAI22_X1 port map( A1 => n17837, A2 => n14523, B1 => n17845, B2 => 
                           n16809, ZN => n9270);
   U4140 : OAI22_X1 port map( A1 => n17859, A2 => n15140, B1 => n17866, B2 => 
                           n16809, ZN => n9271);
   U4141 : OAI22_X1 port map( A1 => n17881, A2 => n15651, B1 => n17888, B2 => 
                           n16809, ZN => n9272);
   U4142 : OAI22_X1 port map( A1 => n17903, A2 => n14660, B1 => n17910, B2 => 
                           n16809, ZN => n9273);
   U4143 : OAI22_X1 port map( A1 => n17837, A2 => n14524, B1 => n17844, B2 => 
                           n16815, ZN => n9342);
   U4144 : OAI22_X1 port map( A1 => n17859, A2 => n15141, B1 => n17866, B2 => 
                           n16815, ZN => n9343);
   U4145 : OAI22_X1 port map( A1 => n17881, A2 => n15652, B1 => n17888, B2 => 
                           n16815, ZN => n9344);
   U4146 : OAI22_X1 port map( A1 => n17903, A2 => n14661, B1 => n17909, B2 => 
                           n16815, ZN => n9345);
   U4147 : OAI22_X1 port map( A1 => n17837, A2 => n14525, B1 => n17844, B2 => 
                           n16821, ZN => n9414);
   U4148 : OAI22_X1 port map( A1 => n17859, A2 => n15142, B1 => n17865, B2 => 
                           n16821, ZN => n9415);
   U4149 : OAI22_X1 port map( A1 => n17881, A2 => n15653, B1 => n17887, B2 => 
                           n16821, ZN => n9416);
   U4150 : OAI22_X1 port map( A1 => n17903, A2 => n14662, B1 => n17909, B2 => 
                           n16821, ZN => n9417);
   U4151 : OAI22_X1 port map( A1 => n17836, A2 => n14526, B1 => n17843, B2 => 
                           n16827, ZN => n9486);
   U4152 : OAI22_X1 port map( A1 => n17858, A2 => n15143, B1 => n17865, B2 => 
                           n16827, ZN => n9487);
   U4153 : OAI22_X1 port map( A1 => n17880, A2 => n15654, B1 => n17887, B2 => 
                           n16827, ZN => n9488);
   U4154 : OAI22_X1 port map( A1 => n17902, A2 => n14663, B1 => n17908, B2 => 
                           n16827, ZN => n9489);
   U4155 : OAI22_X1 port map( A1 => n17836, A2 => n14478, B1 => n17843, B2 => 
                           n16833, ZN => n9558);
   U4156 : OAI22_X1 port map( A1 => n17858, A2 => n15117, B1 => n17864, B2 => 
                           n16833, ZN => n9559);
   U4157 : OAI22_X1 port map( A1 => n17880, A2 => n15655, B1 => n17886, B2 => 
                           n16833, ZN => n9560);
   U4158 : OAI22_X1 port map( A1 => n17902, A2 => n14664, B1 => n17908, B2 => 
                           n16833, ZN => n9561);
   U4159 : OAI22_X1 port map( A1 => n17836, A2 => n14479, B1 => n17842, B2 => 
                           n16839, ZN => n9630);
   U4160 : OAI22_X1 port map( A1 => n17858, A2 => n15118, B1 => n17864, B2 => 
                           n16839, ZN => n9631);
   U4161 : OAI22_X1 port map( A1 => n17880, A2 => n15656, B1 => n17886, B2 => 
                           n16839, ZN => n9632);
   U4162 : OAI22_X1 port map( A1 => n17902, A2 => n14665, B1 => n17907, B2 => 
                           n16839, ZN => n9633);
   U4163 : OAI22_X1 port map( A1 => n17836, A2 => n14480, B1 => n17842, B2 => 
                           n16845, ZN => n9702);
   U4164 : OAI22_X1 port map( A1 => n17858, A2 => n15119, B1 => n17863, B2 => 
                           n16845, ZN => n9703);
   U4165 : OAI22_X1 port map( A1 => n17880, A2 => n15657, B1 => n17885, B2 => 
                           n16845, ZN => n9704);
   U4166 : OAI22_X1 port map( A1 => n17902, A2 => n14666, B1 => n17907, B2 => 
                           n16845, ZN => n9705);
   U4167 : OAI22_X1 port map( A1 => n17836, A2 => n14481, B1 => n17841, B2 => 
                           n16851, ZN => n9774);
   U4168 : OAI22_X1 port map( A1 => n17858, A2 => n15120, B1 => n17863, B2 => 
                           n16851, ZN => n9775);
   U4169 : OAI22_X1 port map( A1 => n17880, A2 => n15658, B1 => n17885, B2 => 
                           n16851, ZN => n9776);
   U4170 : OAI22_X1 port map( A1 => n17902, A2 => n14667, B1 => n17906, B2 => 
                           n16851, ZN => n9777);
   U4171 : OAI22_X1 port map( A1 => n17836, A2 => n14482, B1 => n17841, B2 => 
                           n16857, ZN => n9846);
   U4172 : OAI22_X1 port map( A1 => n17858, A2 => n15121, B1 => n17862, B2 => 
                           n16857, ZN => n9847);
   U4173 : OAI22_X1 port map( A1 => n17880, A2 => n15659, B1 => n17884, B2 => 
                           n16857, ZN => n9848);
   U4174 : OAI22_X1 port map( A1 => n17902, A2 => n14668, B1 => n17906, B2 => 
                           n16857, ZN => n9849);
   U4175 : OAI22_X1 port map( A1 => n17858, A2 => n15122, B1 => n17862, B2 => 
                           n17512, ZN => n9919);
   U4176 : OAI22_X1 port map( A1 => n17880, A2 => n15660, B1 => n17884, B2 => 
                           n17512, ZN => n9920);
   U4177 : OAI22_X1 port map( A1 => n17944, A2 => n14910, B1 => n17960, B2 => 
                           n16436, ZN => n7767);
   U4178 : OAI22_X1 port map( A1 => n17967, A2 => n15243, B1 => n17981, B2 => 
                           n16442, ZN => n7842);
   U4179 : OAI22_X1 port map( A1 => n17925, A2 => n15434, B1 => n17939, B2 => 
                           n16448, ZN => n7916);
   U4180 : OAI22_X1 port map( A1 => n17858, A2 => n15123, B1 => n17874, B2 => 
                           n16436, ZN => n7765);
   U4181 : OAI22_X1 port map( A1 => n17902, A2 => n14669, B1 => n17918, B2 => 
                           n16436, ZN => n7766);
   U4182 : OAI22_X1 port map( A1 => n17882, A2 => n15661, B1 => n17896, B2 => 
                           n16442, ZN => n7840);
   U4183 : OAI22_X1 port map( A1 => n17838, A2 => n14510, B1 => n17852, B2 => 
                           n16731, ZN => n8334);
   U4184 : OAI22_X1 port map( A1 => n16692, A2 => n18027, B1 => n16693, B2 => 
                           n14860, ZN => n8107);
   U4185 : OAI22_X1 port map( A1 => n16692, A2 => n16702, B1 => n16693, B2 => 
                           n14051, ZN => n8109);
   U4186 : OAI22_X1 port map( A1 => n17577, A2 => n18027, B1 => n17578, B2 => 
                           n14052, ZN => n9985);
   U4187 : OAI22_X1 port map( A1 => n18003, A2 => n18026, B1 => n18005, B2 => 
                           n12048, ZN => n9998);
   U4188 : OAI22_X1 port map( A1 => n18016, A2 => n18026, B1 => n18018, B2 => 
                           n14534, ZN => n9999);
   U4189 : OAI22_X1 port map( A1 => n16934, A2 => n18031, B1 => n14279, B2 => 
                           n16936, ZN => n10006);
   U4190 : OAI22_X1 port map( A1 => n17017, A2 => n18030, B1 => n14871, B2 => 
                           n4420, ZN => n10013);
   U4191 : OAI22_X1 port map( A1 => n17036, A2 => n18030, B1 => n14869, B2 => 
                           n17038, ZN => n10015);
   U4192 : OAI22_X1 port map( A1 => n17049, A2 => n18030, B1 => n14056, B2 => 
                           n17051, ZN => n10016);
   U4193 : OAI22_X1 port map( A1 => n17577, A2 => n16701, B1 => n17578, B2 => 
                           n14856, ZN => n10057);
   U4194 : OAI22_X1 port map( A1 => n17281, A2 => n18029, B1 => n14057, B2 => 
                           n17283, ZN => n10035);
   U4195 : OAI22_X1 port map( A1 => n17294, A2 => n18028, B1 => n14299, B2 => 
                           n17296, ZN => n10036);
   U4196 : OAI22_X1 port map( A1 => n17346, A2 => n18028, B1 => n14870, B2 => 
                           n17348, ZN => n10040);
   U4197 : OAI22_X1 port map( A1 => n17372, A2 => n18028, B1 => n14060, B2 => 
                           n17374, ZN => n10042);
   U4198 : OAI22_X1 port map( A1 => n17398, A2 => n18028, B1 => n14055, B2 => 
                           n17400, ZN => n10044);
   U4199 : OAI22_X1 port map( A1 => n18004, A2 => n16702, B1 => n18005, B2 => 
                           n12049, ZN => n10070);
   U4200 : OAI22_X1 port map( A1 => n18017, A2 => n16702, B1 => n18018, B2 => 
                           n14535, ZN => n10071);
   U4201 : OAI22_X1 port map( A1 => n16877, A2 => n14938, B1 => n16884, B2 => 
                           n16436, ZN => n7770);
   U4202 : OAI22_X1 port map( A1 => n16920, A2 => n15552, B1 => n16927, B2 => 
                           n16436, ZN => n7772);
   U4203 : OAI22_X1 port map( A1 => n16945, A2 => n11951, B1 => n16952, B2 => 
                           n16437, ZN => n7773);
   U4204 : OAI22_X1 port map( A1 => n16966, A2 => n15466, B1 => n16973, B2 => 
                           n16437, ZN => n7774);
   U4205 : OAI22_X1 port map( A1 => n17009, A2 => n15073, B1 => n17016, B2 => 
                           n16437, ZN => n7776);
   U4206 : OAI22_X1 port map( A1 => n17137, A2 => n14678, B1 => n17144, B2 => 
                           n16437, ZN => n7781);
   U4207 : OAI22_X1 port map( A1 => n17160, A2 => n15004, B1 => n17167, B2 => 
                           n16437, ZN => n7782);
   U4208 : OAI22_X1 port map( A1 => n17182, A2 => n12356, B1 => n17189, B2 => 
                           n16437, ZN => n7783);
   U4209 : OAI22_X1 port map( A1 => n17202, A2 => n15181, B1 => n17209, B2 => 
                           n16437, ZN => n7784);
   U4210 : OAI22_X1 port map( A1 => n16877, A2 => n14939, B1 => n16884, B2 => 
                           n16442, ZN => n7845);
   U4211 : OAI22_X1 port map( A1 => n16910, A2 => n14485, B1 => n16917, B2 => 
                           n16442, ZN => n7846);
   U4212 : OAI22_X1 port map( A1 => n16920, A2 => n15553, B1 => n16927, B2 => 
                           n16442, ZN => n7847);
   U4213 : OAI22_X1 port map( A1 => n16956, A2 => n14774, B1 => n16963, B2 => 
                           n16443, ZN => n7848);
   U4214 : OAI22_X1 port map( A1 => n16966, A2 => n15467, B1 => n16973, B2 => 
                           n16443, ZN => n7849);
   U4215 : OAI22_X1 port map( A1 => n16999, A2 => n14429, B1 => n17006, B2 => 
                           n16443, ZN => n7850);
   U4216 : OAI22_X1 port map( A1 => n17009, A2 => n15075, B1 => n17016, B2 => 
                           n16443, ZN => n7851);
   U4217 : OAI22_X1 port map( A1 => n17160, A2 => n15005, B1 => n17167, B2 => 
                           n16443, ZN => n7857);
   U4218 : OAI22_X1 port map( A1 => n17192, A2 => n14301, B1 => n17199, B2 => 
                           n16443, ZN => n7858);
   U4219 : OAI22_X1 port map( A1 => n17202, A2 => n15182, B1 => n17209, B2 => 
                           n16443, ZN => n7859);
   U4220 : OAI22_X1 port map( A1 => n16887, A2 => n15401, B1 => n16894, B2 => 
                           n16448, ZN => n7920);
   U4221 : OAI22_X1 port map( A1 => n16910, A2 => n14486, B1 => n16917, B2 => 
                           n16448, ZN => n7922);
   U4222 : OAI22_X1 port map( A1 => n16920, A2 => n15554, B1 => n16927, B2 => 
                           n16448, ZN => n7923);
   U4223 : OAI22_X1 port map( A1 => n16976, A2 => n14890, B1 => n16983, B2 => 
                           n16449, ZN => n7924);
   U4224 : OAI22_X1 port map( A1 => n16999, A2 => n14431, B1 => n17006, B2 => 
                           n16449, ZN => n7926);
   U4225 : OAI22_X1 port map( A1 => n17009, A2 => n15077, B1 => n17016, B2 => 
                           n16449, ZN => n7927);
   U4226 : OAI22_X1 port map( A1 => n17171, A2 => n12020, B1 => n17178, B2 => 
                           n16449, ZN => n7932);
   U4227 : OAI22_X1 port map( A1 => n17182, A2 => n12360, B1 => n17189, B2 => 
                           n16449, ZN => n7933);
   U4228 : OAI22_X1 port map( A1 => n17192, A2 => n14302, B1 => n17199, B2 => 
                           n16449, ZN => n7934);
   U4229 : OAI22_X1 port map( A1 => n17202, A2 => n15183, B1 => n17209, B2 => 
                           n16449, ZN => n7935);
   U4230 : OAI22_X1 port map( A1 => n16877, A2 => n14941, B1 => n16884, B2 => 
                           n16456, ZN => n7993);
   U4231 : OAI22_X1 port map( A1 => n16887, A2 => n15402, B1 => n16894, B2 => 
                           n16457, ZN => n7994);
   U4232 : OAI22_X1 port map( A1 => n16910, A2 => n14487, B1 => n16917, B2 => 
                           n16457, ZN => n7996);
   U4233 : OAI22_X1 port map( A1 => n16920, A2 => n15555, B1 => n16927, B2 => 
                           n16457, ZN => n7997);
   U4234 : OAI22_X1 port map( A1 => n16944, A2 => n11997, B1 => n16952, B2 => 
                           n16709, ZN => n8119);
   U4235 : OAI22_X1 port map( A1 => n16956, A2 => n14779, B1 => n16963, B2 => 
                           n16709, ZN => n8120);
   U4236 : OAI22_X1 port map( A1 => n16966, A2 => n15469, B1 => n16973, B2 => 
                           n16709, ZN => n8121);
   U4237 : OAI22_X1 port map( A1 => n16976, A2 => n14891, B1 => n16983, B2 => 
                           n16710, ZN => n8122);
   U4238 : OAI22_X1 port map( A1 => n16999, A2 => n14433, B1 => n17006, B2 => 
                           n16710, ZN => n8124);
   U4239 : OAI22_X1 port map( A1 => n17009, A2 => n15079, B1 => n17016, B2 => 
                           n16710, ZN => n8125);
   U4240 : OAI22_X1 port map( A1 => n17137, A2 => n14681, B1 => n17144, B2 => 
                           n16718, ZN => n8199);
   U4241 : OAI22_X1 port map( A1 => n17160, A2 => n15007, B1 => n17167, B2 => 
                           n16718, ZN => n8201);
   U4242 : OAI22_X1 port map( A1 => n17170, A2 => n12021, B1 => n17178, B2 => 
                           n16719, ZN => n8202);
   U4243 : OAI22_X1 port map( A1 => n17182, A2 => n12364, B1 => n17189, B2 => 
                           n16719, ZN => n8203);
   U4244 : OAI22_X1 port map( A1 => n17192, A2 => n14303, B1 => n17199, B2 => 
                           n16719, ZN => n8204);
   U4245 : OAI22_X1 port map( A1 => n17202, A2 => n15184, B1 => n17209, B2 => 
                           n16719, ZN => n8205);
   U4246 : OAI22_X1 port map( A1 => n17062, A2 => n18030, B1 => n14872, B2 => 
                           n17064, ZN => n10017);
   U4247 : OAI22_X1 port map( A1 => n17210, A2 => n18029, B1 => n14873, B2 => 
                           n4362, ZN => n10029);
   U4248 : OAI22_X1 port map( A1 => n17411, A2 => n18028, B1 => n14874, B2 => 
                           n17413, ZN => n10045);
   U4249 : OAI22_X1 port map( A1 => n16877, A2 => n14942, B1 => n16884, B2 => 
                           n16725, ZN => n8273);
   U4250 : OAI22_X1 port map( A1 => n16887, A2 => n15403, B1 => n16894, B2 => 
                           n16726, ZN => n8274);
   U4251 : OAI22_X1 port map( A1 => n16910, A2 => n14488, B1 => n16917, B2 => 
                           n16726, ZN => n8276);
   U4252 : OAI22_X1 port map( A1 => n4448, A2 => n15556, B1 => n16926, B2 => 
                           n16726, ZN => n8277);
   U4253 : OAI22_X1 port map( A1 => n16945, A2 => n11998, B1 => n16952, B2 => 
                           n16726, ZN => n8279);
   U4254 : OAI22_X1 port map( A1 => n16956, A2 => n14782, B1 => n16963, B2 => 
                           n16726, ZN => n8280);
   U4255 : OAI22_X1 port map( A1 => n4432, A2 => n15470, B1 => n16973, B2 => 
                           n16726, ZN => n8281);
   U4256 : OAI22_X1 port map( A1 => n16976, A2 => n14892, B1 => n16983, B2 => 
                           n16726, ZN => n8282);
   U4257 : OAI22_X1 port map( A1 => n4423, A2 => n14436, B1 => n17006, B2 => 
                           n16726, ZN => n8284);
   U4258 : OAI22_X1 port map( A1 => n17009, A2 => n15082, B1 => n17015, B2 => 
                           n16726, ZN => n8285);
   U4259 : OAI22_X1 port map( A1 => n17137, A2 => n14682, B1 => n17144, B2 => 
                           n16727, ZN => n8295);
   U4260 : OAI22_X1 port map( A1 => n17160, A2 => n15008, B1 => n17167, B2 => 
                           n16727, ZN => n8297);
   U4261 : OAI22_X1 port map( A1 => n17171, A2 => n12022, B1 => n17178, B2 => 
                           n16728, ZN => n8298);
   U4262 : OAI22_X1 port map( A1 => n17182, A2 => n12366, B1 => n17189, B2 => 
                           n16728, ZN => n8299);
   U4263 : OAI22_X1 port map( A1 => n17192, A2 => n14304, B1 => n17199, B2 => 
                           n16728, ZN => n8300);
   U4264 : OAI22_X1 port map( A1 => n17202, A2 => n15185, B1 => n17208, B2 => 
                           n16728, ZN => n8301);
   U4265 : OAI22_X1 port map( A1 => n16877, A2 => n14943, B1 => n16883, B2 => 
                           n16732, ZN => n8345);
   U4266 : OAI22_X1 port map( A1 => n16887, A2 => n15404, B1 => n16894, B2 => 
                           n16732, ZN => n8346);
   U4267 : OAI22_X1 port map( A1 => n16910, A2 => n14489, B1 => n16916, B2 => 
                           n16732, ZN => n8348);
   U4268 : OAI22_X1 port map( A1 => n4448, A2 => n15557, B1 => n16926, B2 => 
                           n16732, ZN => n8349);
   U4269 : OAI22_X1 port map( A1 => n16945, A2 => n11999, B1 => n16952, B2 => 
                           n16733, ZN => n8351);
   U4270 : OAI22_X1 port map( A1 => n16956, A2 => n14784, B1 => n16963, B2 => 
                           n16733, ZN => n8352);
   U4271 : OAI22_X1 port map( A1 => n4432, A2 => n15471, B1 => n16972, B2 => 
                           n16733, ZN => n8353);
   U4272 : OAI22_X1 port map( A1 => n16976, A2 => n14893, B1 => n16983, B2 => 
                           n16733, ZN => n8354);
   U4273 : OAI22_X1 port map( A1 => n4423, A2 => n14438, B1 => n17005, B2 => 
                           n16733, ZN => n8356);
   U4274 : OAI22_X1 port map( A1 => n17009, A2 => n15084, B1 => n17015, B2 => 
                           n16733, ZN => n8357);
   U4275 : OAI22_X1 port map( A1 => n17137, A2 => n14683, B1 => n17144, B2 => 
                           n16734, ZN => n8367);
   U4276 : OAI22_X1 port map( A1 => n17160, A2 => n15009, B1 => n17166, B2 => 
                           n16734, ZN => n8369);
   U4277 : OAI22_X1 port map( A1 => n17171, A2 => n12023, B1 => n17178, B2 => 
                           n16734, ZN => n8370);
   U4278 : OAI22_X1 port map( A1 => n17182, A2 => n12368, B1 => n17188, B2 => 
                           n16734, ZN => n8371);
   U4279 : OAI22_X1 port map( A1 => n17192, A2 => n14305, B1 => n17198, B2 => 
                           n16734, ZN => n8372);
   U4280 : OAI22_X1 port map( A1 => n17202, A2 => n15186, B1 => n17208, B2 => 
                           n16734, ZN => n8373);
   U4281 : OAI22_X1 port map( A1 => n16877, A2 => n14944, B1 => n16883, B2 => 
                           n16738, ZN => n8417);
   U4282 : OAI22_X1 port map( A1 => n16887, A2 => n15405, B1 => n16893, B2 => 
                           n16738, ZN => n8418);
   U4283 : OAI22_X1 port map( A1 => n16910, A2 => n14490, B1 => n16916, B2 => 
                           n16738, ZN => n8420);
   U4284 : OAI22_X1 port map( A1 => n4448, A2 => n15558, B1 => n16926, B2 => 
                           n16738, ZN => n8421);
   U4285 : OAI22_X1 port map( A1 => n16945, A2 => n12000, B1 => n16951, B2 => 
                           n16739, ZN => n8423);
   U4286 : OAI22_X1 port map( A1 => n16956, A2 => n14786, B1 => n16962, B2 => 
                           n16739, ZN => n8424);
   U4287 : OAI22_X1 port map( A1 => n4432, A2 => n15472, B1 => n16972, B2 => 
                           n16739, ZN => n8425);
   U4288 : OAI22_X1 port map( A1 => n16976, A2 => n14894, B1 => n16982, B2 => 
                           n16739, ZN => n8426);
   U4289 : OAI22_X1 port map( A1 => n4423, A2 => n14440, B1 => n17005, B2 => 
                           n16739, ZN => n8428);
   U4290 : OAI22_X1 port map( A1 => n17009, A2 => n15086, B1 => n17015, B2 => 
                           n16739, ZN => n8429);
   U4291 : OAI22_X1 port map( A1 => n17137, A2 => n14684, B1 => n17143, B2 => 
                           n16740, ZN => n8439);
   U4292 : OAI22_X1 port map( A1 => n17160, A2 => n15010, B1 => n17166, B2 => 
                           n16740, ZN => n8441);
   U4293 : OAI22_X1 port map( A1 => n17171, A2 => n12024, B1 => n17177, B2 => 
                           n16740, ZN => n8442);
   U4294 : OAI22_X1 port map( A1 => n17182, A2 => n12407, B1 => n17188, B2 => 
                           n16740, ZN => n8443);
   U4295 : OAI22_X1 port map( A1 => n17192, A2 => n14306, B1 => n17198, B2 => 
                           n16740, ZN => n8444);
   U4296 : OAI22_X1 port map( A1 => n17202, A2 => n15187, B1 => n17208, B2 => 
                           n16740, ZN => n8445);
   U4297 : OAI22_X1 port map( A1 => n16877, A2 => n14945, B1 => n16883, B2 => 
                           n16744, ZN => n8489);
   U4298 : OAI22_X1 port map( A1 => n16887, A2 => n15406, B1 => n16893, B2 => 
                           n16744, ZN => n8490);
   U4299 : OAI22_X1 port map( A1 => n16910, A2 => n14491, B1 => n16916, B2 => 
                           n16744, ZN => n8492);
   U4300 : OAI22_X1 port map( A1 => n4448, A2 => n15559, B1 => n16926, B2 => 
                           n16744, ZN => n8493);
   U4301 : OAI22_X1 port map( A1 => n16945, A2 => n12001, B1 => n16951, B2 => 
                           n16745, ZN => n8495);
   U4302 : OAI22_X1 port map( A1 => n16956, A2 => n14788, B1 => n16962, B2 => 
                           n16745, ZN => n8496);
   U4303 : OAI22_X1 port map( A1 => n4432, A2 => n15473, B1 => n16972, B2 => 
                           n16745, ZN => n8497);
   U4304 : OAI22_X1 port map( A1 => n16976, A2 => n14895, B1 => n16982, B2 => 
                           n16745, ZN => n8498);
   U4305 : OAI22_X1 port map( A1 => n4423, A2 => n14442, B1 => n17005, B2 => 
                           n16745, ZN => n8500);
   U4306 : OAI22_X1 port map( A1 => n17009, A2 => n15088, B1 => n17015, B2 => 
                           n16745, ZN => n8501);
   U4307 : OAI22_X1 port map( A1 => n17137, A2 => n14685, B1 => n17143, B2 => 
                           n16746, ZN => n8511);
   U4308 : OAI22_X1 port map( A1 => n17160, A2 => n15011, B1 => n17166, B2 => 
                           n16746, ZN => n8513);
   U4309 : OAI22_X1 port map( A1 => n17171, A2 => n12025, B1 => n17177, B2 => 
                           n16746, ZN => n8514);
   U4310 : OAI22_X1 port map( A1 => n17182, A2 => n12409, B1 => n17188, B2 => 
                           n16746, ZN => n8515);
   U4311 : OAI22_X1 port map( A1 => n17192, A2 => n14307, B1 => n17198, B2 => 
                           n16746, ZN => n8516);
   U4312 : OAI22_X1 port map( A1 => n17202, A2 => n15188, B1 => n17208, B2 => 
                           n16746, ZN => n8517);
   U4313 : OAI22_X1 port map( A1 => n16877, A2 => n14946, B1 => n16883, B2 => 
                           n16750, ZN => n8561);
   U4314 : OAI22_X1 port map( A1 => n16887, A2 => n15407, B1 => n16893, B2 => 
                           n16750, ZN => n8562);
   U4315 : OAI22_X1 port map( A1 => n16910, A2 => n14492, B1 => n16916, B2 => 
                           n16750, ZN => n8564);
   U4316 : OAI22_X1 port map( A1 => n4448, A2 => n15560, B1 => n16925, B2 => 
                           n16750, ZN => n8565);
   U4317 : OAI22_X1 port map( A1 => n16945, A2 => n12002, B1 => n16951, B2 => 
                           n16751, ZN => n8567);
   U4318 : OAI22_X1 port map( A1 => n16956, A2 => n14790, B1 => n16962, B2 => 
                           n16751, ZN => n8568);
   U4319 : OAI22_X1 port map( A1 => n4432, A2 => n15474, B1 => n16972, B2 => 
                           n16751, ZN => n8569);
   U4320 : OAI22_X1 port map( A1 => n16976, A2 => n14896, B1 => n16982, B2 => 
                           n16751, ZN => n8570);
   U4321 : OAI22_X1 port map( A1 => n4423, A2 => n14444, B1 => n17005, B2 => 
                           n16751, ZN => n8572);
   U4322 : OAI22_X1 port map( A1 => n17009, A2 => n15090, B1 => n17014, B2 => 
                           n16751, ZN => n8573);
   U4323 : OAI22_X1 port map( A1 => n17137, A2 => n14686, B1 => n17143, B2 => 
                           n16752, ZN => n8583);
   U4324 : OAI22_X1 port map( A1 => n17160, A2 => n15012, B1 => n17166, B2 => 
                           n16752, ZN => n8585);
   U4325 : OAI22_X1 port map( A1 => n17171, A2 => n12026, B1 => n17177, B2 => 
                           n16752, ZN => n8586);
   U4326 : OAI22_X1 port map( A1 => n17182, A2 => n12411, B1 => n17188, B2 => 
                           n16752, ZN => n8587);
   U4327 : OAI22_X1 port map( A1 => n17192, A2 => n14308, B1 => n17198, B2 => 
                           n16752, ZN => n8588);
   U4328 : OAI22_X1 port map( A1 => n17202, A2 => n15189, B1 => n17207, B2 => 
                           n16752, ZN => n8589);
   U4329 : OAI22_X1 port map( A1 => n16877, A2 => n14947, B1 => n16882, B2 => 
                           n16756, ZN => n8633);
   U4330 : OAI22_X1 port map( A1 => n16887, A2 => n15408, B1 => n16893, B2 => 
                           n16756, ZN => n8634);
   U4331 : OAI22_X1 port map( A1 => n16910, A2 => n14493, B1 => n16915, B2 => 
                           n16756, ZN => n8636);
   U4332 : OAI22_X1 port map( A1 => n4448, A2 => n15561, B1 => n16925, B2 => 
                           n16756, ZN => n8637);
   U4333 : OAI22_X1 port map( A1 => n16945, A2 => n12003, B1 => n16951, B2 => 
                           n16757, ZN => n8639);
   U4334 : OAI22_X1 port map( A1 => n16956, A2 => n14792, B1 => n16962, B2 => 
                           n16757, ZN => n8640);
   U4335 : OAI22_X1 port map( A1 => n4432, A2 => n15475, B1 => n16971, B2 => 
                           n16757, ZN => n8641);
   U4336 : OAI22_X1 port map( A1 => n16976, A2 => n14897, B1 => n16982, B2 => 
                           n16757, ZN => n8642);
   U4337 : OAI22_X1 port map( A1 => n4423, A2 => n14446, B1 => n17004, B2 => 
                           n16757, ZN => n8644);
   U4338 : OAI22_X1 port map( A1 => n17009, A2 => n15092, B1 => n17014, B2 => 
                           n16757, ZN => n8645);
   U4339 : OAI22_X1 port map( A1 => n17137, A2 => n14687, B1 => n17143, B2 => 
                           n16758, ZN => n8655);
   U4340 : OAI22_X1 port map( A1 => n17160, A2 => n15013, B1 => n17165, B2 => 
                           n16758, ZN => n8657);
   U4341 : OAI22_X1 port map( A1 => n17171, A2 => n12027, B1 => n17177, B2 => 
                           n16758, ZN => n8658);
   U4342 : OAI22_X1 port map( A1 => n17182, A2 => n12600, B1 => n17187, B2 => 
                           n16758, ZN => n8659);
   U4343 : OAI22_X1 port map( A1 => n17192, A2 => n14309, B1 => n17197, B2 => 
                           n16758, ZN => n8660);
   U4344 : OAI22_X1 port map( A1 => n17202, A2 => n15190, B1 => n17207, B2 => 
                           n16758, ZN => n8661);
   U4345 : OAI22_X1 port map( A1 => n16877, A2 => n14948, B1 => n16882, B2 => 
                           n16762, ZN => n8705);
   U4346 : OAI22_X1 port map( A1 => n16887, A2 => n15409, B1 => n16892, B2 => 
                           n16762, ZN => n8706);
   U4347 : OAI22_X1 port map( A1 => n16910, A2 => n14494, B1 => n16915, B2 => 
                           n16762, ZN => n8708);
   U4348 : OAI22_X1 port map( A1 => n4448, A2 => n15562, B1 => n16925, B2 => 
                           n16762, ZN => n8709);
   U4349 : OAI22_X1 port map( A1 => n16945, A2 => n12004, B1 => n16950, B2 => 
                           n16763, ZN => n8711);
   U4350 : OAI22_X1 port map( A1 => n16956, A2 => n14794, B1 => n16961, B2 => 
                           n16763, ZN => n8712);
   U4351 : OAI22_X1 port map( A1 => n4432, A2 => n15476, B1 => n16971, B2 => 
                           n16763, ZN => n8713);
   U4352 : OAI22_X1 port map( A1 => n16976, A2 => n14898, B1 => n16981, B2 => 
                           n16763, ZN => n8714);
   U4353 : OAI22_X1 port map( A1 => n4423, A2 => n14448, B1 => n17004, B2 => 
                           n16763, ZN => n8716);
   U4354 : OAI22_X1 port map( A1 => n17009, A2 => n15094, B1 => n17014, B2 => 
                           n16763, ZN => n8717);
   U4355 : OAI22_X1 port map( A1 => n17137, A2 => n14688, B1 => n17142, B2 => 
                           n16764, ZN => n8727);
   U4356 : OAI22_X1 port map( A1 => n17160, A2 => n15014, B1 => n17165, B2 => 
                           n16764, ZN => n8729);
   U4357 : OAI22_X1 port map( A1 => n17171, A2 => n12028, B1 => n17176, B2 => 
                           n16764, ZN => n8730);
   U4358 : OAI22_X1 port map( A1 => n17182, A2 => n12652, B1 => n17187, B2 => 
                           n16764, ZN => n8731);
   U4359 : OAI22_X1 port map( A1 => n17192, A2 => n14310, B1 => n17197, B2 => 
                           n16764, ZN => n8732);
   U4360 : OAI22_X1 port map( A1 => n17202, A2 => n15191, B1 => n17207, B2 => 
                           n16764, ZN => n8733);
   U4361 : OAI22_X1 port map( A1 => n16877, A2 => n14949, B1 => n16882, B2 => 
                           n16768, ZN => n8777);
   U4362 : OAI22_X1 port map( A1 => n16887, A2 => n15410, B1 => n16892, B2 => 
                           n16768, ZN => n8778);
   U4363 : OAI22_X1 port map( A1 => n16910, A2 => n14495, B1 => n16915, B2 => 
                           n16768, ZN => n8780);
   U4364 : OAI22_X1 port map( A1 => n16920, A2 => n15563, B1 => n16924, B2 => 
                           n16768, ZN => n8781);
   U4365 : OAI22_X1 port map( A1 => n16945, A2 => n12005, B1 => n16950, B2 => 
                           n16769, ZN => n8783);
   U4366 : OAI22_X1 port map( A1 => n16956, A2 => n14796, B1 => n16961, B2 => 
                           n16769, ZN => n8784);
   U4367 : OAI22_X1 port map( A1 => n16966, A2 => n15477, B1 => n16971, B2 => 
                           n16769, ZN => n8785);
   U4368 : OAI22_X1 port map( A1 => n16976, A2 => n14899, B1 => n16981, B2 => 
                           n16769, ZN => n8786);
   U4369 : OAI22_X1 port map( A1 => n16999, A2 => n14450, B1 => n17004, B2 => 
                           n16769, ZN => n8788);
   U4370 : OAI22_X1 port map( A1 => n17009, A2 => n15096, B1 => n17013, B2 => 
                           n16769, ZN => n8789);
   U4371 : OAI22_X1 port map( A1 => n17137, A2 => n14689, B1 => n17142, B2 => 
                           n16770, ZN => n8799);
   U4372 : OAI22_X1 port map( A1 => n17160, A2 => n15015, B1 => n17165, B2 => 
                           n16770, ZN => n8801);
   U4373 : OAI22_X1 port map( A1 => n17171, A2 => n12030, B1 => n17176, B2 => 
                           n16770, ZN => n8802);
   U4374 : OAI22_X1 port map( A1 => n17182, A2 => n13996, B1 => n17187, B2 => 
                           n16770, ZN => n8803);
   U4375 : OAI22_X1 port map( A1 => n17192, A2 => n14311, B1 => n17197, B2 => 
                           n16770, ZN => n8804);
   U4376 : OAI22_X1 port map( A1 => n17202, A2 => n15192, B1 => n17206, B2 => 
                           n16770, ZN => n8805);
   U4377 : OAI22_X1 port map( A1 => n16877, A2 => n14950, B1 => n16881, B2 => 
                           n16774, ZN => n8849);
   U4378 : OAI22_X1 port map( A1 => n16887, A2 => n15411, B1 => n16892, B2 => 
                           n16774, ZN => n8850);
   U4379 : OAI22_X1 port map( A1 => n16910, A2 => n14496, B1 => n16914, B2 => 
                           n16774, ZN => n8852);
   U4380 : OAI22_X1 port map( A1 => n4448, A2 => n15564, B1 => n16924, B2 => 
                           n16774, ZN => n8853);
   U4381 : OAI22_X1 port map( A1 => n16945, A2 => n12006, B1 => n16950, B2 => 
                           n16775, ZN => n8855);
   U4382 : OAI22_X1 port map( A1 => n16956, A2 => n14798, B1 => n16961, B2 => 
                           n16775, ZN => n8856);
   U4383 : OAI22_X1 port map( A1 => n4432, A2 => n15478, B1 => n16970, B2 => 
                           n16775, ZN => n8857);
   U4384 : OAI22_X1 port map( A1 => n16976, A2 => n14900, B1 => n16981, B2 => 
                           n16775, ZN => n8858);
   U4385 : OAI22_X1 port map( A1 => n4423, A2 => n14452, B1 => n17003, B2 => 
                           n16775, ZN => n8860);
   U4386 : OAI22_X1 port map( A1 => n17009, A2 => n15098, B1 => n17013, B2 => 
                           n16775, ZN => n8861);
   U4387 : OAI22_X1 port map( A1 => n17137, A2 => n14690, B1 => n17142, B2 => 
                           n16776, ZN => n8871);
   U4388 : OAI22_X1 port map( A1 => n17160, A2 => n15016, B1 => n17164, B2 => 
                           n16776, ZN => n8873);
   U4389 : OAI22_X1 port map( A1 => n17171, A2 => n12031, B1 => n17176, B2 => 
                           n16776, ZN => n8874);
   U4390 : OAI22_X1 port map( A1 => n17182, A2 => n14008, B1 => n17186, B2 => 
                           n16776, ZN => n8875);
   U4391 : OAI22_X1 port map( A1 => n17192, A2 => n14312, B1 => n17196, B2 => 
                           n16776, ZN => n8876);
   U4392 : OAI22_X1 port map( A1 => n17202, A2 => n15193, B1 => n17206, B2 => 
                           n16776, ZN => n8877);
   U4393 : OAI22_X1 port map( A1 => n16877, A2 => n14951, B1 => n16881, B2 => 
                           n16780, ZN => n8921);
   U4394 : OAI22_X1 port map( A1 => n16887, A2 => n15412, B1 => n16891, B2 => 
                           n16780, ZN => n8922);
   U4395 : OAI22_X1 port map( A1 => n16910, A2 => n14497, B1 => n16914, B2 => 
                           n16780, ZN => n8924);
   U4396 : OAI22_X1 port map( A1 => n4448, A2 => n15565, B1 => n16924, B2 => 
                           n16780, ZN => n8925);
   U4397 : OAI22_X1 port map( A1 => n16945, A2 => n12007, B1 => n16949, B2 => 
                           n16781, ZN => n8927);
   U4398 : OAI22_X1 port map( A1 => n16956, A2 => n14800, B1 => n16960, B2 => 
                           n16781, ZN => n8928);
   U4399 : OAI22_X1 port map( A1 => n4432, A2 => n15479, B1 => n16970, B2 => 
                           n16781, ZN => n8929);
   U4400 : OAI22_X1 port map( A1 => n16976, A2 => n14901, B1 => n16980, B2 => 
                           n16781, ZN => n8930);
   U4401 : OAI22_X1 port map( A1 => n4423, A2 => n14454, B1 => n17003, B2 => 
                           n16781, ZN => n8932);
   U4402 : OAI22_X1 port map( A1 => n17009, A2 => n15100, B1 => n17013, B2 => 
                           n16781, ZN => n8933);
   U4403 : OAI22_X1 port map( A1 => n17137, A2 => n14691, B1 => n17141, B2 => 
                           n16782, ZN => n8943);
   U4404 : OAI22_X1 port map( A1 => n17160, A2 => n15017, B1 => n17164, B2 => 
                           n16782, ZN => n8945);
   U4405 : OAI22_X1 port map( A1 => n17171, A2 => n12032, B1 => n17175, B2 => 
                           n16782, ZN => n8946);
   U4406 : OAI22_X1 port map( A1 => n17182, A2 => n14015, B1 => n17186, B2 => 
                           n16782, ZN => n8947);
   U4407 : OAI22_X1 port map( A1 => n17192, A2 => n14313, B1 => n17196, B2 => 
                           n16782, ZN => n8948);
   U4408 : OAI22_X1 port map( A1 => n17202, A2 => n15194, B1 => n17206, B2 => 
                           n16782, ZN => n8949);
   U4409 : OAI22_X1 port map( A1 => n16877, A2 => n14952, B1 => n16881, B2 => 
                           n16786, ZN => n8993);
   U4410 : OAI22_X1 port map( A1 => n16887, A2 => n15413, B1 => n16891, B2 => 
                           n16786, ZN => n8994);
   U4411 : OAI22_X1 port map( A1 => n16910, A2 => n14498, B1 => n16914, B2 => 
                           n16786, ZN => n8996);
   U4412 : OAI22_X1 port map( A1 => n4448, A2 => n15566, B1 => n16924, B2 => 
                           n16786, ZN => n8997);
   U4413 : OAI22_X1 port map( A1 => n16945, A2 => n12008, B1 => n16949, B2 => 
                           n16787, ZN => n8999);
   U4414 : OAI22_X1 port map( A1 => n16956, A2 => n14802, B1 => n16960, B2 => 
                           n16787, ZN => n9000);
   U4415 : OAI22_X1 port map( A1 => n4432, A2 => n15480, B1 => n16970, B2 => 
                           n16787, ZN => n9001);
   U4416 : OAI22_X1 port map( A1 => n16976, A2 => n14902, B1 => n16980, B2 => 
                           n16787, ZN => n9002);
   U4417 : OAI22_X1 port map( A1 => n4423, A2 => n14456, B1 => n17003, B2 => 
                           n16787, ZN => n9004);
   U4418 : OAI22_X1 port map( A1 => n17009, A2 => n15102, B1 => n17013, B2 => 
                           n16787, ZN => n9005);
   U4419 : OAI22_X1 port map( A1 => n17137, A2 => n14692, B1 => n17141, B2 => 
                           n16788, ZN => n9015);
   U4420 : OAI22_X1 port map( A1 => n17160, A2 => n15018, B1 => n17164, B2 => 
                           n16788, ZN => n9017);
   U4421 : OAI22_X1 port map( A1 => n17171, A2 => n12033, B1 => n17175, B2 => 
                           n16788, ZN => n9018);
   U4422 : OAI22_X1 port map( A1 => n17182, A2 => n14035, B1 => n17186, B2 => 
                           n16788, ZN => n9019);
   U4423 : OAI22_X1 port map( A1 => n17192, A2 => n14314, B1 => n17196, B2 => 
                           n16788, ZN => n9020);
   U4424 : OAI22_X1 port map( A1 => n17202, A2 => n15195, B1 => n17206, B2 => 
                           n16788, ZN => n9021);
   U4425 : OAI22_X1 port map( A1 => n16877, A2 => n14953, B1 => n16881, B2 => 
                           n16792, ZN => n9065);
   U4426 : OAI22_X1 port map( A1 => n16887, A2 => n15414, B1 => n16891, B2 => 
                           n16792, ZN => n9066);
   U4427 : OAI22_X1 port map( A1 => n16910, A2 => n14499, B1 => n16914, B2 => 
                           n16792, ZN => n9068);
   U4428 : OAI22_X1 port map( A1 => n16920, A2 => n15567, B1 => n16923, B2 => 
                           n16792, ZN => n9069);
   U4429 : OAI22_X1 port map( A1 => n16945, A2 => n12009, B1 => n16949, B2 => 
                           n16793, ZN => n9071);
   U4430 : OAI22_X1 port map( A1 => n16956, A2 => n14804, B1 => n16960, B2 => 
                           n16793, ZN => n9072);
   U4431 : OAI22_X1 port map( A1 => n16966, A2 => n15481, B1 => n16970, B2 => 
                           n16793, ZN => n9073);
   U4432 : OAI22_X1 port map( A1 => n16976, A2 => n14903, B1 => n16980, B2 => 
                           n16793, ZN => n9074);
   U4433 : OAI22_X1 port map( A1 => n16999, A2 => n14458, B1 => n17003, B2 => 
                           n16793, ZN => n9076);
   U4434 : OAI22_X1 port map( A1 => n17009, A2 => n15104, B1 => n17012, B2 => 
                           n16793, ZN => n9077);
   U4435 : OAI22_X1 port map( A1 => n17137, A2 => n14693, B1 => n17141, B2 => 
                           n16794, ZN => n9087);
   U4436 : OAI22_X1 port map( A1 => n17160, A2 => n15019, B1 => n17164, B2 => 
                           n16794, ZN => n9089);
   U4437 : OAI22_X1 port map( A1 => n17171, A2 => n12034, B1 => n17175, B2 => 
                           n16794, ZN => n9090);
   U4438 : OAI22_X1 port map( A1 => n17182, A2 => n14037, B1 => n17186, B2 => 
                           n16794, ZN => n9091);
   U4439 : OAI22_X1 port map( A1 => n17192, A2 => n14315, B1 => n17196, B2 => 
                           n16794, ZN => n9092);
   U4440 : OAI22_X1 port map( A1 => n17202, A2 => n15196, B1 => n17205, B2 => 
                           n16794, ZN => n9093);
   U4441 : OAI22_X1 port map( A1 => n16877, A2 => n14954, B1 => n16880, B2 => 
                           n16798, ZN => n9137);
   U4442 : OAI22_X1 port map( A1 => n16887, A2 => n15415, B1 => n16891, B2 => 
                           n16798, ZN => n9138);
   U4443 : OAI22_X1 port map( A1 => n16910, A2 => n14500, B1 => n16913, B2 => 
                           n16798, ZN => n9140);
   U4444 : OAI22_X1 port map( A1 => n16920, A2 => n15568, B1 => n16923, B2 => 
                           n16798, ZN => n9141);
   U4445 : OAI22_X1 port map( A1 => n16945, A2 => n12010, B1 => n16949, B2 => 
                           n16799, ZN => n9143);
   U4446 : OAI22_X1 port map( A1 => n16956, A2 => n14806, B1 => n16960, B2 => 
                           n16799, ZN => n9144);
   U4447 : OAI22_X1 port map( A1 => n16966, A2 => n15482, B1 => n16969, B2 => 
                           n16799, ZN => n9145);
   U4448 : OAI22_X1 port map( A1 => n16976, A2 => n14904, B1 => n16980, B2 => 
                           n16799, ZN => n9146);
   U4449 : OAI22_X1 port map( A1 => n16999, A2 => n14460, B1 => n17002, B2 => 
                           n16799, ZN => n9148);
   U4450 : OAI22_X1 port map( A1 => n17009, A2 => n15106, B1 => n17012, B2 => 
                           n16799, ZN => n9149);
   U4451 : OAI22_X1 port map( A1 => n17137, A2 => n14694, B1 => n17141, B2 => 
                           n16800, ZN => n9159);
   U4452 : OAI22_X1 port map( A1 => n17160, A2 => n15020, B1 => n17163, B2 => 
                           n16800, ZN => n9161);
   U4453 : OAI22_X1 port map( A1 => n17171, A2 => n12035, B1 => n17175, B2 => 
                           n16800, ZN => n9162);
   U4454 : OAI22_X1 port map( A1 => n17182, A2 => n14039, B1 => n17185, B2 => 
                           n16800, ZN => n9163);
   U4455 : OAI22_X1 port map( A1 => n17192, A2 => n14316, B1 => n17195, B2 => 
                           n16800, ZN => n9164);
   U4456 : OAI22_X1 port map( A1 => n17202, A2 => n15197, B1 => n17205, B2 => 
                           n16800, ZN => n9165);
   U4457 : OAI22_X1 port map( A1 => n16877, A2 => n14955, B1 => n16880, B2 => 
                           n16804, ZN => n9209);
   U4458 : OAI22_X1 port map( A1 => n16887, A2 => n15416, B1 => n16890, B2 => 
                           n16804, ZN => n9210);
   U4459 : OAI22_X1 port map( A1 => n16910, A2 => n14501, B1 => n16913, B2 => 
                           n16804, ZN => n9212);
   U4460 : OAI22_X1 port map( A1 => n4448, A2 => n15569, B1 => n16923, B2 => 
                           n16804, ZN => n9213);
   U4461 : OAI22_X1 port map( A1 => n16945, A2 => n12011, B1 => n16948, B2 => 
                           n16805, ZN => n9215);
   U4462 : OAI22_X1 port map( A1 => n16956, A2 => n14808, B1 => n16959, B2 => 
                           n16805, ZN => n9216);
   U4463 : OAI22_X1 port map( A1 => n4432, A2 => n15483, B1 => n16969, B2 => 
                           n16805, ZN => n9217);
   U4464 : OAI22_X1 port map( A1 => n16976, A2 => n14905, B1 => n16979, B2 => 
                           n16805, ZN => n9218);
   U4465 : OAI22_X1 port map( A1 => n4423, A2 => n14462, B1 => n17002, B2 => 
                           n16805, ZN => n9220);
   U4466 : OAI22_X1 port map( A1 => n17009, A2 => n15108, B1 => n17012, B2 => 
                           n16805, ZN => n9221);
   U4467 : OAI22_X1 port map( A1 => n17137, A2 => n14695, B1 => n17140, B2 => 
                           n16806, ZN => n9231);
   U4468 : OAI22_X1 port map( A1 => n17160, A2 => n15021, B1 => n17163, B2 => 
                           n16806, ZN => n9233);
   U4469 : OAI22_X1 port map( A1 => n17171, A2 => n12036, B1 => n17174, B2 => 
                           n16806, ZN => n9234);
   U4470 : OAI22_X1 port map( A1 => n17182, A2 => n14041, B1 => n17185, B2 => 
                           n16806, ZN => n9235);
   U4471 : OAI22_X1 port map( A1 => n17192, A2 => n14317, B1 => n17195, B2 => 
                           n16806, ZN => n9236);
   U4472 : OAI22_X1 port map( A1 => n17202, A2 => n15198, B1 => n17205, B2 => 
                           n16806, ZN => n9237);
   U4473 : OAI22_X1 port map( A1 => n4462, A2 => n14956, B1 => n16880, B2 => 
                           n16810, ZN => n9281);
   U4474 : OAI22_X1 port map( A1 => n4459, A2 => n15417, B1 => n16890, B2 => 
                           n16810, ZN => n9282);
   U4475 : OAI22_X1 port map( A1 => n4451, A2 => n14502, B1 => n16913, B2 => 
                           n16810, ZN => n9284);
   U4476 : OAI22_X1 port map( A1 => n16920, A2 => n15570, B1 => n16923, B2 => 
                           n16810, ZN => n9285);
   U4477 : OAI22_X1 port map( A1 => n4438, A2 => n12012, B1 => n16948, B2 => 
                           n16811, ZN => n9287);
   U4478 : OAI22_X1 port map( A1 => n4435, A2 => n14810, B1 => n16959, B2 => 
                           n16811, ZN => n9288);
   U4479 : OAI22_X1 port map( A1 => n16966, A2 => n15484, B1 => n16969, B2 => 
                           n16811, ZN => n9289);
   U4480 : OAI22_X1 port map( A1 => n4429, A2 => n14906, B1 => n16979, B2 => 
                           n16811, ZN => n9290);
   U4481 : OAI22_X1 port map( A1 => n16999, A2 => n14464, B1 => n17002, B2 => 
                           n16811, ZN => n9292);
   U4482 : OAI22_X1 port map( A1 => n4420, A2 => n15110, B1 => n17012, B2 => 
                           n16811, ZN => n9293);
   U4483 : OAI22_X1 port map( A1 => n4382, A2 => n14696, B1 => n17140, B2 => 
                           n16812, ZN => n9303);
   U4484 : OAI22_X1 port map( A1 => n4376, A2 => n15022, B1 => n17163, B2 => 
                           n16812, ZN => n9305);
   U4485 : OAI22_X1 port map( A1 => n4373, A2 => n12037, B1 => n17174, B2 => 
                           n16812, ZN => n9306);
   U4486 : OAI22_X1 port map( A1 => n4370, A2 => n14043, B1 => n17185, B2 => 
                           n16812, ZN => n9307);
   U4487 : OAI22_X1 port map( A1 => n4367, A2 => n14318, B1 => n17195, B2 => 
                           n16812, ZN => n9308);
   U4488 : OAI22_X1 port map( A1 => n4362, A2 => n15199, B1 => n17205, B2 => 
                           n16812, ZN => n9309);
   U4489 : OAI22_X1 port map( A1 => n4462, A2 => n14957, B1 => n16880, B2 => 
                           n16816, ZN => n9353);
   U4490 : OAI22_X1 port map( A1 => n4459, A2 => n15418, B1 => n16890, B2 => 
                           n16816, ZN => n9354);
   U4491 : OAI22_X1 port map( A1 => n4451, A2 => n14503, B1 => n16913, B2 => 
                           n16816, ZN => n9356);
   U4492 : OAI22_X1 port map( A1 => n16920, A2 => n15571, B1 => n16922, B2 => 
                           n16816, ZN => n9357);
   U4493 : OAI22_X1 port map( A1 => n4438, A2 => n12013, B1 => n16948, B2 => 
                           n16817, ZN => n9359);
   U4494 : OAI22_X1 port map( A1 => n4435, A2 => n14812, B1 => n16959, B2 => 
                           n16817, ZN => n9360);
   U4495 : OAI22_X1 port map( A1 => n16966, A2 => n15485, B1 => n16969, B2 => 
                           n16817, ZN => n9361);
   U4496 : OAI22_X1 port map( A1 => n4429, A2 => n14907, B1 => n16979, B2 => 
                           n16817, ZN => n9362);
   U4497 : OAI22_X1 port map( A1 => n16999, A2 => n14466, B1 => n17002, B2 => 
                           n16817, ZN => n9364);
   U4498 : OAI22_X1 port map( A1 => n4420, A2 => n15112, B1 => n17011, B2 => 
                           n16817, ZN => n9365);
   U4499 : OAI22_X1 port map( A1 => n4382, A2 => n14697, B1 => n17140, B2 => 
                           n16818, ZN => n9375);
   U4500 : OAI22_X1 port map( A1 => n4376, A2 => n15023, B1 => n17163, B2 => 
                           n16818, ZN => n9377);
   U4501 : OAI22_X1 port map( A1 => n4373, A2 => n12038, B1 => n17174, B2 => 
                           n16818, ZN => n9378);
   U4502 : OAI22_X1 port map( A1 => n4370, A2 => n14045, B1 => n17185, B2 => 
                           n16818, ZN => n9379);
   U4503 : OAI22_X1 port map( A1 => n4367, A2 => n14319, B1 => n17195, B2 => 
                           n16818, ZN => n9380);
   U4504 : OAI22_X1 port map( A1 => n4362, A2 => n15200, B1 => n17204, B2 => 
                           n16818, ZN => n9381);
   U4505 : OAI22_X1 port map( A1 => n4462, A2 => n14958, B1 => n16879, B2 => 
                           n16822, ZN => n9425);
   U4506 : OAI22_X1 port map( A1 => n4459, A2 => n15419, B1 => n16890, B2 => 
                           n16822, ZN => n9426);
   U4507 : OAI22_X1 port map( A1 => n4451, A2 => n14504, B1 => n16912, B2 => 
                           n16822, ZN => n9428);
   U4508 : OAI22_X1 port map( A1 => n16920, A2 => n15572, B1 => n16922, B2 => 
                           n16822, ZN => n9429);
   U4509 : OAI22_X1 port map( A1 => n4438, A2 => n12014, B1 => n16948, B2 => 
                           n16823, ZN => n9431);
   U4510 : OAI22_X1 port map( A1 => n4435, A2 => n14814, B1 => n16959, B2 => 
                           n16823, ZN => n9432);
   U4511 : OAI22_X1 port map( A1 => n16966, A2 => n15486, B1 => n16968, B2 => 
                           n16823, ZN => n9433);
   U4512 : OAI22_X1 port map( A1 => n4429, A2 => n14908, B1 => n16979, B2 => 
                           n16823, ZN => n9434);
   U4513 : OAI22_X1 port map( A1 => n16999, A2 => n14468, B1 => n17001, B2 => 
                           n16823, ZN => n9436);
   U4514 : OAI22_X1 port map( A1 => n4420, A2 => n15114, B1 => n17011, B2 => 
                           n16823, ZN => n9437);
   U4515 : OAI22_X1 port map( A1 => n4382, A2 => n14698, B1 => n17140, B2 => 
                           n16824, ZN => n9447);
   U4516 : OAI22_X1 port map( A1 => n4376, A2 => n15024, B1 => n17162, B2 => 
                           n16824, ZN => n9449);
   U4517 : OAI22_X1 port map( A1 => n4373, A2 => n12039, B1 => n17174, B2 => 
                           n16824, ZN => n9450);
   U4518 : OAI22_X1 port map( A1 => n4370, A2 => n14047, B1 => n17184, B2 => 
                           n16824, ZN => n9451);
   U4519 : OAI22_X1 port map( A1 => n4367, A2 => n14320, B1 => n17194, B2 => 
                           n16824, ZN => n9452);
   U4520 : OAI22_X1 port map( A1 => n4362, A2 => n15201, B1 => n17204, B2 => 
                           n16824, ZN => n9453);
   U4521 : OAI22_X1 port map( A1 => n4462, A2 => n14959, B1 => n16879, B2 => 
                           n16828, ZN => n9497);
   U4522 : OAI22_X1 port map( A1 => n4459, A2 => n15420, B1 => n16889, B2 => 
                           n16828, ZN => n9498);
   U4523 : OAI22_X1 port map( A1 => n4451, A2 => n14505, B1 => n16912, B2 => 
                           n16828, ZN => n9500);
   U4524 : OAI22_X1 port map( A1 => n16920, A2 => n15573, B1 => n16922, B2 => 
                           n16828, ZN => n9501);
   U4525 : OAI22_X1 port map( A1 => n4438, A2 => n12015, B1 => n16947, B2 => 
                           n16829, ZN => n9503);
   U4526 : OAI22_X1 port map( A1 => n4435, A2 => n14758, B1 => n16958, B2 => 
                           n16829, ZN => n9504);
   U4527 : OAI22_X1 port map( A1 => n16966, A2 => n15459, B1 => n16968, B2 => 
                           n16829, ZN => n9505);
   U4528 : OAI22_X1 port map( A1 => n4429, A2 => n14909, B1 => n16978, B2 => 
                           n16829, ZN => n9506);
   U4529 : OAI22_X1 port map( A1 => n16999, A2 => n14470, B1 => n17001, B2 => 
                           n16829, ZN => n9508);
   U4530 : OAI22_X1 port map( A1 => n4420, A2 => n15116, B1 => n17011, B2 => 
                           n16829, ZN => n9509);
   U4531 : OAI22_X1 port map( A1 => n4382, A2 => n14671, B1 => n17139, B2 => 
                           n16830, ZN => n9519);
   U4532 : OAI22_X1 port map( A1 => n4376, A2 => n15025, B1 => n17162, B2 => 
                           n16830, ZN => n9521);
   U4533 : OAI22_X1 port map( A1 => n4373, A2 => n12040, B1 => n17173, B2 => 
                           n16830, ZN => n9522);
   U4534 : OAI22_X1 port map( A1 => n4370, A2 => n14049, B1 => n17184, B2 => 
                           n16830, ZN => n9523);
   U4535 : OAI22_X1 port map( A1 => n4367, A2 => n14321, B1 => n17194, B2 => 
                           n16830, ZN => n9524);
   U4536 : OAI22_X1 port map( A1 => n4362, A2 => n15202, B1 => n17204, B2 => 
                           n16830, ZN => n9525);
   U4537 : OAI22_X1 port map( A1 => n4462, A2 => n14931, B1 => n16879, B2 => 
                           n16834, ZN => n9569);
   U4538 : OAI22_X1 port map( A1 => n4459, A2 => n15421, B1 => n16889, B2 => 
                           n16834, ZN => n9570);
   U4539 : OAI22_X1 port map( A1 => n4451, A2 => n14471, B1 => n16912, B2 => 
                           n16834, ZN => n9572);
   U4540 : OAI22_X1 port map( A1 => n16920, A2 => n15545, B1 => n16922, B2 => 
                           n16834, ZN => n9573);
   U4541 : OAI22_X1 port map( A1 => n4438, A2 => n11907, B1 => n16947, B2 => 
                           n16835, ZN => n9575);
   U4542 : OAI22_X1 port map( A1 => n4435, A2 => n14760, B1 => n16958, B2 => 
                           n16835, ZN => n9576);
   U4543 : OAI22_X1 port map( A1 => n16966, A2 => n15460, B1 => n16968, B2 => 
                           n16835, ZN => n9577);
   U4544 : OAI22_X1 port map( A1 => n4429, A2 => n14875, B1 => n16978, B2 => 
                           n16835, ZN => n9578);
   U4545 : OAI22_X1 port map( A1 => n16999, A2 => n14527, B1 => n17001, B2 => 
                           n16835, ZN => n9580);
   U4546 : OAI22_X1 port map( A1 => n4420, A2 => n15144, B1 => n17011, B2 => 
                           n16835, ZN => n9581);
   U4547 : OAI22_X1 port map( A1 => n4382, A2 => n14672, B1 => n17139, B2 => 
                           n16836, ZN => n9591);
   U4548 : OAI22_X1 port map( A1 => n4376, A2 => n15026, B1 => n17162, B2 => 
                           n16836, ZN => n9593);
   U4549 : OAI22_X1 port map( A1 => n4373, A2 => n12041, B1 => n17173, B2 => 
                           n16836, ZN => n9594);
   U4550 : OAI22_X1 port map( A1 => n4370, A2 => n12349, B1 => n17184, B2 => 
                           n16836, ZN => n9595);
   U4551 : OAI22_X1 port map( A1 => n4367, A2 => n14322, B1 => n17194, B2 => 
                           n16836, ZN => n9596);
   U4552 : OAI22_X1 port map( A1 => n4362, A2 => n15203, B1 => n17204, B2 => 
                           n16836, ZN => n9597);
   U4553 : OAI22_X1 port map( A1 => n4462, A2 => n14932, B1 => n16878, B2 => 
                           n16840, ZN => n9641_port);
   U4554 : OAI22_X1 port map( A1 => n4459, A2 => n15422, B1 => n16889, B2 => 
                           n16840, ZN => n9642);
   U4555 : OAI22_X1 port map( A1 => n4451, A2 => n14472, B1 => n16912, B2 => 
                           n16840, ZN => n9644);
   U4556 : OAI22_X1 port map( A1 => n16920, A2 => n15546, B1 => n16921, B2 => 
                           n16840, ZN => n9645);
   U4557 : OAI22_X1 port map( A1 => n4438, A2 => n11945, B1 => n16947, B2 => 
                           n16841, ZN => n9647);
   U4558 : OAI22_X1 port map( A1 => n4435, A2 => n14762, B1 => n16958, B2 => 
                           n16841, ZN => n9648);
   U4559 : OAI22_X1 port map( A1 => n16966, A2 => n15461, B1 => n16967, B2 => 
                           n16841, ZN => n9649);
   U4560 : OAI22_X1 port map( A1 => n4429, A2 => n14877, B1 => n16978, B2 => 
                           n16841, ZN => n9650);
   U4561 : OAI22_X1 port map( A1 => n16999, A2 => n14528, B1 => n17001, B2 => 
                           n16841, ZN => n9652);
   U4562 : OAI22_X1 port map( A1 => n4420, A2 => n15145, B1 => n17010, B2 => 
                           n16841, ZN => n9653);
   U4563 : OAI22_X1 port map( A1 => n4382, A2 => n14673, B1 => n17139, B2 => 
                           n16842, ZN => n9663);
   U4564 : OAI22_X1 port map( A1 => n4376, A2 => n15027, B1 => n17161, B2 => 
                           n16842, ZN => n9665);
   U4565 : OAI22_X1 port map( A1 => n4373, A2 => n12042, B1 => n17173, B2 => 
                           n16842, ZN => n9666);
   U4566 : OAI22_X1 port map( A1 => n4370, A2 => n12350, B1 => n17184, B2 => 
                           n16842, ZN => n9667);
   U4567 : OAI22_X1 port map( A1 => n4367, A2 => n14323, B1 => n17194, B2 => 
                           n16842, ZN => n9668);
   U4568 : OAI22_X1 port map( A1 => n4362, A2 => n15204, B1 => n17203, B2 => 
                           n16842, ZN => n9669);
   U4569 : OAI22_X1 port map( A1 => n4462, A2 => n14933, B1 => n16878, B2 => 
                           n16846, ZN => n9713);
   U4570 : OAI22_X1 port map( A1 => n4459, A2 => n15423, B1 => n16889, B2 => 
                           n16846, ZN => n9714);
   U4571 : OAI22_X1 port map( A1 => n4451, A2 => n14473, B1 => n16911, B2 => 
                           n16846, ZN => n9716);
   U4572 : OAI22_X1 port map( A1 => n16920, A2 => n15547, B1 => n16921, B2 => 
                           n16846, ZN => n9717);
   U4573 : OAI22_X1 port map( A1 => n4438, A2 => n11946, B1 => n16947, B2 => 
                           n16847, ZN => n9719);
   U4574 : OAI22_X1 port map( A1 => n4435, A2 => n14764, B1 => n16958, B2 => 
                           n16847, ZN => n9720);
   U4575 : OAI22_X1 port map( A1 => n16966, A2 => n15462, B1 => n16967, B2 => 
                           n16847, ZN => n9721);
   U4576 : OAI22_X1 port map( A1 => n4429, A2 => n14879, B1 => n16978, B2 => 
                           n16847, ZN => n9722);
   U4577 : OAI22_X1 port map( A1 => n16999, A2 => n14529, B1 => n17000, B2 => 
                           n16847, ZN => n9724);
   U4578 : OAI22_X1 port map( A1 => n4420, A2 => n15146, B1 => n17010, B2 => 
                           n16847, ZN => n9725);
   U4579 : OAI22_X1 port map( A1 => n4382, A2 => n14674, B1 => n17139, B2 => 
                           n16848, ZN => n9735);
   U4580 : OAI22_X1 port map( A1 => n4376, A2 => n15028, B1 => n17161, B2 => 
                           n16848, ZN => n9737);
   U4581 : OAI22_X1 port map( A1 => n4373, A2 => n12043, B1 => n17173, B2 => 
                           n16848, ZN => n9738);
   U4582 : OAI22_X1 port map( A1 => n4370, A2 => n12351, B1 => n17183, B2 => 
                           n16848, ZN => n9739);
   U4583 : OAI22_X1 port map( A1 => n4367, A2 => n14324, B1 => n17193, B2 => 
                           n16848, ZN => n9740);
   U4584 : OAI22_X1 port map( A1 => n4362, A2 => n15205, B1 => n17203, B2 => 
                           n16848, ZN => n9741);
   U4585 : OAI22_X1 port map( A1 => n4462, A2 => n14934, B1 => n16879, B2 => 
                           n16852, ZN => n9785);
   U4586 : OAI22_X1 port map( A1 => n4459, A2 => n15424, B1 => n16888, B2 => 
                           n16852, ZN => n9786);
   U4587 : OAI22_X1 port map( A1 => n4451, A2 => n14474, B1 => n16911, B2 => 
                           n16852, ZN => n9788);
   U4588 : OAI22_X1 port map( A1 => n16920, A2 => n15548, B1 => n16921, B2 => 
                           n16852, ZN => n9789);
   U4589 : OAI22_X1 port map( A1 => n4438, A2 => n11947, B1 => n16946, B2 => 
                           n16853, ZN => n9791);
   U4590 : OAI22_X1 port map( A1 => n4435, A2 => n14766, B1 => n16957, B2 => 
                           n16853, ZN => n9792);
   U4591 : OAI22_X1 port map( A1 => n16966, A2 => n15463, B1 => n16968, B2 => 
                           n16853, ZN => n9793);
   U4592 : OAI22_X1 port map( A1 => n4429, A2 => n14881, B1 => n16977, B2 => 
                           n16853, ZN => n9794);
   U4593 : OAI22_X1 port map( A1 => n16999, A2 => n14530, B1 => n17000, B2 => 
                           n16853, ZN => n9796);
   U4594 : OAI22_X1 port map( A1 => n4420, A2 => n15147, B1 => n17010, B2 => 
                           n16853, ZN => n9797);
   U4595 : OAI22_X1 port map( A1 => n4382, A2 => n14675, B1 => n17138, B2 => 
                           n16854, ZN => n9807);
   U4596 : OAI22_X1 port map( A1 => n4376, A2 => n15029, B1 => n17162, B2 => 
                           n16854, ZN => n9809);
   U4597 : OAI22_X1 port map( A1 => n4373, A2 => n12044, B1 => n17172, B2 => 
                           n16854, ZN => n9810);
   U4598 : OAI22_X1 port map( A1 => n4370, A2 => n12352, B1 => n17183, B2 => 
                           n16854, ZN => n9811);
   U4599 : OAI22_X1 port map( A1 => n4367, A2 => n14325, B1 => n17193, B2 => 
                           n16854, ZN => n9812);
   U4600 : OAI22_X1 port map( A1 => n4362, A2 => n15206, B1 => n17203, B2 => 
                           n16854, ZN => n9813);
   U4601 : OAI22_X1 port map( A1 => n4462, A2 => n14935, B1 => n16878, B2 => 
                           n16858, ZN => n9857);
   U4602 : OAI22_X1 port map( A1 => n4459, A2 => n15425, B1 => n16888, B2 => 
                           n16858, ZN => n9858);
   U4603 : OAI22_X1 port map( A1 => n4451, A2 => n14475, B1 => n16911, B2 => 
                           n16858, ZN => n9860);
   U4604 : OAI22_X1 port map( A1 => n16920, A2 => n15549, B1 => n16921, B2 => 
                           n16858, ZN => n9861);
   U4605 : OAI22_X1 port map( A1 => n4438, A2 => n11948, B1 => n16946, B2 => 
                           n16859, ZN => n9863);
   U4606 : OAI22_X1 port map( A1 => n4435, A2 => n14768, B1 => n16957, B2 => 
                           n16859, ZN => n9864);
   U4607 : OAI22_X1 port map( A1 => n16966, A2 => n15464, B1 => n16967, B2 => 
                           n16859, ZN => n9865);
   U4608 : OAI22_X1 port map( A1 => n4429, A2 => n14883, B1 => n16977, B2 => 
                           n16859, ZN => n9866);
   U4609 : OAI22_X1 port map( A1 => n16999, A2 => n14531, B1 => n17000, B2 => 
                           n16859, ZN => n9868);
   U4610 : OAI22_X1 port map( A1 => n4420, A2 => n15148, B1 => n17010, B2 => 
                           n16859, ZN => n9869);
   U4611 : OAI22_X1 port map( A1 => n4382, A2 => n14676, B1 => n17138, B2 => 
                           n16860, ZN => n9879);
   U4612 : OAI22_X1 port map( A1 => n4376, A2 => n15030, B1 => n17161, B2 => 
                           n16860, ZN => n9881);
   U4613 : OAI22_X1 port map( A1 => n4373, A2 => n12045, B1 => n17172, B2 => 
                           n16860, ZN => n9882);
   U4614 : OAI22_X1 port map( A1 => n4370, A2 => n12353, B1 => n17183, B2 => 
                           n16860, ZN => n9883);
   U4615 : OAI22_X1 port map( A1 => n4367, A2 => n14326, B1 => n17193, B2 => 
                           n16860, ZN => n9884);
   U4616 : OAI22_X1 port map( A1 => n4362, A2 => n15207, B1 => n17203, B2 => 
                           n16860, ZN => n9885);
   U4617 : OAI22_X1 port map( A1 => n16877, A2 => n14936, B1 => n16882, B2 => 
                           n17513, ZN => n9929);
   U4618 : OAI22_X1 port map( A1 => n16887, A2 => n15426, B1 => n16892, B2 => 
                           n17513, ZN => n9930);
   U4619 : OAI22_X1 port map( A1 => n16910, A2 => n14476, B1 => n16915, B2 => 
                           n17513, ZN => n9932);
   U4620 : OAI22_X1 port map( A1 => n16920, A2 => n15550, B1 => n16925, B2 => 
                           n17513, ZN => n9933);
   U4621 : OAI22_X1 port map( A1 => n16945, A2 => n11949, B1 => n16950, B2 => 
                           n17514, ZN => n9935);
   U4622 : OAI22_X1 port map( A1 => n16956, A2 => n14770, B1 => n16961, B2 => 
                           n17514, ZN => n9936);
   U4623 : OAI22_X1 port map( A1 => n16966, A2 => n15465, B1 => n16971, B2 => 
                           n17514, ZN => n9937);
   U4624 : OAI22_X1 port map( A1 => n16976, A2 => n14885, B1 => n16981, B2 => 
                           n17514, ZN => n9938);
   U4625 : OAI22_X1 port map( A1 => n16999, A2 => n14532, B1 => n17004, B2 => 
                           n17514, ZN => n9940);
   U4626 : OAI22_X1 port map( A1 => n17009, A2 => n15149, B1 => n17014, B2 => 
                           n17514, ZN => n9941);
   U4627 : OAI22_X1 port map( A1 => n17137, A2 => n14677, B1 => n17142, B2 => 
                           n17515, ZN => n9951);
   U4628 : OAI22_X1 port map( A1 => n17160, A2 => n15031, B1 => n17165, B2 => 
                           n17515, ZN => n9953);
   U4629 : OAI22_X1 port map( A1 => n17171, A2 => n12046, B1 => n17176, B2 => 
                           n17515, ZN => n9954);
   U4630 : OAI22_X1 port map( A1 => n17182, A2 => n12354, B1 => n17187, B2 => 
                           n17515, ZN => n9955);
   U4631 : OAI22_X1 port map( A1 => n17192, A2 => n14327, B1 => n17197, B2 => 
                           n17515, ZN => n9956);
   U4632 : OAI22_X1 port map( A1 => n17202, A2 => n15208, B1 => n17207, B2 => 
                           n17515, ZN => n9957);
   U4633 : OAI22_X1 port map( A1 => n16928, A2 => n18031, B1 => n15277, B2 => 
                           n16920, ZN => n10005);
   U4634 : OAI22_X1 port map( A1 => n17023, A2 => n18030, B1 => n12160, B2 => 
                           n17025, ZN => n10014);
   U4635 : OAI22_X1 port map( A1 => n17075, A2 => n18030, B1 => n15278, B2 => 
                           n17077, ZN => n10018);
   U4636 : OAI22_X1 port map( A1 => n17088, A2 => n18030, B1 => n15276, B2 => 
                           n17090, ZN => n10019);
   U4637 : OAI22_X1 port map( A1 => n17101, A2 => n18030, B1 => n11498, B2 => 
                           n17103, ZN => n10020);
   U4638 : OAI22_X1 port map( A1 => n17114, A2 => n18030, B1 => n12163, B2 => 
                           n17116, ZN => n10021);
   U4639 : OAI22_X1 port map( A1 => n17127, A2 => n18030, B1 => n15282, B2 => 
                           n17129, ZN => n10022);
   U4640 : OAI22_X1 port map( A1 => n17229, A2 => n18029, B1 => n15273, B2 => 
                           n17231, ZN => n10031);
   U4641 : OAI22_X1 port map( A1 => n17242, A2 => n18029, B1 => n12161, B2 => 
                           n17244, ZN => n10032);
   U4642 : OAI22_X1 port map( A1 => n17255, A2 => n18029, B1 => n14822, B2 => 
                           n17257, ZN => n10033);
   U4643 : OAI22_X1 port map( A1 => n17307, A2 => n18028, B1 => n15281, B2 => 
                           n17309, ZN => n10037);
   U4644 : OAI22_X1 port map( A1 => n17320, A2 => n18028, B1 => n15270, B2 => 
                           n17322, ZN => n10038);
   U4645 : OAI22_X1 port map( A1 => n17333, A2 => n18028, B1 => n11541, B2 => 
                           n17335, ZN => n10039);
   U4646 : OAI22_X1 port map( A1 => n17359, A2 => n18028, B1 => n15280, B2 => 
                           n17361, ZN => n10041);
   U4647 : OAI22_X1 port map( A1 => n17385, A2 => n18028, B1 => n14629, B2 => 
                           n17387, ZN => n10043);
   U4648 : OAI22_X1 port map( A1 => n17424, A2 => n18028, B1 => n15271, B2 => 
                           n17426, ZN => n10046);
   U4649 : OAI22_X1 port map( A1 => n17437, A2 => n18028, B1 => n12196, B2 => 
                           n17439, ZN => n10047);
   U4650 : OAI22_X1 port map( A1 => n17451, A2 => n18027, B1 => n14632, B2 => 
                           n17452, ZN => n10048);
   U4651 : OAI22_X1 port map( A1 => n17463, A2 => n18027, B1 => n15274, B2 => 
                           n17465, ZN => n10049);
   U4652 : OAI22_X1 port map( A1 => n17476, A2 => n18027, B1 => n15283, B2 => 
                           n17478, ZN => n10050);
   U4653 : OAI22_X1 port map( A1 => n17489, A2 => n18027, B1 => n14630, B2 => 
                           n17491, ZN => n10051);
   U4654 : OAI22_X1 port map( A1 => n17502, A2 => n18027, B1 => n15279, B2 => 
                           n17504, ZN => n10052);
   U4655 : OAI22_X1 port map( A1 => n4462, A2 => n14937, B1 => n16885, B2 => 
                           n16706, ZN => n10073);
   U4656 : OAI22_X1 port map( A1 => n4459, A2 => n15427, B1 => n16895, B2 => 
                           n16706, ZN => n10074);
   U4657 : OAI22_X1 port map( A1 => n4451, A2 => n14477, B1 => n16918, B2 => 
                           n16706, ZN => n10076);
   U4658 : OAI22_X1 port map( A1 => n16920, A2 => n15551, B1 => n16928, B2 => 
                           n16706, ZN => n10077);
   U4659 : OAI22_X1 port map( A1 => n4438, A2 => n11950, B1 => n16953, B2 => 
                           n16706, ZN => n10079);
   U4660 : OAI22_X1 port map( A1 => n4435, A2 => n14816, B1 => n16964, B2 => 
                           n16706, ZN => n10080);
   U4661 : OAI22_X1 port map( A1 => n16966, A2 => n15487, B1 => n16974, B2 => 
                           n16706, ZN => n10081);
   U4662 : OAI22_X1 port map( A1 => n16976, A2 => n14887, B1 => n16984, B2 => 
                           n16706, ZN => n10082);
   U4663 : OAI22_X1 port map( A1 => n16999, A2 => n14533, B1 => n17007, B2 => 
                           n16705, ZN => n10084);
   U4664 : OAI22_X1 port map( A1 => n17009, A2 => n15150, B1 => n17017, B2 => 
                           n16705, ZN => n10085);
   U4665 : OAI22_X1 port map( A1 => n17137, A2 => n14699, B1 => n17145, B2 => 
                           n16705, ZN => n10095);
   U4666 : OAI22_X1 port map( A1 => n17160, A2 => n15032, B1 => n17168, B2 => 
                           n16704, ZN => n10097);
   U4667 : OAI22_X1 port map( A1 => n17170, A2 => n12047, B1 => n17179, B2 => 
                           n16704, ZN => n10098);
   U4668 : OAI22_X1 port map( A1 => n17182, A2 => n12355, B1 => n17190, B2 => 
                           n16704, ZN => n10099);
   U4669 : OAI22_X1 port map( A1 => n17192, A2 => n14328, B1 => n17200, B2 => 
                           n16704, ZN => n10100);
   U4670 : OAI22_X1 port map( A1 => n17202, A2 => n15209, B1 => n17210, B2 => 
                           n16704, ZN => n10101);
   U4671 : INV_X1 port map( A => N46298, ZN => n13978);
   U4672 : INV_X1 port map( A => N45784, ZN => n12497);
   U4673 : NAND2_X1 port map( A1 => n14091, A2 => n14149, ZN => n4175);
   U4674 : NAND2_X1 port map( A1 => n14091, A2 => n14150, ZN => n4186);
   U4675 : NAND2_X1 port map( A1 => n14140, A2 => n14196, ZN => n14120);
   U4676 : NAND2_X1 port map( A1 => n14128, A2 => n14196, ZN => n14166);
   U4677 : NAND2_X1 port map( A1 => n14146, A2 => n14196, ZN => n14163);
   U4678 : NOR2_X1 port map( A1 => n13973, A2 => n13974, ZN => n12624);
   U4679 : NAND2_X1 port map( A1 => n14137, A2 => n14020, ZN => n14117);
   U4680 : NAND2_X1 port map( A1 => n14202, A2 => n14020, ZN => n14125);
   U4681 : NAND2_X1 port map( A1 => n14138, A2 => n14020, ZN => n14123);
   U4682 : NAND2_X1 port map( A1 => n14143, A2 => n14020, ZN => n14160);
   U4683 : NAND2_X1 port map( A1 => n14150, A2 => n14151, ZN => n4173);
   U4684 : NAND2_X1 port map( A1 => n14149, A2 => n14151, ZN => n4242);
   U4685 : NAND2_X1 port map( A1 => datain(0), A2 => n18039, ZN => n12338);
   U4686 : NAND2_X1 port map( A1 => datain(1), A2 => n18039, ZN => n12184);
   U4687 : NAND2_X1 port map( A1 => datain(2), A2 => n18039, ZN => n12029);
   U4688 : NOR2_X1 port map( A1 => n18050, A2 => n14006, ZN => n4090);
   U4689 : OR2_X1 port map( A1 => n14144, A2 => n14020, ZN => n14124);
   U4690 : AND2_X1 port map( A1 => n14143, A2 => N9925, ZN => n14108);
   U4691 : NAND2_X1 port map( A1 => n14130, A2 => n14146, ZN => n14136);
   U4692 : INV_X1 port map( A => N46299, ZN => n13979);
   U4693 : INV_X1 port map( A => N45785, ZN => n12498);
   U4694 : INV_X1 port map( A => N276, ZN => n14234);
   U4695 : AND2_X1 port map( A1 => n14094, A2 => n14105, ZN => n4123);
   U4696 : AND2_X1 port map( A1 => n14104, A2 => n14105, ZN => n4124);
   U4697 : AND2_X1 port map( A1 => n14108, A2 => n14105, ZN => n4130);
   U4698 : AND2_X1 port map( A1 => n14107, A2 => n14105, ZN => n4131);
   U4699 : INV_X1 port map( A => n14263, ZN => n14262);
   U4700 : AND2_X1 port map( A1 => n14194, A2 => n14178, ZN => n14170);
   U4701 : INV_X1 port map( A => n14146, ZN => n14172);
   U4702 : NAND2_X1 port map( A1 => n13903, A2 => n13901, ZN => n12522);
   U4703 : NAND2_X1 port map( A1 => n12422, A2 => n12420, ZN => n10519);
   U4704 : NAND2_X1 port map( A1 => n13901, A2 => n13902, ZN => n12523);
   U4705 : NAND2_X1 port map( A1 => n12420, A2 => n12421, ZN => n10520);
   U4706 : AND2_X1 port map( A1 => n14091, A2 => n14152, ZN => n4170);
   U4707 : AND2_X1 port map( A1 => n14091, A2 => n14092, ZN => n4107);
   U4708 : AND2_X1 port map( A1 => N9921, A2 => n14209, ZN => n14137);
   U4709 : AND2_X1 port map( A1 => n14152, A2 => n14151, ZN => n4171);
   U4710 : OAI21_X1 port map( B1 => n18051, B2 => n14821, A => n13997, ZN => 
                           n10185);
   U4711 : AND2_X1 port map( A1 => N9923, A2 => N9921, ZN => n14143);
   U4712 : NAND2_X1 port map( A1 => datain(4), A2 => n18038, ZN => n10425);
   U4713 : AND2_X1 port map( A1 => n13904, A2 => n13985, ZN => n12524);
   U4714 : AND2_X1 port map( A1 => n13904, A2 => n13902, ZN => n12525);
   U4715 : AND2_X1 port map( A1 => n12423, A2 => n12421, ZN => n10523);
   U4716 : AND2_X1 port map( A1 => n12423, A2 => n12504, ZN => n10522);
   U4717 : AND2_X1 port map( A1 => n13903, A2 => n13904, ZN => n12520);
   U4718 : AND2_X1 port map( A1 => n13905, A2 => n13904, ZN => n12634);
   U4719 : AND2_X1 port map( A1 => n12422, A2 => n12423, ZN => n10517);
   U4720 : AND2_X1 port map( A1 => n12424, A2 => n12423, ZN => n10663);
   U4721 : AND2_X1 port map( A1 => n13901, A2 => n13985, ZN => n12633);
   U4722 : AND2_X1 port map( A1 => n12420, A2 => n12504, ZN => n10662);
   U4723 : AND2_X1 port map( A1 => n13905, A2 => n13901, ZN => n12519);
   U4724 : AND2_X1 port map( A1 => n12424, A2 => n12420, ZN => n10516);
   U4725 : NAND2_X1 port map( A1 => n12492, A2 => n12507, ZN => n12500);
   U4726 : INV_X1 port map( A => n12493, ZN => n12507);
   U4727 : BUF_X1 port map( A => reset, Z => n18032);
   U4728 : NAND2_X1 port map( A1 => n13973, A2 => n13988, ZN => n13981);
   U4729 : INV_X1 port map( A => n13974, ZN => n13988);
   U4730 : INV_X1 port map( A => N9923, ZN => n14209);
   U4731 : INV_X1 port map( A => n14114, ZN => n4150);
   U4732 : OAI22_X1 port map( A1 => n14115, A2 => n14116, B1 => n14117, B2 => 
                           n14118, ZN => n14114);
   U4733 : INV_X1 port map( A => N46300, ZN => n13976);
   U4734 : INV_X1 port map( A => N45786, ZN => n12495);
   U4735 : INV_X1 port map( A => N274, ZN => n14259);
   U4736 : INV_X1 port map( A => N46301, ZN => n13975);
   U4737 : INV_X1 port map( A => N45787, ZN => n12494);
   U4738 : INV_X1 port map( A => N275, ZN => n14257);
   U4739 : INV_X1 port map( A => n14119, ZN => n4148);
   U4740 : OAI22_X1 port map( A1 => n14120, A2 => n14115, B1 => n14121, B2 => 
                           n14117, ZN => n14119);
   U4741 : INV_X1 port map( A => n14195, ZN => n4222);
   U4742 : OAI22_X1 port map( A1 => n14166, A2 => n14115, B1 => n14167, B2 => 
                           n14117, ZN => n14195);
   U4743 : NAND2_X1 port map( A1 => datain(5), A2 => n18038, ZN => n10315);
   U4744 : AND2_X1 port map( A1 => n14147, A2 => n14820, ZN => n14130);
   U4745 : INV_X1 port map( A => n14128, ZN => n14100);
   U4746 : NAND2_X1 port map( A1 => datain(3), A2 => n18038, ZN => n11868);
   U4747 : INV_X1 port map( A => N46303, ZN => n13963);
   U4748 : INV_X1 port map( A => N45789, ZN => n12482);
   U4749 : INV_X1 port map( A => add_73_carry_5_port, ZN => n14265);
   U4750 : INV_X1 port map( A => n14006, ZN => n14233);
   U4751 : INV_X1 port map( A => n14247, ZN => n14239);
   U4752 : INV_X1 port map( A => n14149, ZN => n14186);
   U4753 : INV_X1 port map( A => n14150, ZN => n14184);
   U4754 : INV_X1 port map( A => N45788, ZN => n12499);
   U4755 : INV_X1 port map( A => N46302, ZN => n13980);
   U4756 : NOR2_X1 port map( A1 => N9908, A2 => n14022, ZN => n14017);
   U4757 : NOR2_X1 port map( A1 => n18050, A2 => datain(0), ZN => n12302);
   U4758 : NOR2_X1 port map( A1 => n18050, A2 => datain(1), ZN => n12149);
   U4759 : NOR2_X1 port map( A1 => n18050, A2 => datain(2), ZN => n11996);
   U4760 : INV_X1 port map( A => datain(4), ZN => n10400);
   U4761 : INV_X1 port map( A => datain(5), ZN => n10290);
   U4762 : INV_X1 port map( A => datain(6), ZN => n10285);
   U4763 : INV_X1 port map( A => datain(3), ZN => n11843);
   U4764 : AOI221_X1 port map( B1 => registers_56_1_port, B2 => n16517, C1 => 
                           registers_60_1_port, C2 => n16514, A => n12297, ZN 
                           => n12296);
   U4765 : OAI222_X1 port map( A1 => n16511, A2 => n14570, B1 => n16508, B2 => 
                           n12052, C1 => n16505, C2 => n15243, ZN => n12297);
   U4766 : AOI221_X1 port map( B1 => registers_56_2_port, B2 => n16517, C1 => 
                           registers_60_2_port, C2 => n16514, A => n12144, ZN 
                           => n12143);
   U4767 : OAI222_X1 port map( A1 => n16511, A2 => n14571, B1 => n16508, B2 => 
                           n12053, C1 => n16505, C2 => n15244, ZN => n12144);
   U4768 : AOI221_X1 port map( B1 => registers_56_3_port, B2 => n16517, C1 => 
                           registers_60_3_port, C2 => n16514, A => n11991, ZN 
                           => n11990);
   U4769 : OAI222_X1 port map( A1 => n16511, A2 => n14572, B1 => n16508, B2 => 
                           n12054, C1 => n16505, C2 => n15240, ZN => n11991);
   U4770 : NOR2_X1 port map( A1 => N9910, A2 => n10189, ZN => n14140);
   U4771 : AOI221_X1 port map( B1 => registers_2_0_port, B2 => n16364, C1 => 
                           registers_29_0_port, C2 => n16361, A => n13942, ZN 
                           => n13941);
   U4772 : OAI222_X1 port map( A1 => n16358, A2 => n15004, B1 => n16355, B2 => 
                           n14300, C1 => n16352, C2 => n12018, ZN => n13942);
   U4773 : AOI221_X1 port map( B1 => registers_56_0_port, B2 => n16265, C1 => 
                           registers_60_0_port, C2 => n16262, A => n13968, ZN 
                           => n13967);
   U4774 : OAI222_X1 port map( A1 => n16259, A2 => n14573, B1 => n16256, B2 => 
                           n12055, C1 => n16253, C2 => n15245, ZN => n13968);
   U4775 : AOI221_X1 port map( B1 => registers_2_1_port, B2 => n16364, C1 => 
                           registers_29_1_port, C2 => n16361, A => n13877, ZN 
                           => n13876);
   U4776 : OAI222_X1 port map( A1 => n16358, A2 => n15005, B1 => n16355, B2 => 
                           n14301, C1 => n16352, C2 => n12019, ZN => n13877);
   U4777 : AOI221_X1 port map( B1 => registers_56_1_port, B2 => n16265, C1 => 
                           registers_60_1_port, C2 => n16262, A => n13893, ZN 
                           => n13892);
   U4778 : OAI222_X1 port map( A1 => n16259, A2 => n14570, B1 => n16256, B2 => 
                           n12052, C1 => n16253, C2 => n15243, ZN => n13893);
   U4779 : AOI221_X1 port map( B1 => registers_2_2_port, B2 => n16364, C1 => 
                           registers_29_2_port, C2 => n16361, A => n13835, ZN 
                           => n13834);
   U4780 : OAI222_X1 port map( A1 => n16358, A2 => n15006, B1 => n16355, B2 => 
                           n14302, C1 => n16352, C2 => n12020, ZN => n13835);
   U4781 : AOI221_X1 port map( B1 => registers_56_2_port, B2 => n16265, C1 => 
                           registers_60_2_port, C2 => n16262, A => n13851, ZN 
                           => n13850);
   U4782 : OAI222_X1 port map( A1 => n16259, A2 => n14571, B1 => n16256, B2 => 
                           n12053, C1 => n16253, C2 => n15244, ZN => n13851);
   U4783 : AOI221_X1 port map( B1 => registers_2_3_port, B2 => n16364, C1 => 
                           registers_29_3_port, C2 => n16361, A => n13793, ZN 
                           => n13792);
   U4784 : OAI222_X1 port map( A1 => n16358, A2 => n14989, B1 => n16355, B2 => 
                           n14282, C1 => n16352, C2 => n12016, ZN => n13793);
   U4785 : AOI221_X1 port map( B1 => registers_56_3_port, B2 => n16265, C1 => 
                           registers_60_3_port, C2 => n16262, A => n13809, ZN 
                           => n13808);
   U4786 : OAI222_X1 port map( A1 => n16259, A2 => n14572, B1 => n16256, B2 => 
                           n12054, C1 => n16253, C2 => n15240, ZN => n13809);
   U4787 : AOI221_X1 port map( B1 => registers_2_4_port, B2 => n16364, C1 => 
                           registers_29_4_port, C2 => n16361, A => n13751, ZN 
                           => n13750);
   U4788 : OAI222_X1 port map( A1 => n16358, A2 => n14990, B1 => n16355, B2 => 
                           n14283, C1 => n16352, C2 => n12017, ZN => n13751);
   U4789 : AOI221_X1 port map( B1 => registers_56_4_port, B2 => n16265, C1 => 
                           registers_60_4_port, C2 => n16262, A => n13767, ZN 
                           => n13766);
   U4790 : OAI222_X1 port map( A1 => n16259, A2 => n14538, B1 => n16256, B2 => 
                           n12050, C1 => n16253, C2 => n15241, ZN => n13767);
   U4791 : AOI221_X1 port map( B1 => registers_2_5_port, B2 => n16364, C1 => 
                           registers_29_5_port, C2 => n16361, A => n13709, ZN 
                           => n13708);
   U4792 : OAI222_X1 port map( A1 => n16358, A2 => n15007, B1 => n16355, B2 => 
                           n14303, C1 => n16352, C2 => n12021, ZN => n13709);
   U4793 : AOI221_X1 port map( B1 => registers_56_5_port, B2 => n16265, C1 => 
                           registers_60_5_port, C2 => n16262, A => n13725, ZN 
                           => n13724);
   U4794 : OAI222_X1 port map( A1 => n16259, A2 => n14539, B1 => n16256, B2 => 
                           n12051, C1 => n16253, C2 => n15242, ZN => n13725);
   U4795 : AOI221_X1 port map( B1 => registers_2_6_port, B2 => n16364, C1 => 
                           registers_29_6_port, C2 => n16361, A => n13667, ZN 
                           => n13666);
   U4796 : OAI222_X1 port map( A1 => n16358, A2 => n15008, B1 => n16355, B2 => 
                           n14304, C1 => n16352, C2 => n12022, ZN => n13667);
   U4797 : AOI221_X1 port map( B1 => registers_56_6_port, B2 => n16265, C1 => 
                           registers_60_6_port, C2 => n16262, A => n13683, ZN 
                           => n13682);
   U4798 : OAI222_X1 port map( A1 => n16259, A2 => n14574, B1 => n16256, B2 => 
                           n12056, C1 => n16253, C2 => n15246, ZN => n13683);
   U4799 : AOI221_X1 port map( B1 => registers_2_7_port, B2 => n16364, C1 => 
                           registers_29_7_port, C2 => n16361, A => n13625, ZN 
                           => n13624);
   U4800 : OAI222_X1 port map( A1 => n16358, A2 => n15009, B1 => n16355, B2 => 
                           n14305, C1 => n16352, C2 => n12023, ZN => n13625);
   U4801 : AOI221_X1 port map( B1 => registers_56_7_port, B2 => n16265, C1 => 
                           registers_60_7_port, C2 => n16262, A => n13641, ZN 
                           => n13640);
   U4802 : OAI222_X1 port map( A1 => n16259, A2 => n14575, B1 => n16256, B2 => 
                           n12057, C1 => n16253, C2 => n15247, ZN => n13641);
   U4803 : AOI221_X1 port map( B1 => registers_2_8_port, B2 => n16364, C1 => 
                           registers_29_8_port, C2 => n16361, A => n13583, ZN 
                           => n13582);
   U4804 : OAI222_X1 port map( A1 => n16358, A2 => n15010, B1 => n16355, B2 => 
                           n14306, C1 => n16352, C2 => n12024, ZN => n13583);
   U4805 : AOI221_X1 port map( B1 => registers_56_8_port, B2 => n16265, C1 => 
                           registers_60_8_port, C2 => n16262, A => n13599, ZN 
                           => n13598);
   U4806 : OAI222_X1 port map( A1 => n16259, A2 => n14576, B1 => n16256, B2 => 
                           n12058, C1 => n16253, C2 => n15248, ZN => n13599);
   U4807 : AOI221_X1 port map( B1 => registers_2_9_port, B2 => n16364, C1 => 
                           registers_29_9_port, C2 => n16361, A => n13541, ZN 
                           => n13540);
   U4808 : OAI222_X1 port map( A1 => n16358, A2 => n15011, B1 => n16355, B2 => 
                           n14307, C1 => n16352, C2 => n12025, ZN => n13541);
   U4809 : AOI221_X1 port map( B1 => registers_56_9_port, B2 => n16265, C1 => 
                           registers_60_9_port, C2 => n16262, A => n13557, ZN 
                           => n13556);
   U4810 : OAI222_X1 port map( A1 => n16259, A2 => n14577, B1 => n16256, B2 => 
                           n12059, C1 => n16253, C2 => n15249, ZN => n13557);
   U4811 : AOI221_X1 port map( B1 => registers_2_10_port, B2 => n16364, C1 => 
                           registers_29_10_port, C2 => n16361, A => n13499, ZN 
                           => n13498);
   U4812 : OAI222_X1 port map( A1 => n16358, A2 => n15012, B1 => n16355, B2 => 
                           n14308, C1 => n16352, C2 => n12026, ZN => n13499);
   U4813 : AOI221_X1 port map( B1 => registers_56_10_port, B2 => n16265, C1 => 
                           registers_60_10_port, C2 => n16262, A => n13515, ZN 
                           => n13514);
   U4814 : OAI222_X1 port map( A1 => n16259, A2 => n14578, B1 => n16256, B2 => 
                           n12060, C1 => n16253, C2 => n15250, ZN => n13515);
   U4815 : AOI221_X1 port map( B1 => registers_2_11_port, B2 => n16364, C1 => 
                           registers_29_11_port, C2 => n16361, A => n13457, ZN 
                           => n13456);
   U4816 : OAI222_X1 port map( A1 => n16358, A2 => n15013, B1 => n16355, B2 => 
                           n14309, C1 => n16352, C2 => n12027, ZN => n13457);
   U4817 : AOI221_X1 port map( B1 => registers_56_11_port, B2 => n16265, C1 => 
                           registers_60_11_port, C2 => n16262, A => n13473, ZN 
                           => n13472);
   U4818 : OAI222_X1 port map( A1 => n16259, A2 => n14579, B1 => n16256, B2 => 
                           n12098, C1 => n16253, C2 => n15251, ZN => n13473);
   U4819 : AOI221_X1 port map( B1 => registers_2_12_port, B2 => n16365, C1 => 
                           registers_29_12_port, C2 => n16362, A => n13415, ZN 
                           => n13414);
   U4820 : OAI222_X1 port map( A1 => n16359, A2 => n15014, B1 => n16356, B2 => 
                           n14310, C1 => n16353, C2 => n12028, ZN => n13415);
   U4821 : AOI221_X1 port map( B1 => registers_56_12_port, B2 => n16266, C1 => 
                           registers_60_12_port, C2 => n16263, A => n13431, ZN 
                           => n13430);
   U4822 : OAI222_X1 port map( A1 => n16260, A2 => n14580, B1 => n16257, B2 => 
                           n12099, C1 => n16254, C2 => n15252, ZN => n13431);
   U4823 : AOI221_X1 port map( B1 => registers_2_13_port, B2 => n16365, C1 => 
                           registers_29_13_port, C2 => n16362, A => n13373, ZN 
                           => n13372);
   U4824 : OAI222_X1 port map( A1 => n16359, A2 => n15015, B1 => n16356, B2 => 
                           n14311, C1 => n16353, C2 => n12030, ZN => n13373);
   U4825 : AOI221_X1 port map( B1 => registers_56_13_port, B2 => n16266, C1 => 
                           registers_60_13_port, C2 => n16263, A => n13389, ZN 
                           => n13388);
   U4826 : OAI222_X1 port map( A1 => n16260, A2 => n14581, B1 => n16257, B2 => 
                           n12100, C1 => n16254, C2 => n15253, ZN => n13389);
   U4827 : AOI221_X1 port map( B1 => registers_2_14_port, B2 => n16365, C1 => 
                           registers_29_14_port, C2 => n16362, A => n13331, ZN 
                           => n13330);
   U4828 : OAI222_X1 port map( A1 => n16359, A2 => n15016, B1 => n16356, B2 => 
                           n14312, C1 => n16353, C2 => n12031, ZN => n13331);
   U4829 : AOI221_X1 port map( B1 => registers_56_14_port, B2 => n16266, C1 => 
                           registers_60_14_port, C2 => n16263, A => n13347, ZN 
                           => n13346);
   U4830 : OAI222_X1 port map( A1 => n16260, A2 => n14582, B1 => n16257, B2 => 
                           n12101, C1 => n16254, C2 => n15254, ZN => n13347);
   U4831 : AOI221_X1 port map( B1 => registers_2_15_port, B2 => n16365, C1 => 
                           registers_29_15_port, C2 => n16362, A => n13289, ZN 
                           => n13288);
   U4832 : OAI222_X1 port map( A1 => n16359, A2 => n15017, B1 => n16356, B2 => 
                           n14313, C1 => n16353, C2 => n12032, ZN => n13289);
   U4833 : AOI221_X1 port map( B1 => registers_56_15_port, B2 => n16266, C1 => 
                           registers_60_15_port, C2 => n16263, A => n13305, ZN 
                           => n13304);
   U4834 : OAI222_X1 port map( A1 => n16260, A2 => n14583, B1 => n16257, B2 => 
                           n12102, C1 => n16254, C2 => n15255, ZN => n13305);
   U4835 : AOI221_X1 port map( B1 => registers_2_16_port, B2 => n16365, C1 => 
                           registers_29_16_port, C2 => n16362, A => n13247, ZN 
                           => n13246);
   U4836 : OAI222_X1 port map( A1 => n16359, A2 => n15018, B1 => n16356, B2 => 
                           n14314, C1 => n16353, C2 => n12033, ZN => n13247);
   U4837 : AOI221_X1 port map( B1 => registers_56_16_port, B2 => n16266, C1 => 
                           registers_60_16_port, C2 => n16263, A => n13263, ZN 
                           => n13262);
   U4838 : OAI222_X1 port map( A1 => n16260, A2 => n14584, B1 => n16257, B2 => 
                           n12103, C1 => n16254, C2 => n15256, ZN => n13263);
   U4839 : AOI221_X1 port map( B1 => registers_2_17_port, B2 => n16365, C1 => 
                           registers_29_17_port, C2 => n16362, A => n13205, ZN 
                           => n13204);
   U4840 : OAI222_X1 port map( A1 => n16359, A2 => n15019, B1 => n16356, B2 => 
                           n14315, C1 => n16353, C2 => n12034, ZN => n13205);
   U4841 : AOI221_X1 port map( B1 => registers_56_17_port, B2 => n16266, C1 => 
                           registers_60_17_port, C2 => n16263, A => n13221, ZN 
                           => n13220);
   U4842 : OAI222_X1 port map( A1 => n16260, A2 => n14585, B1 => n16257, B2 => 
                           n12104, C1 => n16254, C2 => n15257, ZN => n13221);
   U4843 : AOI221_X1 port map( B1 => registers_2_18_port, B2 => n16365, C1 => 
                           registers_29_18_port, C2 => n16362, A => n13163, ZN 
                           => n13162);
   U4844 : OAI222_X1 port map( A1 => n16359, A2 => n15020, B1 => n16356, B2 => 
                           n14316, C1 => n16353, C2 => n12035, ZN => n13163);
   U4845 : AOI221_X1 port map( B1 => registers_56_18_port, B2 => n16266, C1 => 
                           registers_60_18_port, C2 => n16263, A => n13179, ZN 
                           => n13178);
   U4846 : OAI222_X1 port map( A1 => n16260, A2 => n14586, B1 => n16257, B2 => 
                           n12105, C1 => n16254, C2 => n15258, ZN => n13179);
   U4847 : AOI221_X1 port map( B1 => registers_2_19_port, B2 => n16365, C1 => 
                           registers_29_19_port, C2 => n16362, A => n13121, ZN 
                           => n13120);
   U4848 : OAI222_X1 port map( A1 => n16359, A2 => n15021, B1 => n16356, B2 => 
                           n14317, C1 => n16353, C2 => n12036, ZN => n13121);
   U4849 : AOI221_X1 port map( B1 => registers_56_19_port, B2 => n16266, C1 => 
                           registers_60_19_port, C2 => n16263, A => n13137, ZN 
                           => n13136);
   U4850 : OAI222_X1 port map( A1 => n16260, A2 => n14587, B1 => n16257, B2 => 
                           n12148, C1 => n16254, C2 => n15259, ZN => n13137);
   U4851 : AOI221_X1 port map( B1 => registers_2_20_port, B2 => n16365, C1 => 
                           registers_29_20_port, C2 => n16362, A => n13079, ZN 
                           => n13078);
   U4852 : OAI222_X1 port map( A1 => n16359, A2 => n15022, B1 => n16356, B2 => 
                           n14318, C1 => n16353, C2 => n12037, ZN => n13079);
   U4853 : AOI221_X1 port map( B1 => registers_56_20_port, B2 => n16266, C1 => 
                           registers_60_20_port, C2 => n16263, A => n13095, ZN 
                           => n13094);
   U4854 : OAI222_X1 port map( A1 => n16260, A2 => n14588, B1 => n16257, B2 => 
                           n12150, C1 => n16254, C2 => n15260, ZN => n13095);
   U4855 : AOI221_X1 port map( B1 => registers_2_21_port, B2 => n16365, C1 => 
                           registers_29_21_port, C2 => n16362, A => n13037, ZN 
                           => n13036);
   U4856 : OAI222_X1 port map( A1 => n16359, A2 => n15023, B1 => n16356, B2 => 
                           n14319, C1 => n16353, C2 => n12038, ZN => n13037);
   U4857 : AOI221_X1 port map( B1 => registers_56_21_port, B2 => n16266, C1 => 
                           registers_60_21_port, C2 => n16263, A => n13053, ZN 
                           => n13052);
   U4858 : OAI222_X1 port map( A1 => n16260, A2 => n14589, B1 => n16257, B2 => 
                           n12151, C1 => n16254, C2 => n15261, ZN => n13053);
   U4859 : AOI221_X1 port map( B1 => registers_2_22_port, B2 => n16365, C1 => 
                           registers_29_22_port, C2 => n16362, A => n12995, ZN 
                           => n12994);
   U4860 : OAI222_X1 port map( A1 => n16359, A2 => n15024, B1 => n16356, B2 => 
                           n14320, C1 => n16353, C2 => n12039, ZN => n12995);
   U4861 : AOI221_X1 port map( B1 => registers_56_22_port, B2 => n16266, C1 => 
                           registers_60_22_port, C2 => n16263, A => n13011, ZN 
                           => n13010);
   U4862 : OAI222_X1 port map( A1 => n16260, A2 => n14590, B1 => n16257, B2 => 
                           n12152, C1 => n16254, C2 => n15262, ZN => n13011);
   U4863 : AOI221_X1 port map( B1 => registers_2_23_port, B2 => n16365, C1 => 
                           registers_29_23_port, C2 => n16362, A => n12953, ZN 
                           => n12952);
   U4864 : OAI222_X1 port map( A1 => n16359, A2 => n15025, B1 => n16356, B2 => 
                           n14321, C1 => n16353, C2 => n12040, ZN => n12953);
   U4865 : AOI221_X1 port map( B1 => registers_56_23_port, B2 => n16266, C1 => 
                           registers_60_23_port, C2 => n16263, A => n12969, ZN 
                           => n12968);
   U4866 : OAI222_X1 port map( A1 => n16260, A2 => n14591, B1 => n16257, B2 => 
                           n12153, C1 => n16254, C2 => n15263, ZN => n12969);
   U4867 : AOI221_X1 port map( B1 => registers_2_24_port, B2 => n16366, C1 => 
                           registers_29_24_port, C2 => n16363, A => n12911, ZN 
                           => n12910);
   U4868 : OAI222_X1 port map( A1 => n16360, A2 => n15026, B1 => n16357, B2 => 
                           n14322, C1 => n16354, C2 => n12041, ZN => n12911);
   U4869 : AOI221_X1 port map( B1 => registers_12_24_port, B2 => n16411, C1 => 
                           registers_17_24_port, C2 => n16408, A => n12903, ZN 
                           => n12902);
   U4870 : OAI22_X1 port map( A1 => n16405, A2 => n15065, B1 => n16402, B2 => 
                           n14419, ZN => n12903);
   U4871 : AOI221_X1 port map( B1 => registers_56_24_port, B2 => n16267, C1 => 
                           registers_60_24_port, C2 => n16264, A => n12927, ZN 
                           => n12926);
   U4872 : OAI222_X1 port map( A1 => n16261, A2 => n14592, B1 => n16258, B2 => 
                           n12154, C1 => n16255, C2 => n15264, ZN => n12927);
   U4873 : AOI221_X1 port map( B1 => registers_2_25_port, B2 => n16366, C1 => 
                           registers_29_25_port, C2 => n16363, A => n12869, ZN 
                           => n12868);
   U4874 : OAI222_X1 port map( A1 => n16360, A2 => n15027, B1 => n16357, B2 => 
                           n14323, C1 => n16354, C2 => n12042, ZN => n12869);
   U4875 : AOI221_X1 port map( B1 => registers_12_25_port, B2 => n16411, C1 => 
                           registers_17_25_port, C2 => n16408, A => n12861, ZN 
                           => n12860);
   U4876 : OAI22_X1 port map( A1 => n16405, A2 => n15066, B1 => n16402, B2 => 
                           n14420, ZN => n12861);
   U4877 : AOI221_X1 port map( B1 => registers_56_25_port, B2 => n16267, C1 => 
                           registers_60_25_port, C2 => n16264, A => n12885, ZN 
                           => n12884);
   U4878 : OAI222_X1 port map( A1 => n16261, A2 => n14593, B1 => n16258, B2 => 
                           n12155, C1 => n16255, C2 => n15265, ZN => n12885);
   U4879 : AOI221_X1 port map( B1 => registers_2_26_port, B2 => n16366, C1 => 
                           registers_29_26_port, C2 => n16363, A => n12827, ZN 
                           => n12826);
   U4880 : OAI222_X1 port map( A1 => n16360, A2 => n15028, B1 => n16357, B2 => 
                           n14324, C1 => n16354, C2 => n12043, ZN => n12827);
   U4881 : AOI221_X1 port map( B1 => registers_12_26_port, B2 => n16411, C1 => 
                           registers_17_26_port, C2 => n16408, A => n12819, ZN 
                           => n12818);
   U4882 : OAI22_X1 port map( A1 => n16405, A2 => n15067, B1 => n16402, B2 => 
                           n14421, ZN => n12819);
   U4883 : AOI221_X1 port map( B1 => registers_56_26_port, B2 => n16267, C1 => 
                           registers_60_26_port, C2 => n16264, A => n12843, ZN 
                           => n12842);
   U4884 : OAI222_X1 port map( A1 => n16261, A2 => n14594, B1 => n16258, B2 => 
                           n12156, C1 => n16255, C2 => n15266, ZN => n12843);
   U4885 : AOI221_X1 port map( B1 => registers_2_27_port, B2 => n16366, C1 => 
                           registers_29_27_port, C2 => n16363, A => n12785, ZN 
                           => n12784);
   U4886 : OAI222_X1 port map( A1 => n16360, A2 => n15029, B1 => n16357, B2 => 
                           n14325, C1 => n16354, C2 => n12044, ZN => n12785);
   U4887 : AOI221_X1 port map( B1 => registers_12_27_port, B2 => n16411, C1 => 
                           registers_17_27_port, C2 => n16408, A => n12777, ZN 
                           => n12776);
   U4888 : OAI22_X1 port map( A1 => n16405, A2 => n15068, B1 => n16402, B2 => 
                           n14422, ZN => n12777);
   U4889 : AOI221_X1 port map( B1 => registers_56_27_port, B2 => n16267, C1 => 
                           registers_60_27_port, C2 => n16264, A => n12801, ZN 
                           => n12800);
   U4890 : OAI222_X1 port map( A1 => n16261, A2 => n14595, B1 => n16258, B2 => 
                           n12157, C1 => n16255, C2 => n15267, ZN => n12801);
   U4891 : AOI221_X1 port map( B1 => registers_2_28_port, B2 => n16366, C1 => 
                           registers_29_28_port, C2 => n16363, A => n12743, ZN 
                           => n12742);
   U4892 : OAI222_X1 port map( A1 => n16360, A2 => n15030, B1 => n16357, B2 => 
                           n14326, C1 => n16354, C2 => n12045, ZN => n12743);
   U4893 : AOI221_X1 port map( B1 => registers_12_28_port, B2 => n16411, C1 => 
                           registers_17_28_port, C2 => n16408, A => n12735, ZN 
                           => n12734);
   U4894 : OAI22_X1 port map( A1 => n16405, A2 => n15069, B1 => n16402, B2 => 
                           n14423, ZN => n12735);
   U4895 : AOI221_X1 port map( B1 => registers_56_28_port, B2 => n16267, C1 => 
                           registers_60_28_port, C2 => n16264, A => n12759, ZN 
                           => n12758);
   U4896 : OAI222_X1 port map( A1 => n16261, A2 => n14596, B1 => n16258, B2 => 
                           n12158, C1 => n16255, C2 => n15268, ZN => n12759);
   U4897 : AOI221_X1 port map( B1 => registers_2_29_port, B2 => n16366, C1 => 
                           registers_29_29_port, C2 => n16363, A => n12701, ZN 
                           => n12700);
   U4898 : OAI222_X1 port map( A1 => n16360, A2 => n15031, B1 => n16357, B2 => 
                           n14327, C1 => n16354, C2 => n12046, ZN => n12701);
   U4899 : AOI221_X1 port map( B1 => registers_12_29_port, B2 => n16411, C1 => 
                           registers_17_29_port, C2 => n16408, A => n12693, ZN 
                           => n12692);
   U4900 : OAI22_X1 port map( A1 => n16405, A2 => n15070, B1 => n16402, B2 => 
                           n14424, ZN => n12693);
   U4901 : AOI221_X1 port map( B1 => registers_56_29_port, B2 => n16267, C1 => 
                           registers_60_29_port, C2 => n16264, A => n12717, ZN 
                           => n12716);
   U4902 : OAI222_X1 port map( A1 => n16261, A2 => n14597, B1 => n16258, B2 => 
                           n12159, C1 => n16255, C2 => n15269, ZN => n12717);
   U4903 : AOI221_X1 port map( B1 => registers_2_30_port, B2 => n16366, C1 => 
                           registers_29_30_port, C2 => n16363, A => n12658, ZN 
                           => n12657);
   U4904 : OAI222_X1 port map( A1 => n16360, A2 => n14857, B1 => n16357, B2 => 
                           n14054, C1 => n16354, C2 => n11904, ZN => n12658);
   U4905 : AOI221_X1 port map( B1 => registers_12_30_port, B2 => n16411, C1 => 
                           registers_17_30_port, C2 => n16408, A => n12649, ZN 
                           => n12648);
   U4906 : OAI22_X1 port map( A1 => n16405, A2 => n14870, B1 => n16402, B2 => 
                           n14060, ZN => n12649);
   U4907 : AOI221_X1 port map( B1 => registers_56_30_port, B2 => n16267, C1 => 
                           registers_60_30_port, C2 => n16264, A => n12675, ZN 
                           => n12674);
   U4908 : OAI222_X1 port map( A1 => n16261, A2 => n14534, B1 => n16258, B2 => 
                           n12048, C1 => n16255, C2 => n15033, ZN => n12675);
   U4909 : AOI221_X1 port map( B1 => registers_2_31_port, B2 => n16366, C1 => 
                           registers_29_31_port, C2 => n16363, A => n12563, ZN 
                           => n12560);
   U4910 : OAI222_X1 port map( A1 => n16360, A2 => n15032, B1 => n16357, B2 => 
                           n14328, C1 => n16354, C2 => n12047, ZN => n12563);
   U4911 : AOI221_X1 port map( B1 => registers_12_31_port, B2 => n16411, C1 => 
                           registers_17_31_port, C2 => n16408, A => n12539, ZN 
                           => n12536);
   U4912 : OAI22_X1 port map( A1 => n16405, A2 => n15071, B1 => n16402, B2 => 
                           n14425, ZN => n12539);
   U4913 : AOI221_X1 port map( B1 => registers_56_31_port, B2 => n16267, C1 => 
                           registers_60_31_port, C2 => n16264, A => n12614, ZN 
                           => n12611);
   U4914 : OAI222_X1 port map( A1 => n16261, A2 => n14535, B1 => n16258, B2 => 
                           n12049, C1 => n16255, C2 => n15034, ZN => n12614);
   U4915 : AOI221_X1 port map( B1 => registers_2_0_port, B2 => n16616, C1 => 
                           registers_29_0_port, C2 => n16613, A => n12461, ZN 
                           => n12460);
   U4916 : OAI222_X1 port map( A1 => n16610, A2 => n15004, B1 => n16607, B2 => 
                           n14300, C1 => n16604, C2 => n12018, ZN => n12461);
   U4917 : AOI221_X1 port map( B1 => registers_56_0_port, B2 => n16517, C1 => 
                           registers_60_0_port, C2 => n16514, A => n12487, ZN 
                           => n12486);
   U4918 : OAI222_X1 port map( A1 => n16511, A2 => n14573, B1 => n16508, B2 => 
                           n12055, C1 => n16505, C2 => n15245, ZN => n12487);
   U4919 : AOI221_X1 port map( B1 => registers_2_1_port, B2 => n16616, C1 => 
                           registers_29_1_port, C2 => n16613, A => n12281, ZN 
                           => n12280);
   U4920 : OAI222_X1 port map( A1 => n16610, A2 => n15005, B1 => n16607, B2 => 
                           n14301, C1 => n16604, C2 => n12019, ZN => n12281);
   U4921 : AOI221_X1 port map( B1 => registers_2_2_port, B2 => n16616, C1 => 
                           registers_29_2_port, C2 => n16613, A => n12128, ZN 
                           => n12127);
   U4922 : OAI222_X1 port map( A1 => n16610, A2 => n15006, B1 => n16607, B2 => 
                           n14302, C1 => n16604, C2 => n12020, ZN => n12128);
   U4923 : AOI221_X1 port map( B1 => registers_2_3_port, B2 => n16616, C1 => 
                           registers_29_3_port, C2 => n16613, A => n11975, ZN 
                           => n11974);
   U4924 : OAI222_X1 port map( A1 => n16610, A2 => n14989, B1 => n16607, B2 => 
                           n14282, C1 => n16604, C2 => n12016, ZN => n11975);
   U4925 : AOI221_X1 port map( B1 => registers_2_4_port, B2 => n16616, C1 => 
                           registers_29_4_port, C2 => n16613, A => n11822, ZN 
                           => n11821);
   U4926 : OAI222_X1 port map( A1 => n16610, A2 => n14990, B1 => n16607, B2 => 
                           n14283, C1 => n16604, C2 => n12017, ZN => n11822);
   U4927 : AOI221_X1 port map( B1 => registers_56_4_port, B2 => n16517, C1 => 
                           registers_60_4_port, C2 => n16514, A => n11838, ZN 
                           => n11837);
   U4928 : OAI222_X1 port map( A1 => n16511, A2 => n14538, B1 => n16508, B2 => 
                           n12050, C1 => n16505, C2 => n15241, ZN => n11838);
   U4929 : AOI221_X1 port map( B1 => registers_2_5_port, B2 => n16616, C1 => 
                           registers_29_5_port, C2 => n16613, A => n11779, ZN 
                           => n11778);
   U4930 : OAI222_X1 port map( A1 => n16610, A2 => n15007, B1 => n16607, B2 => 
                           n14303, C1 => n16604, C2 => n12021, ZN => n11779);
   U4931 : AOI221_X1 port map( B1 => registers_56_5_port, B2 => n16517, C1 => 
                           registers_60_5_port, C2 => n16514, A => n11795, ZN 
                           => n11794);
   U4932 : OAI222_X1 port map( A1 => n16511, A2 => n14539, B1 => n16508, B2 => 
                           n12051, C1 => n16505, C2 => n15242, ZN => n11795);
   U4933 : AOI221_X1 port map( B1 => registers_2_6_port, B2 => n16616, C1 => 
                           registers_29_6_port, C2 => n16613, A => n11736, ZN 
                           => n11735);
   U4934 : OAI222_X1 port map( A1 => n16610, A2 => n15008, B1 => n16607, B2 => 
                           n14304, C1 => n16604, C2 => n12022, ZN => n11736);
   U4935 : AOI221_X1 port map( B1 => registers_56_6_port, B2 => n16517, C1 => 
                           registers_60_6_port, C2 => n16514, A => n11752, ZN 
                           => n11751);
   U4936 : OAI222_X1 port map( A1 => n16511, A2 => n14574, B1 => n16508, B2 => 
                           n12056, C1 => n16505, C2 => n15246, ZN => n11752);
   U4937 : AOI221_X1 port map( B1 => registers_2_7_port, B2 => n16616, C1 => 
                           registers_29_7_port, C2 => n16613, A => n11693, ZN 
                           => n11692);
   U4938 : OAI222_X1 port map( A1 => n16610, A2 => n15009, B1 => n16607, B2 => 
                           n14305, C1 => n16604, C2 => n12023, ZN => n11693);
   U4939 : AOI221_X1 port map( B1 => registers_56_7_port, B2 => n16517, C1 => 
                           registers_60_7_port, C2 => n16514, A => n11709, ZN 
                           => n11708);
   U4940 : OAI222_X1 port map( A1 => n16511, A2 => n14575, B1 => n16508, B2 => 
                           n12057, C1 => n16505, C2 => n15247, ZN => n11709);
   U4941 : AOI221_X1 port map( B1 => registers_2_8_port, B2 => n16616, C1 => 
                           registers_29_8_port, C2 => n16613, A => n11650, ZN 
                           => n11649);
   U4942 : OAI222_X1 port map( A1 => n16610, A2 => n15010, B1 => n16607, B2 => 
                           n14306, C1 => n16604, C2 => n12024, ZN => n11650);
   U4943 : AOI221_X1 port map( B1 => registers_56_8_port, B2 => n16517, C1 => 
                           registers_60_8_port, C2 => n16514, A => n11666, ZN 
                           => n11665);
   U4944 : OAI222_X1 port map( A1 => n16511, A2 => n14576, B1 => n16508, B2 => 
                           n12058, C1 => n16505, C2 => n15248, ZN => n11666);
   U4945 : AOI221_X1 port map( B1 => registers_2_9_port, B2 => n16616, C1 => 
                           registers_29_9_port, C2 => n16613, A => n11607, ZN 
                           => n11606);
   U4946 : OAI222_X1 port map( A1 => n16610, A2 => n15011, B1 => n16607, B2 => 
                           n14307, C1 => n16604, C2 => n12025, ZN => n11607);
   U4947 : AOI221_X1 port map( B1 => registers_56_9_port, B2 => n16517, C1 => 
                           registers_60_9_port, C2 => n16514, A => n11623, ZN 
                           => n11622);
   U4948 : OAI222_X1 port map( A1 => n16511, A2 => n14577, B1 => n16508, B2 => 
                           n12059, C1 => n16505, C2 => n15249, ZN => n11623);
   U4949 : AOI221_X1 port map( B1 => registers_2_10_port, B2 => n16616, C1 => 
                           registers_29_10_port, C2 => n16613, A => n11564, ZN 
                           => n11563);
   U4950 : OAI222_X1 port map( A1 => n16610, A2 => n15012, B1 => n16607, B2 => 
                           n14308, C1 => n16604, C2 => n12026, ZN => n11564);
   U4951 : AOI221_X1 port map( B1 => registers_56_10_port, B2 => n16517, C1 => 
                           registers_60_10_port, C2 => n16514, A => n11580, ZN 
                           => n11579);
   U4952 : OAI222_X1 port map( A1 => n16511, A2 => n14578, B1 => n16508, B2 => 
                           n12060, C1 => n16505, C2 => n15250, ZN => n11580);
   U4953 : AOI221_X1 port map( B1 => registers_2_11_port, B2 => n16616, C1 => 
                           registers_29_11_port, C2 => n16613, A => n11521, ZN 
                           => n11520);
   U4954 : OAI222_X1 port map( A1 => n16610, A2 => n15013, B1 => n16607, B2 => 
                           n14309, C1 => n16604, C2 => n12027, ZN => n11521);
   U4955 : AOI221_X1 port map( B1 => registers_56_11_port, B2 => n16517, C1 => 
                           registers_60_11_port, C2 => n16514, A => n11537, ZN 
                           => n11536);
   U4956 : OAI222_X1 port map( A1 => n16511, A2 => n14579, B1 => n16508, B2 => 
                           n12098, C1 => n16505, C2 => n15251, ZN => n11537);
   U4957 : AOI221_X1 port map( B1 => registers_2_12_port, B2 => n16617, C1 => 
                           registers_29_12_port, C2 => n16614, A => n11478, ZN 
                           => n11477);
   U4958 : OAI222_X1 port map( A1 => n16611, A2 => n15014, B1 => n16608, B2 => 
                           n14310, C1 => n16605, C2 => n12028, ZN => n11478);
   U4959 : AOI221_X1 port map( B1 => registers_56_12_port, B2 => n16518, C1 => 
                           registers_60_12_port, C2 => n16515, A => n11494, ZN 
                           => n11493);
   U4960 : OAI222_X1 port map( A1 => n16512, A2 => n14580, B1 => n16509, B2 => 
                           n12099, C1 => n16506, C2 => n15252, ZN => n11494);
   U4961 : AOI221_X1 port map( B1 => registers_2_13_port, B2 => n16617, C1 => 
                           registers_29_13_port, C2 => n16614, A => n11434, ZN 
                           => n11433);
   U4962 : OAI222_X1 port map( A1 => n16611, A2 => n15015, B1 => n16608, B2 => 
                           n14311, C1 => n16605, C2 => n12030, ZN => n11434);
   U4963 : AOI221_X1 port map( B1 => registers_56_13_port, B2 => n16518, C1 => 
                           registers_60_13_port, C2 => n16515, A => n11450, ZN 
                           => n11449);
   U4964 : OAI222_X1 port map( A1 => n16512, A2 => n14581, B1 => n16509, B2 => 
                           n12100, C1 => n16506, C2 => n15253, ZN => n11450);
   U4965 : AOI221_X1 port map( B1 => registers_2_14_port, B2 => n16617, C1 => 
                           registers_29_14_port, C2 => n16614, A => n11391, ZN 
                           => n11390);
   U4966 : OAI222_X1 port map( A1 => n16611, A2 => n15016, B1 => n16608, B2 => 
                           n14312, C1 => n16605, C2 => n12031, ZN => n11391);
   U4967 : AOI221_X1 port map( B1 => registers_56_14_port, B2 => n16518, C1 => 
                           registers_60_14_port, C2 => n16515, A => n11407, ZN 
                           => n11406);
   U4968 : OAI222_X1 port map( A1 => n16512, A2 => n14582, B1 => n16509, B2 => 
                           n12101, C1 => n16506, C2 => n15254, ZN => n11407);
   U4969 : AOI221_X1 port map( B1 => registers_2_15_port, B2 => n16617, C1 => 
                           registers_29_15_port, C2 => n16614, A => n11348, ZN 
                           => n11347);
   U4970 : OAI222_X1 port map( A1 => n16611, A2 => n15017, B1 => n16608, B2 => 
                           n14313, C1 => n16605, C2 => n12032, ZN => n11348);
   U4971 : AOI221_X1 port map( B1 => registers_56_15_port, B2 => n16518, C1 => 
                           registers_60_15_port, C2 => n16515, A => n11364, ZN 
                           => n11363);
   U4972 : OAI222_X1 port map( A1 => n16512, A2 => n14583, B1 => n16509, B2 => 
                           n12102, C1 => n16506, C2 => n15255, ZN => n11364);
   U4973 : AOI221_X1 port map( B1 => registers_2_16_port, B2 => n16617, C1 => 
                           registers_29_16_port, C2 => n16614, A => n11305, ZN 
                           => n11304);
   U4974 : OAI222_X1 port map( A1 => n16611, A2 => n15018, B1 => n16608, B2 => 
                           n14314, C1 => n16605, C2 => n12033, ZN => n11305);
   U4975 : AOI221_X1 port map( B1 => registers_56_16_port, B2 => n16518, C1 => 
                           registers_60_16_port, C2 => n16515, A => n11321, ZN 
                           => n11320);
   U4976 : OAI222_X1 port map( A1 => n16512, A2 => n14584, B1 => n16509, B2 => 
                           n12103, C1 => n16506, C2 => n15256, ZN => n11321);
   U4977 : AOI221_X1 port map( B1 => registers_2_17_port, B2 => n16617, C1 => 
                           registers_29_17_port, C2 => n16614, A => n11262, ZN 
                           => n11261);
   U4978 : OAI222_X1 port map( A1 => n16611, A2 => n15019, B1 => n16608, B2 => 
                           n14315, C1 => n16605, C2 => n12034, ZN => n11262);
   U4979 : AOI221_X1 port map( B1 => registers_56_17_port, B2 => n16518, C1 => 
                           registers_60_17_port, C2 => n16515, A => n11278, ZN 
                           => n11277);
   U4980 : OAI222_X1 port map( A1 => n16512, A2 => n14585, B1 => n16509, B2 => 
                           n12104, C1 => n16506, C2 => n15257, ZN => n11278);
   U4981 : AOI221_X1 port map( B1 => registers_2_18_port, B2 => n16617, C1 => 
                           registers_29_18_port, C2 => n16614, A => n11219, ZN 
                           => n11218);
   U4982 : OAI222_X1 port map( A1 => n16611, A2 => n15020, B1 => n16608, B2 => 
                           n14316, C1 => n16605, C2 => n12035, ZN => n11219);
   U4983 : AOI221_X1 port map( B1 => registers_56_18_port, B2 => n16518, C1 => 
                           registers_60_18_port, C2 => n16515, A => n11235, ZN 
                           => n11234);
   U4984 : OAI222_X1 port map( A1 => n16512, A2 => n14586, B1 => n16509, B2 => 
                           n12105, C1 => n16506, C2 => n15258, ZN => n11235);
   U4985 : AOI221_X1 port map( B1 => registers_2_19_port, B2 => n16617, C1 => 
                           registers_29_19_port, C2 => n16614, A => n11176, ZN 
                           => n11175);
   U4986 : OAI222_X1 port map( A1 => n16611, A2 => n15021, B1 => n16608, B2 => 
                           n14317, C1 => n16605, C2 => n12036, ZN => n11176);
   U4987 : AOI221_X1 port map( B1 => registers_56_19_port, B2 => n16518, C1 => 
                           registers_60_19_port, C2 => n16515, A => n11192, ZN 
                           => n11191);
   U4988 : OAI222_X1 port map( A1 => n16512, A2 => n14587, B1 => n16509, B2 => 
                           n12148, C1 => n16506, C2 => n15259, ZN => n11192);
   U4989 : AOI221_X1 port map( B1 => registers_2_20_port, B2 => n16617, C1 => 
                           registers_29_20_port, C2 => n16614, A => n11133, ZN 
                           => n11132);
   U4990 : OAI222_X1 port map( A1 => n16611, A2 => n15022, B1 => n16608, B2 => 
                           n14318, C1 => n16605, C2 => n12037, ZN => n11133);
   U4991 : AOI221_X1 port map( B1 => registers_56_20_port, B2 => n16518, C1 => 
                           registers_60_20_port, C2 => n16515, A => n11149, ZN 
                           => n11148);
   U4992 : OAI222_X1 port map( A1 => n16512, A2 => n14588, B1 => n16509, B2 => 
                           n12150, C1 => n16506, C2 => n15260, ZN => n11149);
   U4993 : AOI221_X1 port map( B1 => registers_2_21_port, B2 => n16617, C1 => 
                           registers_29_21_port, C2 => n16614, A => n11090, ZN 
                           => n11089);
   U4994 : OAI222_X1 port map( A1 => n16611, A2 => n15023, B1 => n16608, B2 => 
                           n14319, C1 => n16605, C2 => n12038, ZN => n11090);
   U4995 : AOI221_X1 port map( B1 => registers_56_21_port, B2 => n16518, C1 => 
                           registers_60_21_port, C2 => n16515, A => n11106, ZN 
                           => n11105);
   U4996 : OAI222_X1 port map( A1 => n16512, A2 => n14589, B1 => n16509, B2 => 
                           n12151, C1 => n16506, C2 => n15261, ZN => n11106);
   U4997 : AOI221_X1 port map( B1 => registers_2_22_port, B2 => n16617, C1 => 
                           registers_29_22_port, C2 => n16614, A => n11047, ZN 
                           => n11046);
   U4998 : OAI222_X1 port map( A1 => n16611, A2 => n15024, B1 => n16608, B2 => 
                           n14320, C1 => n16605, C2 => n12039, ZN => n11047);
   U4999 : AOI221_X1 port map( B1 => registers_56_22_port, B2 => n16518, C1 => 
                           registers_60_22_port, C2 => n16515, A => n11063, ZN 
                           => n11062);
   U5000 : OAI222_X1 port map( A1 => n16512, A2 => n14590, B1 => n16509, B2 => 
                           n12152, C1 => n16506, C2 => n15262, ZN => n11063);
   U5001 : AOI221_X1 port map( B1 => registers_2_23_port, B2 => n16617, C1 => 
                           registers_29_23_port, C2 => n16614, A => n11004, ZN 
                           => n11003);
   U5002 : OAI222_X1 port map( A1 => n16611, A2 => n15025, B1 => n16608, B2 => 
                           n14321, C1 => n16605, C2 => n12040, ZN => n11004);
   U5003 : AOI221_X1 port map( B1 => registers_56_23_port, B2 => n16518, C1 => 
                           registers_60_23_port, C2 => n16515, A => n11020, ZN 
                           => n11019);
   U5004 : OAI222_X1 port map( A1 => n16512, A2 => n14591, B1 => n16509, B2 => 
                           n12153, C1 => n16506, C2 => n15263, ZN => n11020);
   U5005 : AOI221_X1 port map( B1 => registers_2_24_port, B2 => n16618, C1 => 
                           registers_29_24_port, C2 => n16615, A => n10961, ZN 
                           => n10960);
   U5006 : OAI222_X1 port map( A1 => n16612, A2 => n15026, B1 => n16609, B2 => 
                           n14322, C1 => n16606, C2 => n12041, ZN => n10961);
   U5007 : AOI221_X1 port map( B1 => registers_12_24_port, B2 => n16663, C1 => 
                           registers_15_24_port, C2 => n16660, A => n10953, ZN 
                           => n10952);
   U5008 : OAI22_X1 port map( A1 => n16657, A2 => n15065, B1 => n16654, B2 => 
                           n14419, ZN => n10953);
   U5009 : AOI221_X1 port map( B1 => net227344, B2 => n16567, C1 => 
                           registers_44_24_port, C2 => n16564, A => n10969, ZN 
                           => n10968);
   U5010 : OAI22_X1 port map( A1 => n16561, A2 => n15144, B1 => n16558, B2 => 
                           n14527, ZN => n10969);
   U5011 : AOI221_X1 port map( B1 => registers_56_24_port, B2 => n16519, C1 => 
                           registers_60_24_port, C2 => n16516, A => n10977, ZN 
                           => n10976);
   U5012 : OAI222_X1 port map( A1 => n16513, A2 => n14592, B1 => n16510, B2 => 
                           n12154, C1 => n16507, C2 => n15264, ZN => n10977);
   U5013 : AOI221_X1 port map( B1 => registers_2_25_port, B2 => n16618, C1 => 
                           registers_29_25_port, C2 => n16615, A => n10918, ZN 
                           => n10917);
   U5014 : OAI222_X1 port map( A1 => n16612, A2 => n15027, B1 => n16609, B2 => 
                           n14323, C1 => n16606, C2 => n12042, ZN => n10918);
   U5015 : AOI221_X1 port map( B1 => registers_12_25_port, B2 => n16663, C1 => 
                           registers_15_25_port, C2 => n16660, A => n10910, ZN 
                           => n10909);
   U5016 : OAI22_X1 port map( A1 => n16657, A2 => n15066, B1 => n16654, B2 => 
                           n14420, ZN => n10910);
   U5017 : AOI221_X1 port map( B1 => net227362, B2 => n16567, C1 => 
                           registers_44_25_port, C2 => n16564, A => n10926, ZN 
                           => n10925);
   U5018 : OAI22_X1 port map( A1 => n16561, A2 => n15145, B1 => n16558, B2 => 
                           n14528, ZN => n10926);
   U5019 : AOI221_X1 port map( B1 => registers_56_25_port, B2 => n16519, C1 => 
                           registers_60_25_port, C2 => n16516, A => n10934, ZN 
                           => n10933);
   U5020 : OAI222_X1 port map( A1 => n16513, A2 => n14593, B1 => n16510, B2 => 
                           n12155, C1 => n16507, C2 => n15265, ZN => n10934);
   U5021 : AOI221_X1 port map( B1 => registers_2_26_port, B2 => n16618, C1 => 
                           registers_29_26_port, C2 => n16615, A => n10875, ZN 
                           => n10874);
   U5022 : OAI222_X1 port map( A1 => n16612, A2 => n15028, B1 => n16609, B2 => 
                           n14324, C1 => n16606, C2 => n12043, ZN => n10875);
   U5023 : AOI221_X1 port map( B1 => registers_12_26_port, B2 => n16663, C1 => 
                           registers_15_26_port, C2 => n16660, A => n10867, ZN 
                           => n10866);
   U5024 : OAI22_X1 port map( A1 => n16657, A2 => n15067, B1 => n16654, B2 => 
                           n14421, ZN => n10867);
   U5025 : AOI221_X1 port map( B1 => net227380, B2 => n16567, C1 => 
                           registers_44_26_port, C2 => n16564, A => n10883, ZN 
                           => n10882);
   U5026 : OAI22_X1 port map( A1 => n16561, A2 => n15146, B1 => n16558, B2 => 
                           n14529, ZN => n10883);
   U5027 : AOI221_X1 port map( B1 => registers_56_26_port, B2 => n16519, C1 => 
                           registers_60_26_port, C2 => n16516, A => n10891, ZN 
                           => n10890);
   U5028 : OAI222_X1 port map( A1 => n16513, A2 => n14594, B1 => n16510, B2 => 
                           n12156, C1 => n16507, C2 => n15266, ZN => n10891);
   U5029 : AOI221_X1 port map( B1 => registers_2_27_port, B2 => n16618, C1 => 
                           registers_29_27_port, C2 => n16615, A => n10832, ZN 
                           => n10831);
   U5030 : OAI222_X1 port map( A1 => n16612, A2 => n15029, B1 => n16609, B2 => 
                           n14325, C1 => n16606, C2 => n12044, ZN => n10832);
   U5031 : AOI221_X1 port map( B1 => registers_12_27_port, B2 => n16663, C1 => 
                           registers_15_27_port, C2 => n16660, A => n10824, ZN 
                           => n10823);
   U5032 : OAI22_X1 port map( A1 => n16657, A2 => n15068, B1 => n16654, B2 => 
                           n14422, ZN => n10824);
   U5033 : AOI221_X1 port map( B1 => net227398, B2 => n16567, C1 => 
                           registers_44_27_port, C2 => n16564, A => n10840, ZN 
                           => n10839);
   U5034 : OAI22_X1 port map( A1 => n16561, A2 => n15147, B1 => n16558, B2 => 
                           n14530, ZN => n10840);
   U5035 : AOI221_X1 port map( B1 => registers_56_27_port, B2 => n16519, C1 => 
                           registers_60_27_port, C2 => n16516, A => n10848, ZN 
                           => n10847);
   U5036 : OAI222_X1 port map( A1 => n16513, A2 => n14595, B1 => n16510, B2 => 
                           n12157, C1 => n16507, C2 => n15267, ZN => n10848);
   U5037 : AOI221_X1 port map( B1 => registers_2_28_port, B2 => n16618, C1 => 
                           registers_29_28_port, C2 => n16615, A => n10789, ZN 
                           => n10788);
   U5038 : OAI222_X1 port map( A1 => n16612, A2 => n15030, B1 => n16609, B2 => 
                           n14326, C1 => n16606, C2 => n12045, ZN => n10789);
   U5039 : AOI221_X1 port map( B1 => registers_12_28_port, B2 => n16663, C1 => 
                           registers_15_28_port, C2 => n16660, A => n10781, ZN 
                           => n10780);
   U5040 : OAI22_X1 port map( A1 => n16657, A2 => n15069, B1 => n16654, B2 => 
                           n14423, ZN => n10781);
   U5041 : AOI221_X1 port map( B1 => net227416, B2 => n16567, C1 => 
                           registers_44_28_port, C2 => n16564, A => n10797, ZN 
                           => n10796);
   U5042 : OAI22_X1 port map( A1 => n16561, A2 => n15148, B1 => n16558, B2 => 
                           n14531, ZN => n10797);
   U5043 : AOI221_X1 port map( B1 => registers_56_28_port, B2 => n16519, C1 => 
                           registers_60_28_port, C2 => n16516, A => n10805, ZN 
                           => n10804);
   U5044 : OAI222_X1 port map( A1 => n16513, A2 => n14596, B1 => n16510, B2 => 
                           n12158, C1 => n16507, C2 => n15268, ZN => n10805);
   U5045 : AOI221_X1 port map( B1 => registers_2_29_port, B2 => n16618, C1 => 
                           registers_29_29_port, C2 => n16615, A => n10746, ZN 
                           => n10745);
   U5046 : OAI222_X1 port map( A1 => n16612, A2 => n15031, B1 => n16609, B2 => 
                           n14327, C1 => n16606, C2 => n12046, ZN => n10746);
   U5047 : AOI221_X1 port map( B1 => registers_12_29_port, B2 => n16663, C1 => 
                           registers_15_29_port, C2 => n16660, A => n10738, ZN 
                           => n10737);
   U5048 : OAI22_X1 port map( A1 => n16657, A2 => n15070, B1 => n16654, B2 => 
                           n14424, ZN => n10738);
   U5049 : AOI221_X1 port map( B1 => net227434, B2 => n16567, C1 => 
                           registers_44_29_port, C2 => n16564, A => n10754, ZN 
                           => n10753);
   U5050 : OAI22_X1 port map( A1 => n16561, A2 => n15149, B1 => n16558, B2 => 
                           n14532, ZN => n10754);
   U5051 : AOI221_X1 port map( B1 => registers_56_29_port, B2 => n16519, C1 => 
                           registers_60_29_port, C2 => n16516, A => n10762, ZN 
                           => n10761);
   U5052 : OAI222_X1 port map( A1 => n16513, A2 => n14597, B1 => n16510, B2 => 
                           n12159, C1 => n16507, C2 => n15269, ZN => n10762);
   U5053 : AOI221_X1 port map( B1 => registers_2_30_port, B2 => n16618, C1 => 
                           registers_29_30_port, C2 => n16615, A => n10691, ZN 
                           => n10690);
   U5054 : OAI222_X1 port map( A1 => n16612, A2 => n14857, B1 => n16609, B2 => 
                           n14054, C1 => n16606, C2 => n11904, ZN => n10691);
   U5055 : AOI221_X1 port map( B1 => registers_12_30_port, B2 => n16663, C1 => 
                           registers_15_30_port, C2 => n16660, A => n10679, ZN 
                           => n10678);
   U5056 : OAI22_X1 port map( A1 => n16657, A2 => n14870, B1 => n16654, B2 => 
                           n14060, ZN => n10679);
   U5057 : AOI221_X1 port map( B1 => net227452, B2 => n16567, C1 => 
                           registers_44_30_port, C2 => n16564, A => n10704, ZN 
                           => n10703);
   U5058 : OAI22_X1 port map( A1 => n16561, A2 => n14871, B1 => n16558, B2 => 
                           n14069, ZN => n10704);
   U5059 : AOI221_X1 port map( B1 => registers_56_30_port, B2 => n16519, C1 => 
                           registers_60_30_port, C2 => n16516, A => n10717, ZN 
                           => n10716);
   U5060 : OAI222_X1 port map( A1 => n16513, A2 => n14534, B1 => n16510, B2 => 
                           n12048, C1 => n16507, C2 => n15033, ZN => n10717);
   U5061 : AOI221_X1 port map( B1 => registers_2_31_port, B2 => n16618, C1 => 
                           registers_29_31_port, C2 => n16615, A => n10568, ZN 
                           => n10565);
   U5062 : OAI222_X1 port map( A1 => n16612, A2 => n15032, B1 => n16609, B2 => 
                           n14328, C1 => n16606, C2 => n12047, ZN => n10568);
   U5063 : AOI221_X1 port map( B1 => registers_12_31_port, B2 => n16663, C1 => 
                           registers_15_31_port, C2 => n16660, A => n10537, ZN 
                           => n10534);
   U5064 : OAI22_X1 port map( A1 => n16657, A2 => n15071, B1 => n16654, B2 => 
                           n14425, ZN => n10537);
   U5065 : AOI221_X1 port map( B1 => net227470, B2 => n16567, C1 => 
                           registers_44_31_port, C2 => n16564, A => n10602, ZN 
                           => n10599);
   U5066 : OAI22_X1 port map( A1 => n16561, A2 => n15150, B1 => n16558, B2 => 
                           n14533, ZN => n10602);
   U5067 : AOI221_X1 port map( B1 => registers_56_31_port, B2 => n16519, C1 => 
                           registers_60_31_port, C2 => n16516, A => n10634, ZN 
                           => n10631);
   U5068 : OAI222_X1 port map( A1 => n16513, A2 => n14535, B1 => n16510, B2 => 
                           n12049, C1 => n16507, C2 => n15034, ZN => n10634);
   U5069 : AOI221_X1 port map( B1 => registers_37_23_port, B2 => n17819, C1 => 
                           registers_0_23_port, C2 => n17816, A => n5281, ZN =>
                           n5280);
   U5070 : OAI22_X1 port map( A1 => n17813, A2 => n15662, B1 => n17810, B2 => 
                           n14700, ZN => n5281);
   U5071 : AOI221_X1 port map( B1 => registers_37_24_port, B2 => n17819, C1 => 
                           registers_0_24_port, C2 => n17816, A => n5116, ZN =>
                           n5115);
   U5072 : OAI22_X1 port map( A1 => n17813, A2 => n15663, B1 => n17810, B2 => 
                           n14701, ZN => n5116);
   U5073 : AOI221_X1 port map( B1 => registers_37_25_port, B2 => n17819, C1 => 
                           registers_0_25_port, C2 => n17816, A => n5002, ZN =>
                           n5001);
   U5074 : OAI22_X1 port map( A1 => n17813, A2 => n15664, B1 => n17810, B2 => 
                           n14702, ZN => n5002);
   U5075 : AOI221_X1 port map( B1 => registers_56_26_port, B2 => n17675, C1 => 
                           registers_55_26_port, C2 => n17672, A => n4910, ZN 
                           => n4909);
   U5076 : OAI22_X1 port map( A1 => n17669, A2 => n15428, B1 => n17666, B2 => 
                           n14703, ZN => n4910);
   U5077 : AOI221_X1 port map( B1 => registers_37_26_port, B2 => n17819, C1 => 
                           registers_0_26_port, C2 => n17816, A => n4880, ZN =>
                           n4879);
   U5078 : OAI22_X1 port map( A1 => n17813, A2 => n15665, B1 => n17810, B2 => 
                           n14704, ZN => n4880);
   U5079 : AOI221_X1 port map( B1 => registers_56_27_port, B2 => n17675, C1 => 
                           registers_55_27_port, C2 => n17672, A => n4779, ZN 
                           => n4778);
   U5080 : OAI22_X1 port map( A1 => n17669, A2 => n15429, B1 => n17666, B2 => 
                           n14705, ZN => n4779);
   U5081 : AOI221_X1 port map( B1 => registers_37_27_port, B2 => n17819, C1 => 
                           registers_0_27_port, C2 => n17816, A => n4751, ZN =>
                           n4750);
   U5082 : OAI22_X1 port map( A1 => n17813, A2 => n15666, B1 => n17810, B2 => 
                           n14706, ZN => n4751);
   U5083 : AOI221_X1 port map( B1 => registers_56_28_port, B2 => n17675, C1 => 
                           registers_55_28_port, C2 => n17672, A => n4650, ZN 
                           => n4649);
   U5084 : OAI22_X1 port map( A1 => n17669, A2 => n15430, B1 => n17666, B2 => 
                           n14707, ZN => n4650);
   U5085 : AOI221_X1 port map( B1 => registers_37_28_port, B2 => n17819, C1 => 
                           registers_0_28_port, C2 => n17816, A => n4622, ZN =>
                           n4621);
   U5086 : OAI22_X1 port map( A1 => n17813, A2 => n15667, B1 => n17810, B2 => 
                           n14708, ZN => n4622);
   U5087 : AOI221_X1 port map( B1 => registers_56_29_port, B2 => n17675, C1 => 
                           registers_55_29_port, C2 => n17672, A => n4521, ZN 
                           => n4520);
   U5088 : OAI22_X1 port map( A1 => n17669, A2 => n15431, B1 => n17666, B2 => 
                           n14709, ZN => n4521);
   U5089 : AOI221_X1 port map( B1 => registers_37_29_port, B2 => n17819, C1 => 
                           registers_0_29_port, C2 => n17816, A => n4489, ZN =>
                           n4488);
   U5090 : OAI22_X1 port map( A1 => n17813, A2 => n15668, B1 => n17810, B2 => 
                           n14710, ZN => n4489);
   U5091 : AOI221_X1 port map( B1 => registers_37_30_port, B2 => n17819, C1 => 
                           registers_0_30_port, C2 => n17816, A => n4109, ZN =>
                           n4106);
   U5092 : OAI22_X1 port map( A1 => n17813, A2 => n15280, B1 => n17810, B2 => 
                           n14629, ZN => n4109);
   U5093 : AOI221_X1 port map( B1 => registers_12_0_port, B2 => n16409, C1 => 
                           registers_17_0_port, C2 => n16406, A => n13916, ZN 
                           => n13915);
   U5094 : OAI22_X1 port map( A1 => n16403, A2 => n15072, B1 => n16400, B2 => 
                           n14426, ZN => n13916);
   U5095 : AOI221_X1 port map( B1 => net226850, B2 => n16313, C1 => 
                           registers_44_0_port, C2 => n16310, A => n13952, ZN 
                           => n13951);
   U5096 : OAI22_X1 port map( A1 => n16307, A2 => n15073, B1 => n16304, B2 => 
                           n14427, ZN => n13952);
   U5097 : AOI221_X1 port map( B1 => registers_12_1_port, B2 => n16409, C1 => 
                           registers_17_1_port, C2 => n16406, A => n13869, ZN 
                           => n13868);
   U5098 : OAI22_X1 port map( A1 => n16403, A2 => n15074, B1 => n16400, B2 => 
                           n14428, ZN => n13869);
   U5099 : AOI221_X1 port map( B1 => net226870, B2 => n16313, C1 => 
                           registers_44_1_port, C2 => n16310, A => n13885, ZN 
                           => n13884);
   U5100 : OAI22_X1 port map( A1 => n16307, A2 => n15075, B1 => n16304, B2 => 
                           n14429, ZN => n13885);
   U5101 : AOI221_X1 port map( B1 => registers_12_2_port, B2 => n16409, C1 => 
                           registers_17_2_port, C2 => n16406, A => n13827, ZN 
                           => n13826);
   U5102 : OAI22_X1 port map( A1 => n16403, A2 => n15076, B1 => n16400, B2 => 
                           n14430, ZN => n13827);
   U5103 : AOI221_X1 port map( B1 => net226883, B2 => n16313, C1 => 
                           registers_44_2_port, C2 => n16310, A => n13843, ZN 
                           => n13842);
   U5104 : OAI22_X1 port map( A1 => n16307, A2 => n15077, B1 => n16304, B2 => 
                           n14431, ZN => n13843);
   U5105 : AOI221_X1 port map( B1 => registers_12_3_port, B2 => n16409, C1 => 
                           registers_17_3_port, C2 => n16406, A => n13785, ZN 
                           => n13784);
   U5106 : OAI22_X1 port map( A1 => n16403, A2 => n14994, B1 => n16400, B2 => 
                           n14291, ZN => n13785);
   U5107 : AOI221_X1 port map( B1 => net226903, B2 => n16313, C1 => 
                           registers_44_3_port, C2 => n16310, A => n13801, ZN 
                           => n13800);
   U5108 : OAI22_X1 port map( A1 => n16307, A2 => n14995, B1 => n16304, B2 => 
                           n14292, ZN => n13801);
   U5109 : AOI221_X1 port map( B1 => registers_12_4_port, B2 => n16409, C1 => 
                           registers_17_4_port, C2 => n16406, A => n13743, ZN 
                           => n13742);
   U5110 : OAI22_X1 port map( A1 => n16403, A2 => n15078, B1 => n16400, B2 => 
                           n14432, ZN => n13743);
   U5111 : AOI221_X1 port map( B1 => net226976, B2 => n16313, C1 => 
                           registers_44_4_port, C2 => n16310, A => n13759, ZN 
                           => n13758);
   U5112 : OAI22_X1 port map( A1 => n16307, A2 => n15079, B1 => n16304, B2 => 
                           n14433, ZN => n13759);
   U5113 : AOI221_X1 port map( B1 => registers_12_5_port, B2 => n16409, C1 => 
                           registers_17_5_port, C2 => n16406, A => n13701, ZN 
                           => n13700);
   U5114 : OAI22_X1 port map( A1 => n16403, A2 => n15080, B1 => n16400, B2 => 
                           n14434, ZN => n13701);
   U5115 : AOI221_X1 port map( B1 => net226996, B2 => n16313, C1 => 
                           registers_44_5_port, C2 => n16310, A => n13717, ZN 
                           => n13716);
   U5116 : OAI22_X1 port map( A1 => n16307, A2 => n14996, B1 => n16304, B2 => 
                           n14293, ZN => n13717);
   U5117 : AOI221_X1 port map( B1 => registers_12_6_port, B2 => n16409, C1 => 
                           registers_17_6_port, C2 => n16406, A => n13659, ZN 
                           => n13658);
   U5118 : OAI22_X1 port map( A1 => n16403, A2 => n15081, B1 => n16400, B2 => 
                           n14435, ZN => n13659);
   U5119 : AOI221_X1 port map( B1 => net227020, B2 => n16313, C1 => 
                           registers_44_6_port, C2 => n16310, A => n13675, ZN 
                           => n13674);
   U5120 : OAI22_X1 port map( A1 => n16307, A2 => n15082, B1 => n16304, B2 => 
                           n14436, ZN => n13675);
   U5121 : AOI221_X1 port map( B1 => registers_12_7_port, B2 => n16409, C1 => 
                           registers_17_7_port, C2 => n16406, A => n13617, ZN 
                           => n13616);
   U5122 : OAI22_X1 port map( A1 => n16403, A2 => n15083, B1 => n16400, B2 => 
                           n14437, ZN => n13617);
   U5123 : AOI221_X1 port map( B1 => net227038, B2 => n16313, C1 => 
                           registers_44_7_port, C2 => n16310, A => n13633, ZN 
                           => n13632);
   U5124 : OAI22_X1 port map( A1 => n16307, A2 => n15084, B1 => n16304, B2 => 
                           n14438, ZN => n13633);
   U5125 : AOI221_X1 port map( B1 => registers_12_8_port, B2 => n16409, C1 => 
                           registers_17_8_port, C2 => n16406, A => n13575, ZN 
                           => n13574);
   U5126 : OAI22_X1 port map( A1 => n16403, A2 => n15085, B1 => n16400, B2 => 
                           n14439, ZN => n13575);
   U5127 : AOI221_X1 port map( B1 => net227056, B2 => n16313, C1 => 
                           registers_44_8_port, C2 => n16310, A => n13591, ZN 
                           => n13590);
   U5128 : OAI22_X1 port map( A1 => n16307, A2 => n15086, B1 => n16304, B2 => 
                           n14440, ZN => n13591);
   U5129 : AOI221_X1 port map( B1 => registers_12_9_port, B2 => n16409, C1 => 
                           registers_17_9_port, C2 => n16406, A => n13533, ZN 
                           => n13532);
   U5130 : OAI22_X1 port map( A1 => n16403, A2 => n15087, B1 => n16400, B2 => 
                           n14441, ZN => n13533);
   U5131 : AOI221_X1 port map( B1 => net227074, B2 => n16313, C1 => 
                           registers_44_9_port, C2 => n16310, A => n13549, ZN 
                           => n13548);
   U5132 : OAI22_X1 port map( A1 => n16307, A2 => n15088, B1 => n16304, B2 => 
                           n14442, ZN => n13549);
   U5133 : AOI221_X1 port map( B1 => registers_12_10_port, B2 => n16409, C1 => 
                           registers_17_10_port, C2 => n16406, A => n13491, ZN 
                           => n13490);
   U5134 : OAI22_X1 port map( A1 => n16403, A2 => n15089, B1 => n16400, B2 => 
                           n14443, ZN => n13491);
   U5135 : AOI221_X1 port map( B1 => net227092, B2 => n16313, C1 => 
                           registers_44_10_port, C2 => n16310, A => n13507, ZN 
                           => n13506);
   U5136 : OAI22_X1 port map( A1 => n16307, A2 => n15090, B1 => n16304, B2 => 
                           n14444, ZN => n13507);
   U5137 : AOI221_X1 port map( B1 => registers_12_11_port, B2 => n16409, C1 => 
                           registers_17_11_port, C2 => n16406, A => n13449, ZN 
                           => n13448);
   U5138 : OAI22_X1 port map( A1 => n16403, A2 => n15091, B1 => n16400, B2 => 
                           n14445, ZN => n13449);
   U5139 : AOI221_X1 port map( B1 => net227110, B2 => n16313, C1 => 
                           registers_44_11_port, C2 => n16310, A => n13465, ZN 
                           => n13464);
   U5140 : OAI22_X1 port map( A1 => n16307, A2 => n15092, B1 => n16304, B2 => 
                           n14446, ZN => n13465);
   U5141 : AOI221_X1 port map( B1 => registers_12_12_port, B2 => n16410, C1 => 
                           registers_17_12_port, C2 => n16407, A => n13407, ZN 
                           => n13406);
   U5142 : OAI22_X1 port map( A1 => n16404, A2 => n15093, B1 => n16401, B2 => 
                           n14447, ZN => n13407);
   U5143 : AOI221_X1 port map( B1 => net227128, B2 => n16314, C1 => 
                           registers_44_12_port, C2 => n16311, A => n13423, ZN 
                           => n13422);
   U5144 : OAI22_X1 port map( A1 => n16308, A2 => n15094, B1 => n16305, B2 => 
                           n14448, ZN => n13423);
   U5145 : AOI221_X1 port map( B1 => registers_12_13_port, B2 => n16410, C1 => 
                           registers_17_13_port, C2 => n16407, A => n13365, ZN 
                           => n13364);
   U5146 : OAI22_X1 port map( A1 => n16404, A2 => n15095, B1 => n16401, B2 => 
                           n14449, ZN => n13365);
   U5147 : AOI221_X1 port map( B1 => net227146, B2 => n16314, C1 => 
                           registers_44_13_port, C2 => n16311, A => n13381, ZN 
                           => n13380);
   U5148 : OAI22_X1 port map( A1 => n16308, A2 => n15096, B1 => n16305, B2 => 
                           n14450, ZN => n13381);
   U5149 : AOI221_X1 port map( B1 => registers_12_14_port, B2 => n16410, C1 => 
                           registers_17_14_port, C2 => n16407, A => n13323, ZN 
                           => n13322);
   U5150 : OAI22_X1 port map( A1 => n16404, A2 => n15097, B1 => n16401, B2 => 
                           n14451, ZN => n13323);
   U5151 : AOI221_X1 port map( B1 => net227164, B2 => n16314, C1 => 
                           registers_44_14_port, C2 => n16311, A => n13339, ZN 
                           => n13338);
   U5152 : OAI22_X1 port map( A1 => n16308, A2 => n15098, B1 => n16305, B2 => 
                           n14452, ZN => n13339);
   U5153 : AOI221_X1 port map( B1 => registers_12_15_port, B2 => n16410, C1 => 
                           registers_17_15_port, C2 => n16407, A => n13281, ZN 
                           => n13280);
   U5154 : OAI22_X1 port map( A1 => n16404, A2 => n15099, B1 => n16401, B2 => 
                           n14453, ZN => n13281);
   U5155 : AOI221_X1 port map( B1 => net227182, B2 => n16314, C1 => 
                           registers_44_15_port, C2 => n16311, A => n13297, ZN 
                           => n13296);
   U5156 : OAI22_X1 port map( A1 => n16308, A2 => n15100, B1 => n16305, B2 => 
                           n14454, ZN => n13297);
   U5157 : AOI221_X1 port map( B1 => registers_12_16_port, B2 => n16410, C1 => 
                           registers_17_16_port, C2 => n16407, A => n13239, ZN 
                           => n13238);
   U5158 : OAI22_X1 port map( A1 => n16404, A2 => n15101, B1 => n16401, B2 => 
                           n14455, ZN => n13239);
   U5159 : AOI221_X1 port map( B1 => net227200, B2 => n16314, C1 => 
                           registers_44_16_port, C2 => n16311, A => n13255, ZN 
                           => n13254);
   U5160 : OAI22_X1 port map( A1 => n16308, A2 => n15102, B1 => n16305, B2 => 
                           n14456, ZN => n13255);
   U5161 : AOI221_X1 port map( B1 => registers_12_17_port, B2 => n16410, C1 => 
                           registers_17_17_port, C2 => n16407, A => n13197, ZN 
                           => n13196);
   U5162 : OAI22_X1 port map( A1 => n16404, A2 => n15103, B1 => n16401, B2 => 
                           n14457, ZN => n13197);
   U5163 : AOI221_X1 port map( B1 => net227218, B2 => n16314, C1 => 
                           registers_44_17_port, C2 => n16311, A => n13213, ZN 
                           => n13212);
   U5164 : OAI22_X1 port map( A1 => n16308, A2 => n15104, B1 => n16305, B2 => 
                           n14458, ZN => n13213);
   U5165 : AOI221_X1 port map( B1 => registers_12_18_port, B2 => n16410, C1 => 
                           registers_17_18_port, C2 => n16407, A => n13155, ZN 
                           => n13154);
   U5166 : OAI22_X1 port map( A1 => n16404, A2 => n15105, B1 => n16401, B2 => 
                           n14459, ZN => n13155);
   U5167 : AOI221_X1 port map( B1 => net227236, B2 => n16314, C1 => 
                           registers_44_18_port, C2 => n16311, A => n13171, ZN 
                           => n13170);
   U5168 : OAI22_X1 port map( A1 => n16308, A2 => n15106, B1 => n16305, B2 => 
                           n14460, ZN => n13171);
   U5169 : AOI221_X1 port map( B1 => registers_12_19_port, B2 => n16410, C1 => 
                           registers_17_19_port, C2 => n16407, A => n13113, ZN 
                           => n13112);
   U5170 : OAI22_X1 port map( A1 => n16404, A2 => n15107, B1 => n16401, B2 => 
                           n14461, ZN => n13113);
   U5171 : AOI221_X1 port map( B1 => net227254, B2 => n16314, C1 => 
                           registers_44_19_port, C2 => n16311, A => n13129, ZN 
                           => n13128);
   U5172 : OAI22_X1 port map( A1 => n16308, A2 => n15108, B1 => n16305, B2 => 
                           n14462, ZN => n13129);
   U5173 : AOI221_X1 port map( B1 => registers_12_20_port, B2 => n16410, C1 => 
                           registers_17_20_port, C2 => n16407, A => n13071, ZN 
                           => n13070);
   U5174 : OAI22_X1 port map( A1 => n16404, A2 => n15109, B1 => n16401, B2 => 
                           n14463, ZN => n13071);
   U5175 : AOI221_X1 port map( B1 => net227272, B2 => n16314, C1 => 
                           registers_44_20_port, C2 => n16311, A => n13087, ZN 
                           => n13086);
   U5176 : OAI22_X1 port map( A1 => n16308, A2 => n15110, B1 => n16305, B2 => 
                           n14464, ZN => n13087);
   U5177 : AOI221_X1 port map( B1 => registers_12_21_port, B2 => n16410, C1 => 
                           registers_17_21_port, C2 => n16407, A => n13029, ZN 
                           => n13028);
   U5178 : OAI22_X1 port map( A1 => n16404, A2 => n15111, B1 => n16401, B2 => 
                           n14465, ZN => n13029);
   U5179 : AOI221_X1 port map( B1 => net227290, B2 => n16314, C1 => 
                           registers_44_21_port, C2 => n16311, A => n13045, ZN 
                           => n13044);
   U5180 : OAI22_X1 port map( A1 => n16308, A2 => n15112, B1 => n16305, B2 => 
                           n14466, ZN => n13045);
   U5181 : AOI221_X1 port map( B1 => registers_12_22_port, B2 => n16410, C1 => 
                           registers_17_22_port, C2 => n16407, A => n12987, ZN 
                           => n12986);
   U5182 : OAI22_X1 port map( A1 => n16404, A2 => n15113, B1 => n16401, B2 => 
                           n14467, ZN => n12987);
   U5183 : AOI221_X1 port map( B1 => net227308, B2 => n16314, C1 => 
                           registers_44_22_port, C2 => n16311, A => n13003, ZN 
                           => n13002);
   U5184 : OAI22_X1 port map( A1 => n16308, A2 => n15114, B1 => n16305, B2 => 
                           n14468, ZN => n13003);
   U5185 : AOI221_X1 port map( B1 => registers_12_23_port, B2 => n16410, C1 => 
                           registers_17_23_port, C2 => n16407, A => n12945, ZN 
                           => n12944);
   U5186 : OAI22_X1 port map( A1 => n16404, A2 => n15115, B1 => n16401, B2 => 
                           n14469, ZN => n12945);
   U5187 : AOI221_X1 port map( B1 => net227326, B2 => n16314, C1 => 
                           registers_44_23_port, C2 => n16311, A => n12961, ZN 
                           => n12960);
   U5188 : OAI22_X1 port map( A1 => n16308, A2 => n15116, B1 => n16305, B2 => 
                           n14470, ZN => n12961);
   U5189 : AOI221_X1 port map( B1 => registers_12_0_port, B2 => n16661, C1 => 
                           registers_15_0_port, C2 => n16658, A => n12435, ZN 
                           => n12434);
   U5190 : OAI22_X1 port map( A1 => n16655, A2 => n15072, B1 => n16652, B2 => 
                           n14426, ZN => n12435);
   U5191 : AOI221_X1 port map( B1 => net226850, B2 => n16565, C1 => 
                           registers_44_0_port, C2 => n16562, A => n12471, ZN 
                           => n12470);
   U5192 : OAI22_X1 port map( A1 => n16559, A2 => n15073, B1 => n16556, B2 => 
                           n14427, ZN => n12471);
   U5193 : AOI221_X1 port map( B1 => registers_12_1_port, B2 => n16661, C1 => 
                           registers_15_1_port, C2 => n16658, A => n12273, ZN 
                           => n12272);
   U5194 : OAI22_X1 port map( A1 => n16655, A2 => n15074, B1 => n16652, B2 => 
                           n14428, ZN => n12273);
   U5195 : AOI221_X1 port map( B1 => net226870, B2 => n16565, C1 => 
                           registers_44_1_port, C2 => n16562, A => n12289, ZN 
                           => n12288);
   U5196 : OAI22_X1 port map( A1 => n16559, A2 => n15075, B1 => n16556, B2 => 
                           n14429, ZN => n12289);
   U5197 : AOI221_X1 port map( B1 => registers_12_2_port, B2 => n16661, C1 => 
                           registers_15_2_port, C2 => n16658, A => n12120, ZN 
                           => n12119);
   U5198 : OAI22_X1 port map( A1 => n16655, A2 => n15076, B1 => n16652, B2 => 
                           n14430, ZN => n12120);
   U5199 : AOI221_X1 port map( B1 => net226883, B2 => n16565, C1 => 
                           registers_44_2_port, C2 => n16562, A => n12136, ZN 
                           => n12135);
   U5200 : OAI22_X1 port map( A1 => n16559, A2 => n15077, B1 => n16556, B2 => 
                           n14431, ZN => n12136);
   U5201 : AOI221_X1 port map( B1 => registers_12_3_port, B2 => n16661, C1 => 
                           registers_15_3_port, C2 => n16658, A => n11967, ZN 
                           => n11966);
   U5202 : OAI22_X1 port map( A1 => n16655, A2 => n14994, B1 => n16652, B2 => 
                           n14291, ZN => n11967);
   U5203 : AOI221_X1 port map( B1 => net226903, B2 => n16565, C1 => 
                           registers_44_3_port, C2 => n16562, A => n11983, ZN 
                           => n11982);
   U5204 : OAI22_X1 port map( A1 => n16559, A2 => n14995, B1 => n16556, B2 => 
                           n14292, ZN => n11983);
   U5205 : AOI221_X1 port map( B1 => registers_12_4_port, B2 => n16661, C1 => 
                           registers_15_4_port, C2 => n16658, A => n11814, ZN 
                           => n11813);
   U5206 : OAI22_X1 port map( A1 => n16655, A2 => n15078, B1 => n16652, B2 => 
                           n14432, ZN => n11814);
   U5207 : AOI221_X1 port map( B1 => net226976, B2 => n16565, C1 => 
                           registers_44_4_port, C2 => n16562, A => n11830, ZN 
                           => n11829);
   U5208 : OAI22_X1 port map( A1 => n16559, A2 => n15079, B1 => n16556, B2 => 
                           n14433, ZN => n11830);
   U5209 : AOI221_X1 port map( B1 => registers_12_5_port, B2 => n16661, C1 => 
                           registers_15_5_port, C2 => n16658, A => n11771, ZN 
                           => n11770);
   U5210 : OAI22_X1 port map( A1 => n16655, A2 => n15080, B1 => n16652, B2 => 
                           n14434, ZN => n11771);
   U5211 : AOI221_X1 port map( B1 => net226996, B2 => n16565, C1 => 
                           registers_44_5_port, C2 => n16562, A => n11787, ZN 
                           => n11786);
   U5212 : OAI22_X1 port map( A1 => n16559, A2 => n14996, B1 => n16556, B2 => 
                           n14293, ZN => n11787);
   U5213 : AOI221_X1 port map( B1 => registers_12_6_port, B2 => n16661, C1 => 
                           registers_15_6_port, C2 => n16658, A => n11728, ZN 
                           => n11727);
   U5214 : OAI22_X1 port map( A1 => n16655, A2 => n15081, B1 => n16652, B2 => 
                           n14435, ZN => n11728);
   U5215 : AOI221_X1 port map( B1 => net227020, B2 => n16565, C1 => 
                           registers_44_6_port, C2 => n16562, A => n11744, ZN 
                           => n11743);
   U5216 : OAI22_X1 port map( A1 => n16559, A2 => n15082, B1 => n16556, B2 => 
                           n14436, ZN => n11744);
   U5217 : AOI221_X1 port map( B1 => registers_12_7_port, B2 => n16661, C1 => 
                           registers_15_7_port, C2 => n16658, A => n11685, ZN 
                           => n11684);
   U5218 : OAI22_X1 port map( A1 => n16655, A2 => n15083, B1 => n16652, B2 => 
                           n14437, ZN => n11685);
   U5219 : AOI221_X1 port map( B1 => net227038, B2 => n16565, C1 => 
                           registers_44_7_port, C2 => n16562, A => n11701, ZN 
                           => n11700);
   U5220 : OAI22_X1 port map( A1 => n16559, A2 => n15084, B1 => n16556, B2 => 
                           n14438, ZN => n11701);
   U5221 : AOI221_X1 port map( B1 => registers_12_8_port, B2 => n16661, C1 => 
                           registers_15_8_port, C2 => n16658, A => n11642, ZN 
                           => n11641);
   U5222 : OAI22_X1 port map( A1 => n16655, A2 => n15085, B1 => n16652, B2 => 
                           n14439, ZN => n11642);
   U5223 : AOI221_X1 port map( B1 => net227056, B2 => n16565, C1 => 
                           registers_44_8_port, C2 => n16562, A => n11658, ZN 
                           => n11657);
   U5224 : OAI22_X1 port map( A1 => n16559, A2 => n15086, B1 => n16556, B2 => 
                           n14440, ZN => n11658);
   U5225 : AOI221_X1 port map( B1 => registers_12_9_port, B2 => n16661, C1 => 
                           registers_15_9_port, C2 => n16658, A => n11599, ZN 
                           => n11598);
   U5226 : OAI22_X1 port map( A1 => n16655, A2 => n15087, B1 => n16652, B2 => 
                           n14441, ZN => n11599);
   U5227 : AOI221_X1 port map( B1 => net227074, B2 => n16565, C1 => 
                           registers_44_9_port, C2 => n16562, A => n11615, ZN 
                           => n11614);
   U5228 : OAI22_X1 port map( A1 => n16559, A2 => n15088, B1 => n16556, B2 => 
                           n14442, ZN => n11615);
   U5229 : AOI221_X1 port map( B1 => registers_12_10_port, B2 => n16661, C1 => 
                           registers_15_10_port, C2 => n16658, A => n11556, ZN 
                           => n11555);
   U5230 : OAI22_X1 port map( A1 => n16655, A2 => n15089, B1 => n16652, B2 => 
                           n14443, ZN => n11556);
   U5231 : AOI221_X1 port map( B1 => net227092, B2 => n16565, C1 => 
                           registers_44_10_port, C2 => n16562, A => n11572, ZN 
                           => n11571);
   U5232 : OAI22_X1 port map( A1 => n16559, A2 => n15090, B1 => n16556, B2 => 
                           n14444, ZN => n11572);
   U5233 : AOI221_X1 port map( B1 => registers_12_11_port, B2 => n16661, C1 => 
                           registers_15_11_port, C2 => n16658, A => n11513, ZN 
                           => n11512);
   U5234 : OAI22_X1 port map( A1 => n16655, A2 => n15091, B1 => n16652, B2 => 
                           n14445, ZN => n11513);
   U5235 : AOI221_X1 port map( B1 => net227110, B2 => n16565, C1 => 
                           registers_44_11_port, C2 => n16562, A => n11529, ZN 
                           => n11528);
   U5236 : OAI22_X1 port map( A1 => n16559, A2 => n15092, B1 => n16556, B2 => 
                           n14446, ZN => n11529);
   U5237 : AOI221_X1 port map( B1 => registers_12_12_port, B2 => n16662, C1 => 
                           registers_15_12_port, C2 => n16659, A => n11470, ZN 
                           => n11469);
   U5238 : OAI22_X1 port map( A1 => n16656, A2 => n15093, B1 => n16653, B2 => 
                           n14447, ZN => n11470);
   U5239 : AOI221_X1 port map( B1 => net227128, B2 => n16566, C1 => 
                           registers_44_12_port, C2 => n16563, A => n11486, ZN 
                           => n11485);
   U5240 : OAI22_X1 port map( A1 => n16560, A2 => n15094, B1 => n16557, B2 => 
                           n14448, ZN => n11486);
   U5241 : AOI221_X1 port map( B1 => registers_12_13_port, B2 => n16662, C1 => 
                           registers_15_13_port, C2 => n16659, A => n11426, ZN 
                           => n11425);
   U5242 : OAI22_X1 port map( A1 => n16656, A2 => n15095, B1 => n16653, B2 => 
                           n14449, ZN => n11426);
   U5243 : AOI221_X1 port map( B1 => net227146, B2 => n16566, C1 => 
                           registers_44_13_port, C2 => n16563, A => n11442, ZN 
                           => n11441);
   U5244 : OAI22_X1 port map( A1 => n16560, A2 => n15096, B1 => n16557, B2 => 
                           n14450, ZN => n11442);
   U5245 : AOI221_X1 port map( B1 => registers_12_14_port, B2 => n16662, C1 => 
                           registers_15_14_port, C2 => n16659, A => n11383, ZN 
                           => n11382);
   U5246 : OAI22_X1 port map( A1 => n16656, A2 => n15097, B1 => n16653, B2 => 
                           n14451, ZN => n11383);
   U5247 : AOI221_X1 port map( B1 => net227164, B2 => n16566, C1 => 
                           registers_44_14_port, C2 => n16563, A => n11399, ZN 
                           => n11398);
   U5248 : OAI22_X1 port map( A1 => n16560, A2 => n15098, B1 => n16557, B2 => 
                           n14452, ZN => n11399);
   U5249 : AOI221_X1 port map( B1 => registers_12_15_port, B2 => n16662, C1 => 
                           registers_15_15_port, C2 => n16659, A => n11340, ZN 
                           => n11339);
   U5250 : OAI22_X1 port map( A1 => n16656, A2 => n15099, B1 => n16653, B2 => 
                           n14453, ZN => n11340);
   U5251 : AOI221_X1 port map( B1 => net227182, B2 => n16566, C1 => 
                           registers_44_15_port, C2 => n16563, A => n11356, ZN 
                           => n11355);
   U5252 : OAI22_X1 port map( A1 => n16560, A2 => n15100, B1 => n16557, B2 => 
                           n14454, ZN => n11356);
   U5253 : AOI221_X1 port map( B1 => registers_12_16_port, B2 => n16662, C1 => 
                           registers_15_16_port, C2 => n16659, A => n11297, ZN 
                           => n11296);
   U5254 : OAI22_X1 port map( A1 => n16656, A2 => n15101, B1 => n16653, B2 => 
                           n14455, ZN => n11297);
   U5255 : AOI221_X1 port map( B1 => net227200, B2 => n16566, C1 => 
                           registers_44_16_port, C2 => n16563, A => n11313, ZN 
                           => n11312);
   U5256 : OAI22_X1 port map( A1 => n16560, A2 => n15102, B1 => n16557, B2 => 
                           n14456, ZN => n11313);
   U5257 : AOI221_X1 port map( B1 => registers_12_17_port, B2 => n16662, C1 => 
                           registers_15_17_port, C2 => n16659, A => n11254, ZN 
                           => n11253);
   U5258 : OAI22_X1 port map( A1 => n16656, A2 => n15103, B1 => n16653, B2 => 
                           n14457, ZN => n11254);
   U5259 : AOI221_X1 port map( B1 => net227218, B2 => n16566, C1 => 
                           registers_44_17_port, C2 => n16563, A => n11270, ZN 
                           => n11269);
   U5260 : OAI22_X1 port map( A1 => n16560, A2 => n15104, B1 => n16557, B2 => 
                           n14458, ZN => n11270);
   U5261 : AOI221_X1 port map( B1 => registers_12_18_port, B2 => n16662, C1 => 
                           registers_15_18_port, C2 => n16659, A => n11211, ZN 
                           => n11210);
   U5262 : OAI22_X1 port map( A1 => n16656, A2 => n15105, B1 => n16653, B2 => 
                           n14459, ZN => n11211);
   U5263 : AOI221_X1 port map( B1 => net227236, B2 => n16566, C1 => 
                           registers_44_18_port, C2 => n16563, A => n11227, ZN 
                           => n11226);
   U5264 : OAI22_X1 port map( A1 => n16560, A2 => n15106, B1 => n16557, B2 => 
                           n14460, ZN => n11227);
   U5265 : AOI221_X1 port map( B1 => registers_12_19_port, B2 => n16662, C1 => 
                           registers_15_19_port, C2 => n16659, A => n11168, ZN 
                           => n11167);
   U5266 : OAI22_X1 port map( A1 => n16656, A2 => n15107, B1 => n16653, B2 => 
                           n14461, ZN => n11168);
   U5267 : AOI221_X1 port map( B1 => net227254, B2 => n16566, C1 => 
                           registers_44_19_port, C2 => n16563, A => n11184, ZN 
                           => n11183);
   U5268 : OAI22_X1 port map( A1 => n16560, A2 => n15108, B1 => n16557, B2 => 
                           n14462, ZN => n11184);
   U5269 : AOI221_X1 port map( B1 => registers_12_20_port, B2 => n16662, C1 => 
                           registers_15_20_port, C2 => n16659, A => n11125, ZN 
                           => n11124);
   U5270 : OAI22_X1 port map( A1 => n16656, A2 => n15109, B1 => n16653, B2 => 
                           n14463, ZN => n11125);
   U5271 : AOI221_X1 port map( B1 => net227272, B2 => n16566, C1 => 
                           registers_44_20_port, C2 => n16563, A => n11141, ZN 
                           => n11140);
   U5272 : OAI22_X1 port map( A1 => n16560, A2 => n15110, B1 => n16557, B2 => 
                           n14464, ZN => n11141);
   U5273 : AOI221_X1 port map( B1 => registers_12_21_port, B2 => n16662, C1 => 
                           registers_15_21_port, C2 => n16659, A => n11082, ZN 
                           => n11081);
   U5274 : OAI22_X1 port map( A1 => n16656, A2 => n15111, B1 => n16653, B2 => 
                           n14465, ZN => n11082);
   U5275 : AOI221_X1 port map( B1 => net227290, B2 => n16566, C1 => 
                           registers_44_21_port, C2 => n16563, A => n11098, ZN 
                           => n11097);
   U5276 : OAI22_X1 port map( A1 => n16560, A2 => n15112, B1 => n16557, B2 => 
                           n14466, ZN => n11098);
   U5277 : AOI221_X1 port map( B1 => registers_12_22_port, B2 => n16662, C1 => 
                           registers_15_22_port, C2 => n16659, A => n11039, ZN 
                           => n11038);
   U5278 : OAI22_X1 port map( A1 => n16656, A2 => n15113, B1 => n16653, B2 => 
                           n14467, ZN => n11039);
   U5279 : AOI221_X1 port map( B1 => net227308, B2 => n16566, C1 => 
                           registers_44_22_port, C2 => n16563, A => n11055, ZN 
                           => n11054);
   U5280 : OAI22_X1 port map( A1 => n16560, A2 => n15114, B1 => n16557, B2 => 
                           n14468, ZN => n11055);
   U5281 : AOI221_X1 port map( B1 => registers_12_23_port, B2 => n16662, C1 => 
                           registers_15_23_port, C2 => n16659, A => n10996, ZN 
                           => n10995);
   U5282 : OAI22_X1 port map( A1 => n16656, A2 => n15115, B1 => n16653, B2 => 
                           n14469, ZN => n10996);
   U5283 : AOI221_X1 port map( B1 => net227326, B2 => n16566, C1 => 
                           registers_44_23_port, C2 => n16563, A => n11012, ZN 
                           => n11011);
   U5284 : OAI22_X1 port map( A1 => n16560, A2 => n15116, B1 => n16557, B2 => 
                           n14470, ZN => n11012);
   U5285 : AOI221_X1 port map( B1 => registers_56_0_port, B2 => n17673, C1 => 
                           registers_55_0_port, C2 => n17670, A => n12403, ZN 
                           => n12402);
   U5286 : OAI22_X1 port map( A1 => n17667, A2 => n15432, B1 => n17664, B2 => 
                           n14711, ZN => n12403);
   U5287 : AOI221_X1 port map( B1 => registers_37_0_port, B2 => n17817, C1 => 
                           registers_0_0_port, C2 => n17814, A => n12379, ZN =>
                           n12378);
   U5288 : OAI22_X1 port map( A1 => n17811, A2 => n15669, B1 => n17808, B2 => 
                           n14712, ZN => n12379);
   U5289 : AOI221_X1 port map( B1 => registers_56_1_port, B2 => n17673, C1 => 
                           registers_55_1_port, C2 => n17670, A => n12249, ZN 
                           => n12248);
   U5290 : OAI22_X1 port map( A1 => n17667, A2 => n15433, B1 => n17664, B2 => 
                           n14713, ZN => n12249);
   U5291 : AOI221_X1 port map( B1 => registers_37_1_port, B2 => n17817, C1 => 
                           registers_0_1_port, C2 => n17814, A => n12225, ZN =>
                           n12224);
   U5292 : OAI22_X1 port map( A1 => n17811, A2 => n15670, B1 => n17808, B2 => 
                           n14714, ZN => n12225);
   U5293 : AOI221_X1 port map( B1 => registers_56_2_port, B2 => n17673, C1 => 
                           registers_55_2_port, C2 => n17670, A => n12094, ZN 
                           => n12093);
   U5294 : OAI22_X1 port map( A1 => n17667, A2 => n15434, B1 => n17664, B2 => 
                           n14715, ZN => n12094);
   U5295 : AOI221_X1 port map( B1 => registers_37_2_port, B2 => n17817, C1 => 
                           registers_0_2_port, C2 => n17814, A => n12070, ZN =>
                           n12069);
   U5296 : OAI22_X1 port map( A1 => n17811, A2 => n15671, B1 => n17808, B2 => 
                           n14716, ZN => n12070);
   U5297 : AOI221_X1 port map( B1 => registers_56_3_port, B2 => n17673, C1 => 
                           registers_55_3_port, C2 => n17670, A => n11941, ZN 
                           => n11940);
   U5298 : OAI22_X1 port map( A1 => n17667, A2 => n15353, B1 => n17664, B2 => 
                           n14717, ZN => n11941);
   U5299 : AOI221_X1 port map( B1 => registers_37_3_port, B2 => n17817, C1 => 
                           registers_0_3_port, C2 => n17814, A => n11917, ZN =>
                           n11916);
   U5300 : OAI22_X1 port map( A1 => n17811, A2 => n15365, B1 => n17808, B2 => 
                           n14640, ZN => n11917);
   U5301 : AOI221_X1 port map( B1 => registers_56_4_port, B2 => n17673, C1 => 
                           registers_55_4_port, C2 => n17670, A => n10498, ZN 
                           => n10497);
   U5302 : OAI22_X1 port map( A1 => n17667, A2 => n15354, B1 => n17664, B2 => 
                           n14718, ZN => n10498);
   U5303 : AOI221_X1 port map( B1 => registers_37_4_port, B2 => n17817, C1 => 
                           registers_0_4_port, C2 => n17814, A => n10474, ZN =>
                           n10473);
   U5304 : OAI22_X1 port map( A1 => n17811, A2 => n15672, B1 => n17808, B2 => 
                           n14719, ZN => n10474);
   U5305 : AOI221_X1 port map( B1 => registers_56_5_port, B2 => n17673, C1 => 
                           registers_55_5_port, C2 => n17670, A => n10388, ZN 
                           => n10387);
   U5306 : OAI22_X1 port map( A1 => n17667, A2 => n15355, B1 => n17664, B2 => 
                           n14720, ZN => n10388);
   U5307 : AOI221_X1 port map( B1 => registers_37_5_port, B2 => n17817, C1 => 
                           registers_0_5_port, C2 => n17814, A => n10364, ZN =>
                           n10363);
   U5308 : OAI22_X1 port map( A1 => n17811, A2 => n15673, B1 => n17808, B2 => 
                           n14721, ZN => n10364);
   U5309 : AOI221_X1 port map( B1 => registers_56_6_port, B2 => n17673, C1 => 
                           registers_55_6_port, C2 => n17670, A => n10276, ZN 
                           => n10275);
   U5310 : OAI22_X1 port map( A1 => n17667, A2 => n15435, B1 => n17664, B2 => 
                           n14722, ZN => n10276);
   U5311 : AOI221_X1 port map( B1 => registers_37_6_port, B2 => n17817, C1 => 
                           registers_0_6_port, C2 => n17814, A => n10252, ZN =>
                           n10251);
   U5312 : OAI22_X1 port map( A1 => n17811, A2 => n15674, B1 => n17808, B2 => 
                           n14723, ZN => n10252);
   U5313 : AOI221_X1 port map( B1 => registers_56_7_port, B2 => n17673, C1 => 
                           registers_55_7_port, C2 => n17670, A => n7640, ZN =>
                           n7639);
   U5314 : OAI22_X1 port map( A1 => n17667, A2 => n15436, B1 => n17664, B2 => 
                           n14724, ZN => n7640);
   U5315 : AOI221_X1 port map( B1 => registers_37_7_port, B2 => n17817, C1 => 
                           registers_0_7_port, C2 => n17814, A => n7616, ZN => 
                           n7615);
   U5316 : OAI22_X1 port map( A1 => n17811, A2 => n15675, B1 => n17808, B2 => 
                           n14725, ZN => n7616);
   U5317 : AOI221_X1 port map( B1 => registers_56_8_port, B2 => n17673, C1 => 
                           registers_55_8_port, C2 => n17670, A => n7525, ZN =>
                           n7524);
   U5318 : OAI22_X1 port map( A1 => n17667, A2 => n15437, B1 => n17664, B2 => 
                           n14726, ZN => n7525);
   U5319 : AOI221_X1 port map( B1 => registers_37_8_port, B2 => n17817, C1 => 
                           registers_0_8_port, C2 => n17814, A => n7501, ZN => 
                           n7500);
   U5320 : OAI22_X1 port map( A1 => n17811, A2 => n15676, B1 => n17808, B2 => 
                           n14727, ZN => n7501);
   U5321 : AOI221_X1 port map( B1 => registers_56_9_port, B2 => n17673, C1 => 
                           registers_55_9_port, C2 => n17670, A => n7416, ZN =>
                           n7415);
   U5322 : OAI22_X1 port map( A1 => n17667, A2 => n15438, B1 => n17664, B2 => 
                           n14728, ZN => n7416);
   U5323 : AOI221_X1 port map( B1 => registers_37_9_port, B2 => n17817, C1 => 
                           registers_0_9_port, C2 => n17814, A => n7392, ZN => 
                           n7391);
   U5324 : OAI22_X1 port map( A1 => n17811, A2 => n15677, B1 => n17808, B2 => 
                           n14729, ZN => n7392);
   U5325 : AOI221_X1 port map( B1 => registers_56_10_port, B2 => n17673, C1 => 
                           registers_55_10_port, C2 => n17670, A => n7307, ZN 
                           => n7306);
   U5326 : OAI22_X1 port map( A1 => n17667, A2 => n15439, B1 => n17664, B2 => 
                           n14730, ZN => n7307);
   U5327 : AOI221_X1 port map( B1 => registers_37_10_port, B2 => n17817, C1 => 
                           registers_0_10_port, C2 => n17814, A => n7283, ZN =>
                           n7282);
   U5328 : OAI22_X1 port map( A1 => n17811, A2 => n15678, B1 => n17808, B2 => 
                           n14731, ZN => n7283);
   U5329 : AOI221_X1 port map( B1 => registers_56_11_port, B2 => n17674, C1 => 
                           registers_55_11_port, C2 => n17671, A => n7193, ZN 
                           => n7192);
   U5330 : OAI22_X1 port map( A1 => n17668, A2 => n15440, B1 => n17665, B2 => 
                           n14732, ZN => n7193);
   U5331 : AOI221_X1 port map( B1 => registers_37_11_port, B2 => n17818, C1 => 
                           registers_0_11_port, C2 => n17815, A => n7169, ZN =>
                           n7168);
   U5332 : OAI22_X1 port map( A1 => n17812, A2 => n15679, B1 => n17809, B2 => 
                           n14733, ZN => n7169);
   U5333 : AOI221_X1 port map( B1 => registers_56_12_port, B2 => n17674, C1 => 
                           registers_55_12_port, C2 => n17671, A => n7084, ZN 
                           => n7083);
   U5334 : OAI22_X1 port map( A1 => n17668, A2 => n15441, B1 => n17665, B2 => 
                           n14734, ZN => n7084);
   U5335 : AOI221_X1 port map( B1 => registers_37_12_port, B2 => n17818, C1 => 
                           registers_0_12_port, C2 => n17815, A => n7060, ZN =>
                           n7059);
   U5336 : OAI22_X1 port map( A1 => n17812, A2 => n15680, B1 => n17809, B2 => 
                           n14735, ZN => n7060);
   U5337 : AOI221_X1 port map( B1 => registers_56_13_port, B2 => n17674, C1 => 
                           registers_55_13_port, C2 => n17671, A => n6975, ZN 
                           => n6974);
   U5338 : OAI22_X1 port map( A1 => n17668, A2 => n15442, B1 => n17665, B2 => 
                           n14736, ZN => n6975);
   U5339 : AOI221_X1 port map( B1 => registers_37_13_port, B2 => n17818, C1 => 
                           registers_0_13_port, C2 => n17815, A => n6951, ZN =>
                           n6950);
   U5340 : OAI22_X1 port map( A1 => n17812, A2 => n15681, B1 => n17809, B2 => 
                           n14737, ZN => n6951);
   U5341 : AOI221_X1 port map( B1 => registers_56_14_port, B2 => n17674, C1 => 
                           registers_55_14_port, C2 => n17671, A => n6866, ZN 
                           => n6865);
   U5342 : OAI22_X1 port map( A1 => n17668, A2 => n15443, B1 => n17665, B2 => 
                           n14738, ZN => n6866);
   U5343 : AOI221_X1 port map( B1 => registers_37_14_port, B2 => n17818, C1 => 
                           registers_0_14_port, C2 => n17815, A => n6842, ZN =>
                           n6841);
   U5344 : OAI22_X1 port map( A1 => n17812, A2 => n15682, B1 => n17809, B2 => 
                           n14739, ZN => n6842);
   U5345 : AOI221_X1 port map( B1 => registers_56_15_port, B2 => n17674, C1 => 
                           registers_55_15_port, C2 => n17671, A => n6757, ZN 
                           => n6756);
   U5346 : OAI22_X1 port map( A1 => n17668, A2 => n15444, B1 => n17665, B2 => 
                           n14740, ZN => n6757);
   U5347 : AOI221_X1 port map( B1 => registers_37_15_port, B2 => n17818, C1 => 
                           registers_0_15_port, C2 => n17815, A => n6733, ZN =>
                           n6732);
   U5348 : OAI22_X1 port map( A1 => n17812, A2 => n15683, B1 => n17809, B2 => 
                           n14741, ZN => n6733);
   U5349 : AOI221_X1 port map( B1 => registers_56_16_port, B2 => n17674, C1 => 
                           registers_55_16_port, C2 => n17671, A => n6617, ZN 
                           => n6616);
   U5350 : OAI22_X1 port map( A1 => n17668, A2 => n15445, B1 => n17665, B2 => 
                           n14742, ZN => n6617);
   U5351 : AOI221_X1 port map( B1 => registers_37_16_port, B2 => n17818, C1 => 
                           registers_0_16_port, C2 => n17815, A => n6573, ZN =>
                           n6572);
   U5352 : OAI22_X1 port map( A1 => n17812, A2 => n15684, B1 => n17809, B2 => 
                           n14743, ZN => n6573);
   U5353 : AOI221_X1 port map( B1 => registers_56_17_port, B2 => n17674, C1 => 
                           registers_55_17_port, C2 => n17671, A => n6430, ZN 
                           => n6429);
   U5354 : OAI22_X1 port map( A1 => n17668, A2 => n15446, B1 => n17665, B2 => 
                           n14744, ZN => n6430);
   U5355 : AOI221_X1 port map( B1 => registers_37_17_port, B2 => n17818, C1 => 
                           registers_0_17_port, C2 => n17815, A => n6386, ZN =>
                           n6385);
   U5356 : OAI22_X1 port map( A1 => n17812, A2 => n15685, B1 => n17809, B2 => 
                           n14745, ZN => n6386);
   U5357 : AOI221_X1 port map( B1 => registers_56_18_port, B2 => n17674, C1 => 
                           registers_55_18_port, C2 => n17671, A => n6245, ZN 
                           => n6244);
   U5358 : OAI22_X1 port map( A1 => n17668, A2 => n15447, B1 => n17665, B2 => 
                           n14746, ZN => n6245);
   U5359 : AOI221_X1 port map( B1 => registers_37_18_port, B2 => n17818, C1 => 
                           registers_0_18_port, C2 => n17815, A => n6199, ZN =>
                           n6198);
   U5360 : OAI22_X1 port map( A1 => n17812, A2 => n15686, B1 => n17809, B2 => 
                           n14747, ZN => n6199);
   U5361 : AOI221_X1 port map( B1 => registers_56_19_port, B2 => n17674, C1 => 
                           registers_55_19_port, C2 => n17671, A => n6059, ZN 
                           => n6058);
   U5362 : OAI22_X1 port map( A1 => n17668, A2 => n15448, B1 => n17665, B2 => 
                           n14748, ZN => n6059);
   U5363 : AOI221_X1 port map( B1 => registers_37_19_port, B2 => n17818, C1 => 
                           registers_0_19_port, C2 => n17815, A => n6014, ZN =>
                           n6013);
   U5364 : OAI22_X1 port map( A1 => n17812, A2 => n15687, B1 => n17809, B2 => 
                           n14749, ZN => n6014);
   U5365 : AOI221_X1 port map( B1 => registers_56_20_port, B2 => n17674, C1 => 
                           registers_55_20_port, C2 => n17671, A => n5872, ZN 
                           => n5871);
   U5366 : OAI22_X1 port map( A1 => n17668, A2 => n15449, B1 => n17665, B2 => 
                           n14750, ZN => n5872);
   U5367 : AOI221_X1 port map( B1 => registers_37_20_port, B2 => n17818, C1 => 
                           registers_0_20_port, C2 => n17815, A => n5842, ZN =>
                           n5826);
   U5368 : OAI22_X1 port map( A1 => n17812, A2 => n15688, B1 => n17809, B2 => 
                           n14751, ZN => n5842);
   U5369 : AOI221_X1 port map( B1 => registers_56_21_port, B2 => n17674, C1 => 
                           registers_55_21_port, C2 => n17671, A => n5686, ZN 
                           => n5684);
   U5370 : OAI22_X1 port map( A1 => n17668, A2 => n15450, B1 => n17665, B2 => 
                           n14752, ZN => n5686);
   U5371 : AOI221_X1 port map( B1 => registers_37_21_port, B2 => n17818, C1 => 
                           registers_0_21_port, C2 => n17815, A => n5655, ZN =>
                           n5654);
   U5372 : OAI22_X1 port map( A1 => n17812, A2 => n15689, B1 => n17809, B2 => 
                           n14753, ZN => n5655);
   U5373 : AOI221_X1 port map( B1 => registers_56_22_port, B2 => n17674, C1 => 
                           registers_55_22_port, C2 => n17671, A => n5501, ZN 
                           => n5499);
   U5374 : OAI22_X1 port map( A1 => n17668, A2 => n15451, B1 => n17665, B2 => 
                           n14754, ZN => n5501);
   U5375 : AOI221_X1 port map( B1 => registers_37_22_port, B2 => n17818, C1 => 
                           registers_0_22_port, C2 => n17815, A => n5468, ZN =>
                           n5467);
   U5376 : OAI22_X1 port map( A1 => n17812, A2 => n15690, B1 => n17809, B2 => 
                           n14755, ZN => n5468);
   U5377 : AOI221_X1 port map( B1 => registers_56_31_port, B2 => n17673, C1 => 
                           registers_55_31_port, C2 => n17670, A => n14191, ZN 
                           => n14190);
   U5378 : OAI22_X1 port map( A1 => n17667, A2 => n14670, B1 => n17664, B2 => 
                           n15318, ZN => n14191);
   U5379 : AOI221_X1 port map( B1 => registers_37_31_port, B2 => n17817, C1 => 
                           registers_0_31_port, C2 => n17814, A => n14084, ZN 
                           => n14083);
   U5380 : OAI22_X1 port map( A1 => n17811, A2 => n15691, B1 => n17808, B2 => 
                           n14756, ZN => n14084);
   U5381 : AOI221_X1 port map( B1 => registers_45_24_port, B2 => n16303, C1 => 
                           registers_4_24_port, C2 => n16300, A => n12920, ZN 
                           => n12917);
   U5382 : OAI22_X1 port map( A1 => n16297, A2 => n11907, B1 => n16294, B2 => 
                           n14875, ZN => n12920);
   U5383 : AOI221_X1 port map( B1 => registers_5_24_port, B2 => n16252, C1 => 
                           registers_59_24_port, C2 => n16249, A => n12928, ZN 
                           => n12925);
   U5384 : OAI22_X1 port map( A1 => n16246, A2 => n12342, B1 => n16243, B2 => 
                           n14876, ZN => n12928);
   U5385 : AOI221_X1 port map( B1 => registers_45_25_port, B2 => n16303, C1 => 
                           registers_4_25_port, C2 => n16300, A => n12878, ZN 
                           => n12875);
   U5386 : OAI22_X1 port map( A1 => n16297, A2 => n11945, B1 => n16294, B2 => 
                           n14877, ZN => n12878);
   U5387 : AOI221_X1 port map( B1 => registers_5_25_port, B2 => n16252, C1 => 
                           registers_59_25_port, C2 => n16249, A => n12886, ZN 
                           => n12883);
   U5388 : OAI22_X1 port map( A1 => n16246, A2 => n12343, B1 => n16243, B2 => 
                           n14878, ZN => n12886);
   U5389 : AOI221_X1 port map( B1 => registers_45_26_port, B2 => n16303, C1 => 
                           registers_4_26_port, C2 => n16300, A => n12836, ZN 
                           => n12833);
   U5390 : OAI22_X1 port map( A1 => n16297, A2 => n11946, B1 => n16294, B2 => 
                           n14879, ZN => n12836);
   U5391 : AOI221_X1 port map( B1 => registers_5_26_port, B2 => n16252, C1 => 
                           registers_59_26_port, C2 => n16249, A => n12844, ZN 
                           => n12841);
   U5392 : OAI22_X1 port map( A1 => n16246, A2 => n12344, B1 => n16243, B2 => 
                           n14880, ZN => n12844);
   U5393 : AOI221_X1 port map( B1 => registers_45_27_port, B2 => n16303, C1 => 
                           registers_4_27_port, C2 => n16300, A => n12794, ZN 
                           => n12791);
   U5394 : OAI22_X1 port map( A1 => n16297, A2 => n11947, B1 => n16294, B2 => 
                           n14881, ZN => n12794);
   U5395 : AOI221_X1 port map( B1 => registers_5_27_port, B2 => n16252, C1 => 
                           registers_59_27_port, C2 => n16249, A => n12802, ZN 
                           => n12799);
   U5396 : OAI22_X1 port map( A1 => n16246, A2 => n12345, B1 => n16243, B2 => 
                           n14882, ZN => n12802);
   U5397 : AOI221_X1 port map( B1 => registers_45_28_port, B2 => n16303, C1 => 
                           registers_4_28_port, C2 => n16300, A => n12752, ZN 
                           => n12749);
   U5398 : OAI22_X1 port map( A1 => n16297, A2 => n11948, B1 => n16294, B2 => 
                           n14883, ZN => n12752);
   U5399 : AOI221_X1 port map( B1 => registers_5_28_port, B2 => n16252, C1 => 
                           registers_59_28_port, C2 => n16249, A => n12760, ZN 
                           => n12757);
   U5400 : OAI22_X1 port map( A1 => n16246, A2 => n12346, B1 => n16243, B2 => 
                           n14884, ZN => n12760);
   U5401 : AOI221_X1 port map( B1 => registers_45_29_port, B2 => n16303, C1 => 
                           registers_4_29_port, C2 => n16300, A => n12710, ZN 
                           => n12707);
   U5402 : OAI22_X1 port map( A1 => n16297, A2 => n11949, B1 => n16294, B2 => 
                           n14885, ZN => n12710);
   U5403 : AOI221_X1 port map( B1 => registers_5_29_port, B2 => n16252, C1 => 
                           registers_59_29_port, C2 => n16249, A => n12718, ZN 
                           => n12715);
   U5404 : OAI22_X1 port map( A1 => n16246, A2 => n12347, B1 => n16243, B2 => 
                           n14886, ZN => n12718);
   U5405 : AOI221_X1 port map( B1 => registers_45_30_port, B2 => n16303, C1 => 
                           registers_4_30_port, C2 => n16300, A => n12667, ZN 
                           => n12664);
   U5406 : OAI22_X1 port map( A1 => n16297, A2 => n11670, B1 => n16294, B2 => 
                           n14854, ZN => n12667);
   U5407 : AOI221_X1 port map( B1 => registers_5_30_port, B2 => n16252, C1 => 
                           registers_59_30_port, C2 => n16249, A => n12676, ZN 
                           => n12673);
   U5408 : OAI22_X1 port map( A1 => n16246, A2 => n12196, B1 => n16243, B2 => 
                           n14858, ZN => n12676);
   U5409 : AOI221_X1 port map( B1 => registers_45_31_port, B2 => n16303, C1 => 
                           registers_4_31_port, C2 => n16300, A => n12593, ZN 
                           => n12584);
   U5410 : OAI22_X1 port map( A1 => n16297, A2 => n11950, B1 => n16294, B2 => 
                           n14887, ZN => n12593);
   U5411 : AOI221_X1 port map( B1 => registers_5_31_port, B2 => n16252, C1 => 
                           registers_59_31_port, C2 => n16249, A => n12620, ZN 
                           => n12610);
   U5412 : OAI22_X1 port map( A1 => n16246, A2 => n12348, B1 => n16243, B2 => 
                           n14859, ZN => n12620);
   U5413 : AOI221_X1 port map( B1 => registers_45_24_port, B2 => n16555, C1 => 
                           registers_48_24_port, C2 => n16552, A => n10970, ZN 
                           => n10967);
   U5414 : OAI22_X1 port map( A1 => n16549, A2 => n11907, B1 => n16546, B2 => 
                           n14875, ZN => n10970);
   U5415 : AOI221_X1 port map( B1 => registers_5_24_port, B2 => n16504, C1 => 
                           registers_59_24_port, C2 => n16501, A => n10978, ZN 
                           => n10975);
   U5416 : OAI22_X1 port map( A1 => n16498, A2 => n12342, B1 => n16495, B2 => 
                           n14876, ZN => n10978);
   U5417 : AOI221_X1 port map( B1 => registers_45_25_port, B2 => n16555, C1 => 
                           registers_48_25_port, C2 => n16552, A => n10927, ZN 
                           => n10924);
   U5418 : OAI22_X1 port map( A1 => n16549, A2 => n11945, B1 => n16546, B2 => 
                           n14877, ZN => n10927);
   U5419 : AOI221_X1 port map( B1 => registers_5_25_port, B2 => n16504, C1 => 
                           registers_59_25_port, C2 => n16501, A => n10935, ZN 
                           => n10932);
   U5420 : OAI22_X1 port map( A1 => n16498, A2 => n12343, B1 => n16495, B2 => 
                           n14878, ZN => n10935);
   U5421 : AOI221_X1 port map( B1 => registers_45_26_port, B2 => n16555, C1 => 
                           registers_48_26_port, C2 => n16552, A => n10884, ZN 
                           => n10881);
   U5422 : OAI22_X1 port map( A1 => n16549, A2 => n11946, B1 => n16546, B2 => 
                           n14879, ZN => n10884);
   U5423 : AOI221_X1 port map( B1 => registers_5_26_port, B2 => n16504, C1 => 
                           registers_59_26_port, C2 => n16501, A => n10892, ZN 
                           => n10889);
   U5424 : OAI22_X1 port map( A1 => n16498, A2 => n12344, B1 => n16495, B2 => 
                           n14880, ZN => n10892);
   U5425 : AOI221_X1 port map( B1 => registers_45_27_port, B2 => n16555, C1 => 
                           registers_48_27_port, C2 => n16552, A => n10841, ZN 
                           => n10838);
   U5426 : OAI22_X1 port map( A1 => n16549, A2 => n11947, B1 => n16546, B2 => 
                           n14881, ZN => n10841);
   U5427 : AOI221_X1 port map( B1 => registers_5_27_port, B2 => n16504, C1 => 
                           registers_59_27_port, C2 => n16501, A => n10849, ZN 
                           => n10846);
   U5428 : OAI22_X1 port map( A1 => n16498, A2 => n12345, B1 => n16495, B2 => 
                           n14882, ZN => n10849);
   U5429 : AOI221_X1 port map( B1 => registers_45_28_port, B2 => n16555, C1 => 
                           registers_48_28_port, C2 => n16552, A => n10798, ZN 
                           => n10795);
   U5430 : OAI22_X1 port map( A1 => n16549, A2 => n11948, B1 => n16546, B2 => 
                           n14883, ZN => n10798);
   U5431 : AOI221_X1 port map( B1 => registers_5_28_port, B2 => n16504, C1 => 
                           registers_59_28_port, C2 => n16501, A => n10806, ZN 
                           => n10803);
   U5432 : OAI22_X1 port map( A1 => n16498, A2 => n12346, B1 => n16495, B2 => 
                           n14884, ZN => n10806);
   U5433 : AOI221_X1 port map( B1 => registers_45_29_port, B2 => n16555, C1 => 
                           registers_48_29_port, C2 => n16552, A => n10755, ZN 
                           => n10752);
   U5434 : OAI22_X1 port map( A1 => n16549, A2 => n11949, B1 => n16546, B2 => 
                           n14885, ZN => n10755);
   U5435 : AOI221_X1 port map( B1 => registers_5_29_port, B2 => n16504, C1 => 
                           registers_59_29_port, C2 => n16501, A => n10763, ZN 
                           => n10760);
   U5436 : OAI22_X1 port map( A1 => n16498, A2 => n12347, B1 => n16495, B2 => 
                           n14886, ZN => n10763);
   U5437 : AOI221_X1 port map( B1 => registers_45_30_port, B2 => n16555, C1 => 
                           registers_48_30_port, C2 => n16552, A => n10707, ZN 
                           => n10702);
   U5438 : OAI22_X1 port map( A1 => n16549, A2 => n11670, B1 => n16546, B2 => 
                           n14854, ZN => n10707);
   U5439 : AOI221_X1 port map( B1 => registers_5_30_port, B2 => n16504, C1 => 
                           registers_59_30_port, C2 => n16501, A => n10718, ZN 
                           => n10715);
   U5440 : OAI22_X1 port map( A1 => n16498, A2 => n12196, B1 => n16495, B2 => 
                           n14858, ZN => n10718);
   U5441 : AOI221_X1 port map( B1 => registers_45_31_port, B2 => n16555, C1 => 
                           registers_48_31_port, C2 => n16552, A => n10609, ZN 
                           => n10598);
   U5442 : OAI22_X1 port map( A1 => n16549, A2 => n11950, B1 => n16546, B2 => 
                           n14887, ZN => n10609);
   U5443 : AOI221_X1 port map( B1 => registers_5_31_port, B2 => n16504, C1 => 
                           registers_59_31_port, C2 => n16501, A => n10643, ZN 
                           => n10630);
   U5444 : OAI22_X1 port map( A1 => n16498, A2 => n12348, B1 => n16495, B2 => 
                           n14859, ZN => n10643);
   U5445 : AOI221_X1 port map( B1 => registers_63_23_port, B2 => n17663, C1 => 
                           registers_62_23_port, C2 => n17660, A => n5315, ZN 
                           => n5312);
   U5446 : OAI22_X1 port map( A1 => n17657, A2 => n14050, B1 => n17654, B2 => 
                           n15319, ZN => n5315);
   U5447 : AOI221_X1 port map( B1 => registers_11_23_port, B2 => n17807, C1 => 
                           net227324, C2 => n17804, A => n5282, ZN => n5279);
   U5448 : OAI22_X1 port map( A1 => n17801, A2 => n15692, B1 => n17798, B2 => 
                           n11874, ZN => n5282);
   U5449 : AOI221_X1 port map( B1 => registers_63_24_port, B2 => n17663, C1 => 
                           registers_62_24_port, C2 => n17660, A => n5143, ZN 
                           => n5140);
   U5450 : OAI22_X1 port map( A1 => n17657, A2 => n12342, B1 => n17654, B2 => 
                           n15320, ZN => n5143);
   U5451 : AOI221_X1 port map( B1 => registers_11_24_port, B2 => n17807, C1 => 
                           net227342, C2 => n17804, A => n5117, ZN => n5113);
   U5452 : OAI22_X1 port map( A1 => n17801, A2 => n15693, B1 => n17798, B2 => 
                           n11875, ZN => n5117);
   U5453 : AOI221_X1 port map( B1 => registers_63_25_port, B2 => n17663, C1 => 
                           registers_62_25_port, C2 => n17660, A => n5029, ZN 
                           => n5026);
   U5454 : OAI22_X1 port map( A1 => n17657, A2 => n12343, B1 => n17654, B2 => 
                           n15321, ZN => n5029);
   U5455 : AOI221_X1 port map( B1 => registers_11_25_port, B2 => n17807, C1 => 
                           net227360, C2 => n17804, A => n5003, ZN => n5000);
   U5456 : OAI22_X1 port map( A1 => n17801, A2 => n15694, B1 => n17798, B2 => 
                           n11876, ZN => n5003);
   U5457 : AOI221_X1 port map( B1 => registers_63_26_port, B2 => n17663, C1 => 
                           registers_62_26_port, C2 => n17660, A => n4911, ZN 
                           => n4908);
   U5458 : OAI22_X1 port map( A1 => n17657, A2 => n12344, B1 => n17654, B2 => 
                           n15322, ZN => n4911);
   U5459 : AOI221_X1 port map( B1 => registers_11_26_port, B2 => n17807, C1 => 
                           net227378, C2 => n17804, A => n4881, ZN => n4878);
   U5460 : OAI22_X1 port map( A1 => n17801, A2 => n15695, B1 => n17798, B2 => 
                           n11877, ZN => n4881);
   U5461 : AOI221_X1 port map( B1 => registers_63_27_port, B2 => n17663, C1 => 
                           registers_62_27_port, C2 => n17660, A => n4780, ZN 
                           => n4777);
   U5462 : OAI22_X1 port map( A1 => n17657, A2 => n12345, B1 => n17654, B2 => 
                           n15323, ZN => n4780);
   U5463 : AOI221_X1 port map( B1 => registers_11_27_port, B2 => n17807, C1 => 
                           net227396, C2 => n17804, A => n4752, ZN => n4749);
   U5464 : OAI22_X1 port map( A1 => n17801, A2 => n15696, B1 => n17798, B2 => 
                           n11878, ZN => n4752);
   U5465 : AOI221_X1 port map( B1 => registers_63_28_port, B2 => n17663, C1 => 
                           registers_62_28_port, C2 => n17660, A => n4651, ZN 
                           => n4648);
   U5466 : OAI22_X1 port map( A1 => n17657, A2 => n12346, B1 => n17654, B2 => 
                           n15324, ZN => n4651);
   U5467 : AOI221_X1 port map( B1 => registers_11_28_port, B2 => n17807, C1 => 
                           net227414, C2 => n17804, A => n4623, ZN => n4620);
   U5468 : OAI22_X1 port map( A1 => n17801, A2 => n15697, B1 => n17798, B2 => 
                           n11879, ZN => n4623);
   U5469 : AOI221_X1 port map( B1 => registers_63_29_port, B2 => n17663, C1 => 
                           registers_62_29_port, C2 => n17660, A => n4522, ZN 
                           => n4519);
   U5470 : OAI22_X1 port map( A1 => n17657, A2 => n12347, B1 => n17654, B2 => 
                           n15325, ZN => n4522);
   U5471 : AOI221_X1 port map( B1 => registers_11_29_port, B2 => n17807, C1 => 
                           net227432, C2 => n17804, A => n4490, ZN => n4487);
   U5472 : OAI22_X1 port map( A1 => n17801, A2 => n15698, B1 => n17798, B2 => 
                           n11880, ZN => n4490);
   U5473 : AOI221_X1 port map( B1 => registers_63_30_port, B2 => n17663, C1 => 
                           registers_62_30_port, C2 => n17660, A => n4227, ZN 
                           => n4217);
   U5474 : OAI22_X1 port map( A1 => n17657, A2 => n12196, B1 => n17654, B2 => 
                           n15271, ZN => n4227);
   U5475 : AOI221_X1 port map( B1 => registers_11_30_port, B2 => n17807, C1 => 
                           net227450, C2 => n17804, A => n4118, ZN => n4103);
   U5476 : OAI22_X1 port map( A1 => n17801, A2 => n15281, B1 => n17798, B2 => 
                           n11541, ZN => n4118);
   U5477 : AOI221_X1 port map( B1 => registers_45_0_port, B2 => n16301, C1 => 
                           registers_4_0_port, C2 => n16298, A => n13954, ZN =>
                           n13950);
   U5478 : OAI22_X1 port map( A1 => n16295, A2 => n11951, B1 => n16292, B2 => 
                           n14888, ZN => n13954);
   U5479 : AOI221_X1 port map( B1 => registers_45_1_port, B2 => n16301, C1 => 
                           registers_4_1_port, C2 => n16298, A => n13886, ZN =>
                           n13883);
   U5480 : OAI22_X1 port map( A1 => n16295, A2 => n11952, B1 => n16292, B2 => 
                           n14889, ZN => n13886);
   U5481 : AOI221_X1 port map( B1 => registers_45_2_port, B2 => n16301, C1 => 
                           registers_4_2_port, C2 => n16298, A => n13844, ZN =>
                           n13841);
   U5482 : OAI22_X1 port map( A1 => n16295, A2 => n11995, B1 => n16292, B2 => 
                           n14890, ZN => n13844);
   U5483 : AOI221_X1 port map( B1 => registers_45_3_port, B2 => n16301, C1 => 
                           registers_4_3_port, C2 => n16298, A => n13802, ZN =>
                           n13799);
   U5484 : OAI22_X1 port map( A1 => n16295, A2 => n11905, B1 => n16292, B2 => 
                           n14861, ZN => n13802);
   U5485 : AOI221_X1 port map( B1 => registers_45_4_port, B2 => n16301, C1 => 
                           registers_4_4_port, C2 => n16298, A => n13760, ZN =>
                           n13757);
   U5486 : OAI22_X1 port map( A1 => n16295, A2 => n11997, B1 => n16292, B2 => 
                           n14891, ZN => n13760);
   U5487 : AOI221_X1 port map( B1 => registers_45_5_port, B2 => n16301, C1 => 
                           registers_4_5_port, C2 => n16298, A => n13718, ZN =>
                           n13715);
   U5488 : OAI22_X1 port map( A1 => n16295, A2 => n11906, B1 => n16292, B2 => 
                           n14862, ZN => n13718);
   U5489 : AOI221_X1 port map( B1 => registers_45_6_port, B2 => n16301, C1 => 
                           registers_4_6_port, C2 => n16298, A => n13676, ZN =>
                           n13673);
   U5490 : OAI22_X1 port map( A1 => n16295, A2 => n11998, B1 => n16292, B2 => 
                           n14892, ZN => n13676);
   U5491 : AOI221_X1 port map( B1 => registers_45_7_port, B2 => n16301, C1 => 
                           registers_4_7_port, C2 => n16298, A => n13634, ZN =>
                           n13631);
   U5492 : OAI22_X1 port map( A1 => n16295, A2 => n11999, B1 => n16292, B2 => 
                           n14893, ZN => n13634);
   U5493 : AOI221_X1 port map( B1 => registers_45_8_port, B2 => n16301, C1 => 
                           registers_4_8_port, C2 => n16298, A => n13592, ZN =>
                           n13589);
   U5494 : OAI22_X1 port map( A1 => n16295, A2 => n12000, B1 => n16292, B2 => 
                           n14894, ZN => n13592);
   U5495 : AOI221_X1 port map( B1 => registers_45_9_port, B2 => n16301, C1 => 
                           registers_4_9_port, C2 => n16298, A => n13550, ZN =>
                           n13547);
   U5496 : OAI22_X1 port map( A1 => n16295, A2 => n12001, B1 => n16292, B2 => 
                           n14895, ZN => n13550);
   U5497 : AOI221_X1 port map( B1 => registers_45_10_port, B2 => n16301, C1 => 
                           registers_4_10_port, C2 => n16298, A => n13508, ZN 
                           => n13505);
   U5498 : OAI22_X1 port map( A1 => n16295, A2 => n12002, B1 => n16292, B2 => 
                           n14896, ZN => n13508);
   U5499 : AOI221_X1 port map( B1 => registers_45_11_port, B2 => n16301, C1 => 
                           registers_4_11_port, C2 => n16298, A => n13466, ZN 
                           => n13463);
   U5500 : OAI22_X1 port map( A1 => n16295, A2 => n12003, B1 => n16292, B2 => 
                           n14897, ZN => n13466);
   U5501 : AOI221_X1 port map( B1 => registers_45_12_port, B2 => n16302, C1 => 
                           registers_4_12_port, C2 => n16299, A => n13424, ZN 
                           => n13421);
   U5502 : OAI22_X1 port map( A1 => n16296, A2 => n12004, B1 => n16293, B2 => 
                           n14898, ZN => n13424);
   U5503 : AOI221_X1 port map( B1 => registers_45_13_port, B2 => n16302, C1 => 
                           registers_4_13_port, C2 => n16299, A => n13382, ZN 
                           => n13379);
   U5504 : OAI22_X1 port map( A1 => n16296, A2 => n12005, B1 => n16293, B2 => 
                           n14899, ZN => n13382);
   U5505 : AOI221_X1 port map( B1 => registers_45_14_port, B2 => n16302, C1 => 
                           registers_4_14_port, C2 => n16299, A => n13340, ZN 
                           => n13337);
   U5506 : OAI22_X1 port map( A1 => n16296, A2 => n12006, B1 => n16293, B2 => 
                           n14900, ZN => n13340);
   U5507 : AOI221_X1 port map( B1 => registers_45_15_port, B2 => n16302, C1 => 
                           registers_4_15_port, C2 => n16299, A => n13298, ZN 
                           => n13295);
   U5508 : OAI22_X1 port map( A1 => n16296, A2 => n12007, B1 => n16293, B2 => 
                           n14901, ZN => n13298);
   U5509 : AOI221_X1 port map( B1 => registers_45_16_port, B2 => n16302, C1 => 
                           registers_4_16_port, C2 => n16299, A => n13256, ZN 
                           => n13253);
   U5510 : OAI22_X1 port map( A1 => n16296, A2 => n12008, B1 => n16293, B2 => 
                           n14902, ZN => n13256);
   U5511 : AOI221_X1 port map( B1 => registers_45_17_port, B2 => n16302, C1 => 
                           registers_4_17_port, C2 => n16299, A => n13214, ZN 
                           => n13211);
   U5512 : OAI22_X1 port map( A1 => n16296, A2 => n12009, B1 => n16293, B2 => 
                           n14903, ZN => n13214);
   U5513 : AOI221_X1 port map( B1 => registers_45_18_port, B2 => n16302, C1 => 
                           registers_4_18_port, C2 => n16299, A => n13172, ZN 
                           => n13169);
   U5514 : OAI22_X1 port map( A1 => n16296, A2 => n12010, B1 => n16293, B2 => 
                           n14904, ZN => n13172);
   U5515 : AOI221_X1 port map( B1 => registers_45_19_port, B2 => n16302, C1 => 
                           registers_4_19_port, C2 => n16299, A => n13130, ZN 
                           => n13127);
   U5516 : OAI22_X1 port map( A1 => n16296, A2 => n12011, B1 => n16293, B2 => 
                           n14905, ZN => n13130);
   U5517 : AOI221_X1 port map( B1 => registers_45_20_port, B2 => n16302, C1 => 
                           registers_4_20_port, C2 => n16299, A => n13088, ZN 
                           => n13085);
   U5518 : OAI22_X1 port map( A1 => n16296, A2 => n12012, B1 => n16293, B2 => 
                           n14906, ZN => n13088);
   U5519 : AOI221_X1 port map( B1 => registers_45_21_port, B2 => n16302, C1 => 
                           registers_4_21_port, C2 => n16299, A => n13046, ZN 
                           => n13043);
   U5520 : OAI22_X1 port map( A1 => n16296, A2 => n12013, B1 => n16293, B2 => 
                           n14907, ZN => n13046);
   U5521 : AOI221_X1 port map( B1 => registers_45_22_port, B2 => n16302, C1 => 
                           registers_4_22_port, C2 => n16299, A => n13004, ZN 
                           => n13001);
   U5522 : OAI22_X1 port map( A1 => n16296, A2 => n12014, B1 => n16293, B2 => 
                           n14908, ZN => n13004);
   U5523 : AOI221_X1 port map( B1 => registers_45_23_port, B2 => n16302, C1 => 
                           registers_4_23_port, C2 => n16299, A => n12962, ZN 
                           => n12959);
   U5524 : OAI22_X1 port map( A1 => n16296, A2 => n12015, B1 => n16293, B2 => 
                           n14909, ZN => n12962);
   U5525 : AOI221_X1 port map( B1 => registers_45_0_port, B2 => n16553, C1 => 
                           registers_48_0_port, C2 => n16550, A => n12473, ZN 
                           => n12469);
   U5526 : OAI22_X1 port map( A1 => n16547, A2 => n11951, B1 => n16544, B2 => 
                           n14888, ZN => n12473);
   U5527 : AOI221_X1 port map( B1 => registers_5_0_port, B2 => n16502, C1 => 
                           registers_59_0_port, C2 => n16499, A => n12490, ZN 
                           => n12485);
   U5528 : OAI22_X1 port map( A1 => n16496, A2 => n12357, B1 => n16493, B2 => 
                           n14910, ZN => n12490);
   U5529 : AOI221_X1 port map( B1 => registers_45_1_port, B2 => n16553, C1 => 
                           registers_48_1_port, C2 => n16550, A => n12290, ZN 
                           => n12287);
   U5530 : OAI22_X1 port map( A1 => n16547, A2 => n11952, B1 => n16544, B2 => 
                           n14889, ZN => n12290);
   U5531 : AOI221_X1 port map( B1 => registers_5_1_port, B2 => n16502, C1 => 
                           registers_59_1_port, C2 => n16499, A => n12298, ZN 
                           => n12295);
   U5532 : OAI22_X1 port map( A1 => n16496, A2 => n12359, B1 => n16493, B2 => 
                           n14911, ZN => n12298);
   U5533 : AOI221_X1 port map( B1 => registers_45_2_port, B2 => n16553, C1 => 
                           registers_48_2_port, C2 => n16550, A => n12137, ZN 
                           => n12134);
   U5534 : OAI22_X1 port map( A1 => n16547, A2 => n11995, B1 => n16544, B2 => 
                           n14890, ZN => n12137);
   U5535 : AOI221_X1 port map( B1 => registers_5_2_port, B2 => n16502, C1 => 
                           registers_59_2_port, C2 => n16499, A => n12145, ZN 
                           => n12142);
   U5536 : OAI22_X1 port map( A1 => n16496, A2 => n12361, B1 => n16493, B2 => 
                           n14912, ZN => n12145);
   U5537 : AOI221_X1 port map( B1 => registers_45_3_port, B2 => n16553, C1 => 
                           registers_48_3_port, C2 => n16550, A => n11984, ZN 
                           => n11981);
   U5538 : OAI22_X1 port map( A1 => n16547, A2 => n11905, B1 => n16544, B2 => 
                           n14861, ZN => n11984);
   U5539 : AOI221_X1 port map( B1 => registers_5_3_port, B2 => n16502, C1 => 
                           registers_59_3_port, C2 => n16499, A => n11992, ZN 
                           => n11989);
   U5540 : OAI22_X1 port map( A1 => n16496, A2 => n12362, B1 => n16493, B2 => 
                           n14863, ZN => n11992);
   U5541 : AOI221_X1 port map( B1 => registers_45_4_port, B2 => n16553, C1 => 
                           registers_48_4_port, C2 => n16550, A => n11831, ZN 
                           => n11828);
   U5542 : OAI22_X1 port map( A1 => n16547, A2 => n11997, B1 => n16544, B2 => 
                           n14891, ZN => n11831);
   U5543 : AOI221_X1 port map( B1 => registers_5_4_port, B2 => n16502, C1 => 
                           registers_59_4_port, C2 => n16499, A => n11839, ZN 
                           => n11836);
   U5544 : OAI22_X1 port map( A1 => n16496, A2 => n12363, B1 => n16493, B2 => 
                           n14864, ZN => n11839);
   U5545 : AOI221_X1 port map( B1 => registers_45_5_port, B2 => n16553, C1 => 
                           registers_48_5_port, C2 => n16550, A => n11788, ZN 
                           => n11785);
   U5546 : OAI22_X1 port map( A1 => n16547, A2 => n11906, B1 => n16544, B2 => 
                           n14862, ZN => n11788);
   U5547 : AOI221_X1 port map( B1 => registers_5_5_port, B2 => n16502, C1 => 
                           registers_59_5_port, C2 => n16499, A => n11796, ZN 
                           => n11793);
   U5548 : OAI22_X1 port map( A1 => n16496, A2 => n12365, B1 => n16493, B2 => 
                           n14865, ZN => n11796);
   U5549 : AOI221_X1 port map( B1 => registers_45_6_port, B2 => n16553, C1 => 
                           registers_48_6_port, C2 => n16550, A => n11745, ZN 
                           => n11742);
   U5550 : OAI22_X1 port map( A1 => n16547, A2 => n11998, B1 => n16544, B2 => 
                           n14892, ZN => n11745);
   U5551 : AOI221_X1 port map( B1 => registers_5_6_port, B2 => n16502, C1 => 
                           registers_59_6_port, C2 => n16499, A => n11753, ZN 
                           => n11750);
   U5552 : OAI22_X1 port map( A1 => n16496, A2 => n12367, B1 => n16493, B2 => 
                           n14913, ZN => n11753);
   U5553 : AOI221_X1 port map( B1 => registers_45_7_port, B2 => n16553, C1 => 
                           registers_48_7_port, C2 => n16550, A => n11702, ZN 
                           => n11699);
   U5554 : OAI22_X1 port map( A1 => n16547, A2 => n11999, B1 => n16544, B2 => 
                           n14893, ZN => n11702);
   U5555 : AOI221_X1 port map( B1 => registers_5_7_port, B2 => n16502, C1 => 
                           registers_59_7_port, C2 => n16499, A => n11710, ZN 
                           => n11707);
   U5556 : OAI22_X1 port map( A1 => n16496, A2 => n12369, B1 => n16493, B2 => 
                           n14914, ZN => n11710);
   U5557 : AOI221_X1 port map( B1 => registers_45_8_port, B2 => n16553, C1 => 
                           registers_48_8_port, C2 => n16550, A => n11659, ZN 
                           => n11656);
   U5558 : OAI22_X1 port map( A1 => n16547, A2 => n12000, B1 => n16544, B2 => 
                           n14894, ZN => n11659);
   U5559 : AOI221_X1 port map( B1 => registers_5_8_port, B2 => n16502, C1 => 
                           registers_59_8_port, C2 => n16499, A => n11667, ZN 
                           => n11664);
   U5560 : OAI22_X1 port map( A1 => n16496, A2 => n12408, B1 => n16493, B2 => 
                           n14915, ZN => n11667);
   U5561 : AOI221_X1 port map( B1 => registers_45_9_port, B2 => n16553, C1 => 
                           registers_48_9_port, C2 => n16550, A => n11616, ZN 
                           => n11613);
   U5562 : OAI22_X1 port map( A1 => n16547, A2 => n12001, B1 => n16544, B2 => 
                           n14895, ZN => n11616);
   U5563 : AOI221_X1 port map( B1 => registers_5_9_port, B2 => n16502, C1 => 
                           registers_59_9_port, C2 => n16499, A => n11624, ZN 
                           => n11621);
   U5564 : OAI22_X1 port map( A1 => n16496, A2 => n12410, B1 => n16493, B2 => 
                           n14916, ZN => n11624);
   U5565 : AOI221_X1 port map( B1 => registers_45_10_port, B2 => n16553, C1 => 
                           registers_48_10_port, C2 => n16550, A => n11573, ZN 
                           => n11570);
   U5566 : OAI22_X1 port map( A1 => n16547, A2 => n12002, B1 => n16544, B2 => 
                           n14896, ZN => n11573);
   U5567 : AOI221_X1 port map( B1 => registers_5_10_port, B2 => n16502, C1 => 
                           registers_59_10_port, C2 => n16499, A => n11581, ZN 
                           => n11578);
   U5568 : OAI22_X1 port map( A1 => n16496, A2 => n12551, B1 => n16493, B2 => 
                           n14917, ZN => n11581);
   U5569 : AOI221_X1 port map( B1 => registers_45_11_port, B2 => n16553, C1 => 
                           registers_48_11_port, C2 => n16550, A => n11530, ZN 
                           => n11527);
   U5570 : OAI22_X1 port map( A1 => n16547, A2 => n12003, B1 => n16544, B2 => 
                           n14897, ZN => n11530);
   U5571 : AOI221_X1 port map( B1 => registers_5_11_port, B2 => n16502, C1 => 
                           registers_59_11_port, C2 => n16499, A => n11538, ZN 
                           => n11535);
   U5572 : OAI22_X1 port map( A1 => n16496, A2 => n12602, B1 => n16493, B2 => 
                           n14918, ZN => n11538);
   U5573 : AOI221_X1 port map( B1 => registers_45_12_port, B2 => n16554, C1 => 
                           registers_48_12_port, C2 => n16551, A => n11487, ZN 
                           => n11484);
   U5574 : OAI22_X1 port map( A1 => n16548, A2 => n12004, B1 => n16545, B2 => 
                           n14898, ZN => n11487);
   U5575 : AOI221_X1 port map( B1 => registers_5_12_port, B2 => n16503, C1 => 
                           registers_59_12_port, C2 => n16500, A => n11495, ZN 
                           => n11492);
   U5576 : OAI22_X1 port map( A1 => n16497, A2 => n12669, B1 => n16494, B2 => 
                           n14919, ZN => n11495);
   U5577 : AOI221_X1 port map( B1 => registers_45_13_port, B2 => n16554, C1 => 
                           registers_48_13_port, C2 => n16551, A => n11443, ZN 
                           => n11440);
   U5578 : OAI22_X1 port map( A1 => n16548, A2 => n12005, B1 => n16545, B2 => 
                           n14899, ZN => n11443);
   U5579 : AOI221_X1 port map( B1 => registers_5_13_port, B2 => n16503, C1 => 
                           registers_59_13_port, C2 => n16500, A => n11451, ZN 
                           => n11448);
   U5580 : OAI22_X1 port map( A1 => n16497, A2 => n13999, B1 => n16494, B2 => 
                           n14920, ZN => n11451);
   U5581 : AOI221_X1 port map( B1 => registers_45_14_port, B2 => n16554, C1 => 
                           registers_48_14_port, C2 => n16551, A => n11400, ZN 
                           => n11397);
   U5582 : OAI22_X1 port map( A1 => n16548, A2 => n12006, B1 => n16545, B2 => 
                           n14900, ZN => n11400);
   U5583 : AOI221_X1 port map( B1 => registers_5_14_port, B2 => n16503, C1 => 
                           registers_59_14_port, C2 => n16500, A => n11408, ZN 
                           => n11405);
   U5584 : OAI22_X1 port map( A1 => n16497, A2 => n14014, B1 => n16494, B2 => 
                           n14921, ZN => n11408);
   U5585 : AOI221_X1 port map( B1 => registers_45_15_port, B2 => n16554, C1 => 
                           registers_48_15_port, C2 => n16551, A => n11357, ZN 
                           => n11354);
   U5586 : OAI22_X1 port map( A1 => n16548, A2 => n12007, B1 => n16545, B2 => 
                           n14901, ZN => n11357);
   U5587 : AOI221_X1 port map( B1 => registers_5_15_port, B2 => n16503, C1 => 
                           registers_59_15_port, C2 => n16500, A => n11365, ZN 
                           => n11362);
   U5588 : OAI22_X1 port map( A1 => n16497, A2 => n14032, B1 => n16494, B2 => 
                           n14922, ZN => n11365);
   U5589 : AOI221_X1 port map( B1 => registers_45_16_port, B2 => n16554, C1 => 
                           registers_48_16_port, C2 => n16551, A => n11314, ZN 
                           => n11311);
   U5590 : OAI22_X1 port map( A1 => n16548, A2 => n12008, B1 => n16545, B2 => 
                           n14902, ZN => n11314);
   U5591 : AOI221_X1 port map( B1 => registers_5_16_port, B2 => n16503, C1 => 
                           registers_59_16_port, C2 => n16500, A => n11322, ZN 
                           => n11319);
   U5592 : OAI22_X1 port map( A1 => n16497, A2 => n14036, B1 => n16494, B2 => 
                           n14923, ZN => n11322);
   U5593 : AOI221_X1 port map( B1 => registers_45_17_port, B2 => n16554, C1 => 
                           registers_48_17_port, C2 => n16551, A => n11271, ZN 
                           => n11268);
   U5594 : OAI22_X1 port map( A1 => n16548, A2 => n12009, B1 => n16545, B2 => 
                           n14903, ZN => n11271);
   U5595 : AOI221_X1 port map( B1 => registers_5_17_port, B2 => n16503, C1 => 
                           registers_59_17_port, C2 => n16500, A => n11279, ZN 
                           => n11276);
   U5596 : OAI22_X1 port map( A1 => n16497, A2 => n14038, B1 => n16494, B2 => 
                           n14924, ZN => n11279);
   U5597 : AOI221_X1 port map( B1 => registers_45_18_port, B2 => n16554, C1 => 
                           registers_48_18_port, C2 => n16551, A => n11228, ZN 
                           => n11225);
   U5598 : OAI22_X1 port map( A1 => n16548, A2 => n12010, B1 => n16545, B2 => 
                           n14904, ZN => n11228);
   U5599 : AOI221_X1 port map( B1 => registers_5_18_port, B2 => n16503, C1 => 
                           registers_59_18_port, C2 => n16500, A => n11236, ZN 
                           => n11233);
   U5600 : OAI22_X1 port map( A1 => n16497, A2 => n14040, B1 => n16494, B2 => 
                           n14925, ZN => n11236);
   U5601 : AOI221_X1 port map( B1 => registers_45_19_port, B2 => n16554, C1 => 
                           registers_48_19_port, C2 => n16551, A => n11185, ZN 
                           => n11182);
   U5602 : OAI22_X1 port map( A1 => n16548, A2 => n12011, B1 => n16545, B2 => 
                           n14905, ZN => n11185);
   U5603 : AOI221_X1 port map( B1 => registers_5_19_port, B2 => n16503, C1 => 
                           registers_59_19_port, C2 => n16500, A => n11193, ZN 
                           => n11190);
   U5604 : OAI22_X1 port map( A1 => n16497, A2 => n14042, B1 => n16494, B2 => 
                           n14926, ZN => n11193);
   U5605 : AOI221_X1 port map( B1 => registers_45_20_port, B2 => n16554, C1 => 
                           registers_48_20_port, C2 => n16551, A => n11142, ZN 
                           => n11139);
   U5606 : OAI22_X1 port map( A1 => n16548, A2 => n12012, B1 => n16545, B2 => 
                           n14906, ZN => n11142);
   U5607 : AOI221_X1 port map( B1 => registers_5_20_port, B2 => n16503, C1 => 
                           registers_59_20_port, C2 => n16500, A => n11150, ZN 
                           => n11147);
   U5608 : OAI22_X1 port map( A1 => n16497, A2 => n14044, B1 => n16494, B2 => 
                           n14927, ZN => n11150);
   U5609 : AOI221_X1 port map( B1 => registers_45_21_port, B2 => n16554, C1 => 
                           registers_48_21_port, C2 => n16551, A => n11099, ZN 
                           => n11096);
   U5610 : OAI22_X1 port map( A1 => n16548, A2 => n12013, B1 => n16545, B2 => 
                           n14907, ZN => n11099);
   U5611 : AOI221_X1 port map( B1 => registers_5_21_port, B2 => n16503, C1 => 
                           registers_59_21_port, C2 => n16500, A => n11107, ZN 
                           => n11104);
   U5612 : OAI22_X1 port map( A1 => n16497, A2 => n14046, B1 => n16494, B2 => 
                           n14928, ZN => n11107);
   U5613 : AOI221_X1 port map( B1 => registers_45_22_port, B2 => n16554, C1 => 
                           registers_48_22_port, C2 => n16551, A => n11056, ZN 
                           => n11053);
   U5614 : OAI22_X1 port map( A1 => n16548, A2 => n12014, B1 => n16545, B2 => 
                           n14908, ZN => n11056);
   U5615 : AOI221_X1 port map( B1 => registers_5_22_port, B2 => n16503, C1 => 
                           registers_59_22_port, C2 => n16500, A => n11064, ZN 
                           => n11061);
   U5616 : OAI22_X1 port map( A1 => n16497, A2 => n14048, B1 => n16494, B2 => 
                           n14929, ZN => n11064);
   U5617 : AOI221_X1 port map( B1 => registers_45_23_port, B2 => n16554, C1 => 
                           registers_48_23_port, C2 => n16551, A => n11013, ZN 
                           => n11010);
   U5618 : OAI22_X1 port map( A1 => n16548, A2 => n12015, B1 => n16545, B2 => 
                           n14909, ZN => n11013);
   U5619 : AOI221_X1 port map( B1 => registers_5_23_port, B2 => n16503, C1 => 
                           registers_59_23_port, C2 => n16500, A => n11021, ZN 
                           => n11018);
   U5620 : OAI22_X1 port map( A1 => n16497, A2 => n14050, B1 => n16494, B2 => 
                           n14930, ZN => n11021);
   U5621 : AOI221_X1 port map( B1 => registers_63_0_port, B2 => n17661, C1 => 
                           registers_62_0_port, C2 => n17658, A => n12404, ZN 
                           => n12401);
   U5622 : OAI22_X1 port map( A1 => n17655, A2 => n12357, B1 => n17652, B2 => 
                           n15326, ZN => n12404);
   U5623 : AOI221_X1 port map( B1 => registers_11_0_port, B2 => n17805, C1 => 
                           net226849, C2 => n17802, A => n12380, ZN => n12377);
   U5624 : OAI22_X1 port map( A1 => n17799, A2 => n15699, B1 => n17796, B2 => 
                           n11881, ZN => n12380);
   U5625 : AOI221_X1 port map( B1 => registers_63_1_port, B2 => n17661, C1 => 
                           registers_62_1_port, C2 => n17658, A => n12250, ZN 
                           => n12247);
   U5626 : OAI22_X1 port map( A1 => n17655, A2 => n12359, B1 => n17652, B2 => 
                           n15327, ZN => n12250);
   U5627 : AOI221_X1 port map( B1 => registers_11_1_port, B2 => n17805, C1 => 
                           net226863, C2 => n17802, A => n12226, ZN => n12223);
   U5628 : OAI22_X1 port map( A1 => n17799, A2 => n15700, B1 => n17796, B2 => 
                           n11882, ZN => n12226);
   U5629 : AOI221_X1 port map( B1 => registers_63_2_port, B2 => n17661, C1 => 
                           registers_62_2_port, C2 => n17658, A => n12095, ZN 
                           => n12092);
   U5630 : OAI22_X1 port map( A1 => n17655, A2 => n12361, B1 => n17652, B2 => 
                           n15328, ZN => n12095);
   U5631 : AOI221_X1 port map( B1 => registers_11_2_port, B2 => n17805, C1 => 
                           net226890, C2 => n17802, A => n12071, ZN => n12068);
   U5632 : OAI22_X1 port map( A1 => n17799, A2 => n15701, B1 => n17796, B2 => 
                           n11883, ZN => n12071);
   U5633 : AOI221_X1 port map( B1 => registers_63_3_port, B2 => n17661, C1 => 
                           registers_62_3_port, C2 => n17658, A => n11942, ZN 
                           => n11939);
   U5634 : OAI22_X1 port map( A1 => n17655, A2 => n12362, B1 => n17652, B2 => 
                           n15329, ZN => n11942);
   U5635 : AOI221_X1 port map( B1 => registers_11_3_port, B2 => n17805, C1 => 
                           net226901, C2 => n17802, A => n11918, ZN => n11915);
   U5636 : OAI22_X1 port map( A1 => n17799, A2 => n15702, B1 => n17796, B2 => 
                           n11627, ZN => n11918);
   U5637 : AOI221_X1 port map( B1 => registers_63_4_port, B2 => n17661, C1 => 
                           registers_62_4_port, C2 => n17658, A => n10499, ZN 
                           => n10496);
   U5638 : OAI22_X1 port map( A1 => n17655, A2 => n12363, B1 => n17652, B2 => 
                           n15330, ZN => n10499);
   U5639 : AOI221_X1 port map( B1 => registers_11_4_port, B2 => n17805, C1 => 
                           net226974, C2 => n17802, A => n10475, ZN => n10472);
   U5640 : OAI22_X1 port map( A1 => n17799, A2 => n15366, B1 => n17796, B2 => 
                           n11884, ZN => n10475);
   U5641 : AOI221_X1 port map( B1 => registers_63_5_port, B2 => n17661, C1 => 
                           registers_62_5_port, C2 => n17658, A => n10389, ZN 
                           => n10386);
   U5642 : OAI22_X1 port map( A1 => n17655, A2 => n12365, B1 => n17652, B2 => 
                           n15331, ZN => n10389);
   U5643 : AOI221_X1 port map( B1 => registers_11_5_port, B2 => n17805, C1 => 
                           net226994, C2 => n17802, A => n10365, ZN => n10362);
   U5644 : OAI22_X1 port map( A1 => n17799, A2 => n15703, B1 => n17796, B2 => 
                           n11885, ZN => n10365);
   U5645 : AOI221_X1 port map( B1 => registers_63_6_port, B2 => n17661, C1 => 
                           registers_62_6_port, C2 => n17658, A => n10277, ZN 
                           => n10274);
   U5646 : OAI22_X1 port map( A1 => n17655, A2 => n12367, B1 => n17652, B2 => 
                           n15332, ZN => n10277);
   U5647 : AOI221_X1 port map( B1 => registers_11_6_port, B2 => n17805, C1 => 
                           net227018, C2 => n17802, A => n10253, ZN => n10250);
   U5648 : OAI22_X1 port map( A1 => n17799, A2 => n15704, B1 => n17796, B2 => 
                           n11886, ZN => n10253);
   U5649 : AOI221_X1 port map( B1 => registers_63_7_port, B2 => n17661, C1 => 
                           registers_62_7_port, C2 => n17658, A => n7641, ZN =>
                           n7638);
   U5650 : OAI22_X1 port map( A1 => n17655, A2 => n12369, B1 => n17652, B2 => 
                           n15333, ZN => n7641);
   U5651 : AOI221_X1 port map( B1 => registers_11_7_port, B2 => n17805, C1 => 
                           net227036, C2 => n17802, A => n7617, ZN => n7614);
   U5652 : OAI22_X1 port map( A1 => n17799, A2 => n15705, B1 => n17796, B2 => 
                           n11887, ZN => n7617);
   U5653 : AOI221_X1 port map( B1 => registers_63_8_port, B2 => n17661, C1 => 
                           registers_62_8_port, C2 => n17658, A => n7526, ZN =>
                           n7523);
   U5654 : OAI22_X1 port map( A1 => n17655, A2 => n12408, B1 => n17652, B2 => 
                           n15334, ZN => n7526);
   U5655 : AOI221_X1 port map( B1 => registers_11_8_port, B2 => n17805, C1 => 
                           net227054, C2 => n17802, A => n7502, ZN => n7499);
   U5656 : OAI22_X1 port map( A1 => n17799, A2 => n15706, B1 => n17796, B2 => 
                           n11888, ZN => n7502);
   U5657 : AOI221_X1 port map( B1 => registers_63_9_port, B2 => n17661, C1 => 
                           registers_62_9_port, C2 => n17658, A => n7417, ZN =>
                           n7414);
   U5658 : OAI22_X1 port map( A1 => n17655, A2 => n12410, B1 => n17652, B2 => 
                           n15335, ZN => n7417);
   U5659 : AOI221_X1 port map( B1 => registers_11_9_port, B2 => n17805, C1 => 
                           net227072, C2 => n17802, A => n7393, ZN => n7390);
   U5660 : OAI22_X1 port map( A1 => n17799, A2 => n15707, B1 => n17796, B2 => 
                           n11889, ZN => n7393);
   U5661 : AOI221_X1 port map( B1 => registers_63_10_port, B2 => n17661, C1 => 
                           registers_62_10_port, C2 => n17658, A => n7308, ZN 
                           => n7305);
   U5662 : OAI22_X1 port map( A1 => n17655, A2 => n12551, B1 => n17652, B2 => 
                           n15336, ZN => n7308);
   U5663 : AOI221_X1 port map( B1 => registers_11_10_port, B2 => n17805, C1 => 
                           net227090, C2 => n17802, A => n7284, ZN => n7281);
   U5664 : OAI22_X1 port map( A1 => n17799, A2 => n15708, B1 => n17796, B2 => 
                           n11890, ZN => n7284);
   U5665 : AOI221_X1 port map( B1 => registers_63_11_port, B2 => n17662, C1 => 
                           registers_62_11_port, C2 => n17659, A => n7194, ZN 
                           => n7191);
   U5666 : OAI22_X1 port map( A1 => n17656, A2 => n12602, B1 => n17653, B2 => 
                           n15337, ZN => n7194);
   U5667 : AOI221_X1 port map( B1 => registers_11_11_port, B2 => n17806, C1 => 
                           net227108, C2 => n17803, A => n7170, ZN => n7167);
   U5668 : OAI22_X1 port map( A1 => n17800, A2 => n15709, B1 => n17797, B2 => 
                           n11891, ZN => n7170);
   U5669 : AOI221_X1 port map( B1 => registers_63_12_port, B2 => n17662, C1 => 
                           registers_62_12_port, C2 => n17659, A => n7085, ZN 
                           => n7082);
   U5670 : OAI22_X1 port map( A1 => n17656, A2 => n12669, B1 => n17653, B2 => 
                           n15338, ZN => n7085);
   U5671 : AOI221_X1 port map( B1 => registers_11_12_port, B2 => n17806, C1 => 
                           net227126, C2 => n17803, A => n7061, ZN => n7058);
   U5672 : OAI22_X1 port map( A1 => n17800, A2 => n15710, B1 => n17797, B2 => 
                           n11892, ZN => n7061);
   U5673 : AOI221_X1 port map( B1 => registers_63_13_port, B2 => n17662, C1 => 
                           registers_62_13_port, C2 => n17659, A => n6976, ZN 
                           => n6973);
   U5674 : OAI22_X1 port map( A1 => n17656, A2 => n13999, B1 => n17653, B2 => 
                           n15339, ZN => n6976);
   U5675 : AOI221_X1 port map( B1 => registers_11_13_port, B2 => n17806, C1 => 
                           net227144, C2 => n17803, A => n6952, ZN => n6949);
   U5676 : OAI22_X1 port map( A1 => n17800, A2 => n15711, B1 => n17797, B2 => 
                           n11893, ZN => n6952);
   U5677 : AOI221_X1 port map( B1 => registers_63_14_port, B2 => n17662, C1 => 
                           registers_62_14_port, C2 => n17659, A => n6867, ZN 
                           => n6864);
   U5678 : OAI22_X1 port map( A1 => n17656, A2 => n14014, B1 => n17653, B2 => 
                           n15340, ZN => n6867);
   U5679 : AOI221_X1 port map( B1 => registers_11_14_port, B2 => n17806, C1 => 
                           net227162, C2 => n17803, A => n6843, ZN => n6840);
   U5680 : OAI22_X1 port map( A1 => n17800, A2 => n15712, B1 => n17797, B2 => 
                           n11894, ZN => n6843);
   U5681 : AOI221_X1 port map( B1 => registers_63_15_port, B2 => n17662, C1 => 
                           registers_62_15_port, C2 => n17659, A => n6758, ZN 
                           => n6755);
   U5682 : OAI22_X1 port map( A1 => n17656, A2 => n14032, B1 => n17653, B2 => 
                           n15341, ZN => n6758);
   U5683 : AOI221_X1 port map( B1 => registers_11_15_port, B2 => n17806, C1 => 
                           net227180, C2 => n17803, A => n6734, ZN => n6731);
   U5684 : OAI22_X1 port map( A1 => n17800, A2 => n15713, B1 => n17797, B2 => 
                           n11895, ZN => n6734);
   U5685 : AOI221_X1 port map( B1 => registers_63_16_port, B2 => n17662, C1 => 
                           registers_62_16_port, C2 => n17659, A => n6618, ZN 
                           => n6615);
   U5686 : OAI22_X1 port map( A1 => n17656, A2 => n14036, B1 => n17653, B2 => 
                           n15342, ZN => n6618);
   U5687 : AOI221_X1 port map( B1 => registers_11_16_port, B2 => n17806, C1 => 
                           net227198, C2 => n17803, A => n6574, ZN => n6570);
   U5688 : OAI22_X1 port map( A1 => n17800, A2 => n15714, B1 => n17797, B2 => 
                           n11896, ZN => n6574);
   U5689 : AOI221_X1 port map( B1 => registers_63_17_port, B2 => n17662, C1 => 
                           registers_62_17_port, C2 => n17659, A => n6433, ZN 
                           => n6428);
   U5690 : OAI22_X1 port map( A1 => n17656, A2 => n14038, B1 => n17653, B2 => 
                           n15343, ZN => n6433);
   U5691 : AOI221_X1 port map( B1 => registers_11_17_port, B2 => n17806, C1 => 
                           net227216, C2 => n17803, A => n6387, ZN => n6384);
   U5692 : OAI22_X1 port map( A1 => n17800, A2 => n15715, B1 => n17797, B2 => 
                           n11897, ZN => n6387);
   U5693 : AOI221_X1 port map( B1 => registers_63_18_port, B2 => n17662, C1 => 
                           registers_62_18_port, C2 => n17659, A => n6247, ZN 
                           => n6241);
   U5694 : OAI22_X1 port map( A1 => n17656, A2 => n14040, B1 => n17653, B2 => 
                           n15344, ZN => n6247);
   U5695 : AOI221_X1 port map( B1 => registers_11_18_port, B2 => n17806, C1 => 
                           net227234, C2 => n17803, A => n6202, ZN => n6197);
   U5696 : OAI22_X1 port map( A1 => n17800, A2 => n15716, B1 => n17797, B2 => 
                           n11898, ZN => n6202);
   U5697 : AOI221_X1 port map( B1 => registers_63_19_port, B2 => n17662, C1 => 
                           registers_62_19_port, C2 => n17659, A => n6060, ZN 
                           => n6056);
   U5698 : OAI22_X1 port map( A1 => n17656, A2 => n14042, B1 => n17653, B2 => 
                           n15345, ZN => n6060);
   U5699 : AOI221_X1 port map( B1 => registers_11_19_port, B2 => n17806, C1 => 
                           net227252, C2 => n17803, A => n6015, ZN => n6010);
   U5700 : OAI22_X1 port map( A1 => n17800, A2 => n15717, B1 => n17797, B2 => 
                           n11899, ZN => n6015);
   U5701 : AOI221_X1 port map( B1 => registers_63_20_port, B2 => n17662, C1 => 
                           registers_62_20_port, C2 => n17659, A => n5873, ZN 
                           => n5870);
   U5702 : OAI22_X1 port map( A1 => n17656, A2 => n14044, B1 => n17653, B2 => 
                           n15346, ZN => n5873);
   U5703 : AOI221_X1 port map( B1 => registers_11_20_port, B2 => n17806, C1 => 
                           net227270, C2 => n17803, A => n5843, ZN => n5825);
   U5704 : OAI22_X1 port map( A1 => n17800, A2 => n15718, B1 => n17797, B2 => 
                           n11900, ZN => n5843);
   U5705 : AOI221_X1 port map( B1 => registers_63_21_port, B2 => n17662, C1 => 
                           registers_62_21_port, C2 => n17659, A => n5688, ZN 
                           => n5683);
   U5706 : OAI22_X1 port map( A1 => n17656, A2 => n14046, B1 => n17653, B2 => 
                           n15347, ZN => n5688);
   U5707 : AOI221_X1 port map( B1 => registers_11_21_port, B2 => n17806, C1 => 
                           net227288, C2 => n17803, A => n5656, ZN => n5653);
   U5708 : OAI22_X1 port map( A1 => n17800, A2 => n15719, B1 => n17797, B2 => 
                           n11901, ZN => n5656);
   U5709 : AOI221_X1 port map( B1 => registers_63_22_port, B2 => n17662, C1 => 
                           registers_62_22_port, C2 => n17659, A => n5502, ZN 
                           => n5497);
   U5710 : OAI22_X1 port map( A1 => n17656, A2 => n14048, B1 => n17653, B2 => 
                           n15348, ZN => n5502);
   U5711 : AOI221_X1 port map( B1 => registers_11_22_port, B2 => n17806, C1 => 
                           net227306, C2 => n17803, A => n5469, ZN => n5466);
   U5712 : OAI22_X1 port map( A1 => n17800, A2 => n15720, B1 => n17797, B2 => 
                           n11902, ZN => n5469);
   U5713 : AOI221_X1 port map( B1 => registers_63_31_port, B2 => n17661, C1 => 
                           registers_62_31_port, C2 => n17658, A => n14198, ZN 
                           => n14189);
   U5714 : OAI22_X1 port map( A1 => n17655, A2 => n12348, B1 => n17652, B2 => 
                           n15349, ZN => n14198);
   U5715 : AOI221_X1 port map( B1 => registers_11_31_port, B2 => n17805, C1 => 
                           net227468, C2 => n17802, A => n14093, ZN => n14082);
   U5716 : OAI22_X1 port map( A1 => n17799, A2 => n15721, B1 => n17796, B2 => 
                           n11903, ZN => n14093);
   U5717 : OAI22_X1 port map( A1 => n7699, A2 => n17827, B1 => n4871, B2 => 
                           n17825, ZN => n9701);
   U5718 : NOR4_X1 port map( A1 => n4872, A2 => n4873, A3 => n4874, A4 => n4875
                           , ZN => n4871);
   U5719 : NAND4_X1 port map( A1 => n4876, A2 => n4877, A3 => n4878, A4 => 
                           n4879, ZN => n4875);
   U5720 : NAND4_X1 port map( A1 => n4906, A2 => n4907, A3 => n4908, A4 => 
                           n4909, ZN => n4872);
   U5721 : OAI22_X1 port map( A1 => n7698, A2 => n17826, B1 => n4738, B2 => 
                           n17825, ZN => n9773);
   U5722 : NOR4_X1 port map( A1 => n4739, A2 => n4740, A3 => n4741, A4 => n4742
                           , ZN => n4738);
   U5723 : NAND4_X1 port map( A1 => n4745, A2 => n4748, A3 => n4749, A4 => 
                           n4750, ZN => n4742);
   U5724 : NAND4_X1 port map( A1 => n4775, A2 => n4776, A3 => n4777, A4 => 
                           n4778, ZN => n4739);
   U5725 : OAI22_X1 port map( A1 => n7697, A2 => n17826, B1 => n4611, B2 => 
                           n17825, ZN => n9845);
   U5726 : NOR4_X1 port map( A1 => n4612, A2 => n4613, A3 => n4614, A4 => n4617
                           , ZN => n4611);
   U5727 : NAND4_X1 port map( A1 => n4618, A2 => n4619, A3 => n4620, A4 => 
                           n4621, ZN => n4617);
   U5728 : NAND4_X1 port map( A1 => n4642, A2 => n4645, A3 => n4648, A4 => 
                           n4649, ZN => n4612);
   U5729 : OAI22_X1 port map( A1 => n7696, A2 => n17826, B1 => n4480, B2 => 
                           n17825, ZN => n9917);
   U5730 : NOR4_X1 port map( A1 => n4481, A2 => n4482, A3 => n4483, A4 => n4484
                           , ZN => n4480);
   U5731 : NAND4_X1 port map( A1 => n4485, A2 => n4486, A3 => n4487, A4 => 
                           n4488, ZN => n4484);
   U5732 : NAND4_X1 port map( A1 => n4517, A2 => n4518, A3 => n4519, A4 => 
                           n4520, ZN => n4481);
   U5733 : OAI22_X1 port map( A1 => n7694, A2 => n17833, B1 => n14075, B2 => 
                           n17825, ZN => n10061);
   U5734 : NOR4_X1 port map( A1 => n14076, A2 => n14077, A3 => n14078, A4 => 
                           n14079, ZN => n14075);
   U5735 : NAND4_X1 port map( A1 => n14080, A2 => n14081, A3 => n14082, A4 => 
                           n14083, ZN => n14079);
   U5736 : NAND4_X1 port map( A1 => n14187, A2 => n14188, A3 => n14189, A4 => 
                           n14190, ZN => n14076);
   U5737 : AOI211_X1 port map( C1 => add_wr(4), C2 => add_wr(3), A => n14267, B
                           => n12514, ZN => n14232);
   U5738 : NOR4_X1 port map( A1 => n14213, A2 => add_wr(2), A3 => add_wr(4), A4
                           => add_wr(3), ZN => n14267);
   U5739 : AOI221_X1 port map( B1 => registers_47_24_port, B2 => n16291, C1 => 
                           registers_51_24_port, C2 => n16288, A => n12921, ZN 
                           => n12916);
   U5740 : OAI22_X1 port map( A1 => n16285, A2 => n15545, B1 => n16282, B2 => 
                           n14471, ZN => n12921);
   U5741 : AOI221_X1 port map( B1 => net227332, B2 => n16240, C1 => n16237, C2 
                           => datain(24), A => n12929, ZN => n12924);
   U5742 : OAI22_X1 port map( A1 => n16234, A2 => n15117, B1 => n16231, B2 => 
                           n14478, ZN => n12929);
   U5743 : AOI221_X1 port map( B1 => registers_47_25_port, B2 => n16291, C1 => 
                           registers_51_25_port, C2 => n16288, A => n12879, ZN 
                           => n12874);
   U5744 : OAI22_X1 port map( A1 => n16285, A2 => n15546, B1 => n16282, B2 => 
                           n14472, ZN => n12879);
   U5745 : AOI221_X1 port map( B1 => net227350, B2 => n16240, C1 => n16237, C2 
                           => datain(25), A => n12887, ZN => n12882);
   U5746 : OAI22_X1 port map( A1 => n16234, A2 => n15118, B1 => n16231, B2 => 
                           n14479, ZN => n12887);
   U5747 : AOI221_X1 port map( B1 => registers_47_26_port, B2 => n16291, C1 => 
                           registers_51_26_port, C2 => n16288, A => n12837, ZN 
                           => n12832);
   U5748 : OAI22_X1 port map( A1 => n16285, A2 => n15547, B1 => n16282, B2 => 
                           n14473, ZN => n12837);
   U5749 : AOI221_X1 port map( B1 => net227368, B2 => n16240, C1 => n16237, C2 
                           => datain(26), A => n12845, ZN => n12840);
   U5750 : OAI22_X1 port map( A1 => n16234, A2 => n15119, B1 => n16231, B2 => 
                           n14480, ZN => n12845);
   U5751 : AOI221_X1 port map( B1 => registers_47_27_port, B2 => n16291, C1 => 
                           registers_51_27_port, C2 => n16288, A => n12795, ZN 
                           => n12790);
   U5752 : OAI22_X1 port map( A1 => n16285, A2 => n15548, B1 => n16282, B2 => 
                           n14474, ZN => n12795);
   U5753 : AOI221_X1 port map( B1 => net227386, B2 => n16240, C1 => n16237, C2 
                           => datain(27), A => n12803, ZN => n12798);
   U5754 : OAI22_X1 port map( A1 => n16234, A2 => n15120, B1 => n16231, B2 => 
                           n14481, ZN => n12803);
   U5755 : AOI221_X1 port map( B1 => registers_47_28_port, B2 => n16291, C1 => 
                           registers_51_28_port, C2 => n16288, A => n12753, ZN 
                           => n12748);
   U5756 : OAI22_X1 port map( A1 => n16285, A2 => n15549, B1 => n16282, B2 => 
                           n14475, ZN => n12753);
   U5757 : AOI221_X1 port map( B1 => net227404, B2 => n16240, C1 => n16237, C2 
                           => datain(28), A => n12761, ZN => n12756);
   U5758 : OAI22_X1 port map( A1 => n16234, A2 => n15121, B1 => n16231, B2 => 
                           n14482, ZN => n12761);
   U5759 : AOI221_X1 port map( B1 => registers_47_29_port, B2 => n16291, C1 => 
                           registers_51_29_port, C2 => n16288, A => n12711, ZN 
                           => n12706);
   U5760 : OAI22_X1 port map( A1 => n16285, A2 => n15550, B1 => n16282, B2 => 
                           n14476, ZN => n12711);
   U5761 : AOI221_X1 port map( B1 => net227422, B2 => n16240, C1 => n16237, C2 
                           => datain(29), A => n12719, ZN => n12714);
   U5762 : OAI22_X1 port map( A1 => n16234, A2 => n15122, B1 => n16231, B2 => 
                           n14483, ZN => n12719);
   U5763 : AOI221_X1 port map( B1 => registers_47_30_port, B2 => n16291, C1 => 
                           registers_51_30_port, C2 => n16288, A => n12668, ZN 
                           => n12663);
   U5764 : OAI22_X1 port map( A1 => n16285, A2 => n15277, B1 => n16282, B2 => 
                           n14065, ZN => n12668);
   U5765 : AOI221_X1 port map( B1 => net227440, B2 => n16240, C1 => n16237, C2 
                           => datain(30), A => n12677, ZN => n12672);
   U5766 : OAI22_X1 port map( A1 => n16234, A2 => n14991, B1 => n16231, B2 => 
                           n14280, ZN => n12677);
   U5767 : AOI221_X1 port map( B1 => registers_47_31_port, B2 => n16291, C1 => 
                           registers_51_31_port, C2 => n16288, A => n12598, ZN 
                           => n12583);
   U5768 : OAI22_X1 port map( A1 => n16285, A2 => n15551, B1 => n16282, B2 => 
                           n14477, ZN => n12598);
   U5769 : AOI221_X1 port map( B1 => net227458, B2 => n16240, C1 => n16237, C2 
                           => datain(31), A => n12625, ZN => n12609);
   U5770 : OAI22_X1 port map( A1 => n16234, A2 => n14992, B1 => n16231, B2 => 
                           n14281, ZN => n12625);
   U5771 : AOI221_X1 port map( B1 => registers_49_24_port, B2 => n16543, C1 => 
                           registers_51_24_port, C2 => n16540, A => n10971, ZN 
                           => n10966);
   U5772 : OAI22_X1 port map( A1 => n16537, A2 => n15452, B1 => n16534, B2 => 
                           n14540, ZN => n10971);
   U5773 : AOI221_X1 port map( B1 => net227332, B2 => n16492, C1 => n16488, C2 
                           => datain(24), A => n10979, ZN => n10974);
   U5774 : OAI22_X1 port map( A1 => n16486, A2 => n15117, B1 => n16483, B2 => 
                           n14478, ZN => n10979);
   U5775 : AOI221_X1 port map( B1 => registers_49_25_port, B2 => n16543, C1 => 
                           registers_51_25_port, C2 => n16540, A => n10928, ZN 
                           => n10923);
   U5776 : OAI22_X1 port map( A1 => n16537, A2 => n15453, B1 => n16534, B2 => 
                           n14541, ZN => n10928);
   U5777 : AOI221_X1 port map( B1 => net227350, B2 => n16492, C1 => n16488, C2 
                           => datain(25), A => n10936, ZN => n10931);
   U5778 : OAI22_X1 port map( A1 => n16486, A2 => n15118, B1 => n16483, B2 => 
                           n14479, ZN => n10936);
   U5779 : AOI221_X1 port map( B1 => registers_49_26_port, B2 => n16543, C1 => 
                           registers_51_26_port, C2 => n16540, A => n10885, ZN 
                           => n10880);
   U5780 : OAI22_X1 port map( A1 => n16537, A2 => n15454, B1 => n16534, B2 => 
                           n14542, ZN => n10885);
   U5781 : AOI221_X1 port map( B1 => net227368, B2 => n16492, C1 => n16489, C2 
                           => datain(26), A => n10893, ZN => n10888);
   U5782 : OAI22_X1 port map( A1 => n16486, A2 => n15119, B1 => n16483, B2 => 
                           n14480, ZN => n10893);
   U5783 : AOI221_X1 port map( B1 => registers_49_27_port, B2 => n16543, C1 => 
                           registers_51_27_port, C2 => n16540, A => n10842, ZN 
                           => n10837);
   U5784 : OAI22_X1 port map( A1 => n16537, A2 => n15455, B1 => n16534, B2 => 
                           n14543, ZN => n10842);
   U5785 : AOI221_X1 port map( B1 => net227386, B2 => n16492, C1 => n16489, C2 
                           => datain(27), A => n10850, ZN => n10845);
   U5786 : OAI22_X1 port map( A1 => n16486, A2 => n15120, B1 => n16483, B2 => 
                           n14481, ZN => n10850);
   U5787 : AOI221_X1 port map( B1 => registers_49_28_port, B2 => n16543, C1 => 
                           registers_51_28_port, C2 => n16540, A => n10799, ZN 
                           => n10794);
   U5788 : OAI22_X1 port map( A1 => n16537, A2 => n15456, B1 => n16534, B2 => 
                           n14544, ZN => n10799);
   U5789 : AOI221_X1 port map( B1 => net227404, B2 => n16492, C1 => n16489, C2 
                           => datain(28), A => n10807, ZN => n10802);
   U5790 : OAI22_X1 port map( A1 => n16486, A2 => n15121, B1 => n16483, B2 => 
                           n14482, ZN => n10807);
   U5791 : AOI221_X1 port map( B1 => registers_49_29_port, B2 => n16543, C1 => 
                           registers_51_29_port, C2 => n16540, A => n10756, ZN 
                           => n10751);
   U5792 : OAI22_X1 port map( A1 => n16537, A2 => n15457, B1 => n16534, B2 => 
                           n14545, ZN => n10756);
   U5793 : AOI221_X1 port map( B1 => net227422, B2 => n16492, C1 => n16489, C2 
                           => datain(29), A => n10764, ZN => n10759);
   U5794 : OAI22_X1 port map( A1 => n16486, A2 => n15122, B1 => n16483, B2 => 
                           n14483, ZN => n10764);
   U5795 : AOI221_X1 port map( B1 => registers_49_30_port, B2 => n16543, C1 => 
                           registers_51_30_port, C2 => n16540, A => n10709, ZN 
                           => n10701);
   U5796 : OAI22_X1 port map( A1 => n16537, A2 => n15274, B1 => n16534, B2 => 
                           n14279, ZN => n10709);
   U5797 : AOI221_X1 port map( B1 => net227440, B2 => n16492, C1 => n16489, C2 
                           => datain(30), A => n10719, ZN => n10714);
   U5798 : OAI22_X1 port map( A1 => n16486, A2 => n14991, B1 => n16483, B2 => 
                           n14280, ZN => n10719);
   U5799 : AOI221_X1 port map( B1 => registers_49_31_port, B2 => n16543, C1 => 
                           registers_51_31_port, C2 => n16540, A => n10616, ZN 
                           => n10597);
   U5800 : OAI22_X1 port map( A1 => n16537, A2 => n15458, B1 => n16534, B2 => 
                           n14546, ZN => n10616);
   U5801 : AOI221_X1 port map( B1 => net227458, B2 => n16492, C1 => n16489, C2 
                           => datain(31), A => n10650, ZN => n10629);
   U5802 : OAI22_X1 port map( A1 => n16486, A2 => n14992, B1 => n16483, B2 => 
                           n14281, ZN => n10650);
   U5803 : AOI221_X1 port map( B1 => net227322, B2 => n17747, C1 => 
                           registers_29_23_port, C2 => n17744, A => n5294, ZN 
                           => n5288);
   U5804 : OAI22_X1 port map( A1 => n17741, A2 => n15722, B1 => n17738, B2 => 
                           n14757, ZN => n5294);
   U5805 : AOI221_X1 port map( B1 => net227325, B2 => n17699, C1 => 
                           registers_9_23_port, C2 => n17696, A => n5305, ZN =>
                           n5299);
   U5806 : OAI22_X1 port map( A1 => n17693, A2 => n15723, B1 => n17690, B2 => 
                           n12164, ZN => n5305);
   U5807 : AOI221_X1 port map( B1 => registers_41_23_port, B2 => n17651, C1 => 
                           registers_40_23_port, C2 => n17648, A => n5316, ZN 
                           => n5311);
   U5808 : OAI22_X1 port map( A1 => n17645, A2 => n15459, B1 => n17642, B2 => 
                           n14758, ZN => n5316);
   U5809 : AOI221_X1 port map( B1 => registers_18_23_port, B2 => n17795, C1 => 
                           registers_19_23_port, C2 => n17792, A => n5283, ZN 
                           => n5278);
   U5810 : OAI22_X1 port map( A1 => n17789, A2 => n14598, B1 => n17786, B2 => 
                           n15285, ZN => n5283);
   U5811 : AOI221_X1 port map( B1 => net227340, B2 => n17747, C1 => 
                           registers_29_24_port, C2 => n17744, A => n5128, ZN 
                           => n5121);
   U5812 : OAI22_X1 port map( A1 => n17741, A2 => n15724, B1 => n17738, B2 => 
                           n14759, ZN => n5128);
   U5813 : AOI221_X1 port map( B1 => net227343, B2 => n17699, C1 => 
                           registers_9_24_port, C2 => n17696, A => n5136, ZN =>
                           n5131);
   U5814 : OAI22_X1 port map( A1 => n17693, A2 => n15725, B1 => n17690, B2 => 
                           n12165, ZN => n5136);
   U5815 : AOI221_X1 port map( B1 => registers_41_24_port, B2 => n17651, C1 => 
                           registers_40_24_port, C2 => n17648, A => n5146, ZN 
                           => n5139);
   U5816 : OAI22_X1 port map( A1 => n17645, A2 => n15460, B1 => n17642, B2 => 
                           n14760, ZN => n5146);
   U5817 : AOI221_X1 port map( B1 => registers_18_24_port, B2 => n17795, C1 => 
                           registers_19_24_port, C2 => n17792, A => n5118, ZN 
                           => n5112);
   U5818 : OAI22_X1 port map( A1 => n17789, A2 => n14599, B1 => n17786, B2 => 
                           n15286, ZN => n5118);
   U5819 : AOI221_X1 port map( B1 => net227358, B2 => n17747, C1 => 
                           registers_29_25_port, C2 => n17744, A => n5012, ZN 
                           => n5007);
   U5820 : OAI22_X1 port map( A1 => n17741, A2 => n15726, B1 => n17738, B2 => 
                           n14761, ZN => n5012);
   U5821 : AOI221_X1 port map( B1 => net227361, B2 => n17699, C1 => 
                           registers_9_25_port, C2 => n17696, A => n5022, ZN =>
                           n5015);
   U5822 : OAI22_X1 port map( A1 => n17693, A2 => n15727, B1 => n17690, B2 => 
                           n12166, ZN => n5022);
   U5823 : AOI221_X1 port map( B1 => registers_41_25_port, B2 => n17651, C1 => 
                           registers_40_25_port, C2 => n17648, A => n5030, ZN 
                           => n5025);
   U5824 : OAI22_X1 port map( A1 => n17645, A2 => n15461, B1 => n17642, B2 => 
                           n14762, ZN => n5030);
   U5825 : AOI221_X1 port map( B1 => registers_18_25_port, B2 => n17795, C1 => 
                           registers_19_25_port, C2 => n17792, A => n5004, ZN 
                           => n4999);
   U5826 : OAI22_X1 port map( A1 => n17789, A2 => n14600, B1 => n17786, B2 => 
                           n15287, ZN => n5004);
   U5827 : AOI221_X1 port map( B1 => net227376, B2 => n17747, C1 => 
                           registers_29_26_port, C2 => n17744, A => n4890, ZN 
                           => n4885);
   U5828 : OAI22_X1 port map( A1 => n17741, A2 => n15728, B1 => n17738, B2 => 
                           n14763, ZN => n4890);
   U5829 : AOI221_X1 port map( B1 => net227379, B2 => n17699, C1 => 
                           registers_9_26_port, C2 => n17696, A => n4902, ZN =>
                           n4895);
   U5830 : OAI22_X1 port map( A1 => n17693, A2 => n15729, B1 => n17690, B2 => 
                           n12167, ZN => n4902);
   U5831 : AOI221_X1 port map( B1 => registers_41_26_port, B2 => n17651, C1 => 
                           registers_40_26_port, C2 => n17648, A => n4912, ZN 
                           => n4907);
   U5832 : OAI22_X1 port map( A1 => n17645, A2 => n15462, B1 => n17642, B2 => 
                           n14764, ZN => n4912);
   U5833 : AOI221_X1 port map( B1 => registers_18_26_port, B2 => n17795, C1 => 
                           registers_19_26_port, C2 => n17792, A => n4882, ZN 
                           => n4877);
   U5834 : OAI22_X1 port map( A1 => n17789, A2 => n14601, B1 => n17786, B2 => 
                           n15288, ZN => n4882);
   U5835 : AOI221_X1 port map( B1 => net227394, B2 => n17747, C1 => 
                           registers_29_27_port, C2 => n17744, A => n4763, ZN 
                           => n4758);
   U5836 : OAI22_X1 port map( A1 => n17741, A2 => n15730, B1 => n17738, B2 => 
                           n14765, ZN => n4763);
   U5837 : AOI221_X1 port map( B1 => net227397, B2 => n17699, C1 => 
                           registers_9_27_port, C2 => n17696, A => n4773, ZN =>
                           n4768);
   U5838 : OAI22_X1 port map( A1 => n17693, A2 => n15731, B1 => n17690, B2 => 
                           n12168, ZN => n4773);
   U5839 : AOI221_X1 port map( B1 => registers_41_27_port, B2 => n17651, C1 => 
                           registers_40_27_port, C2 => n17648, A => n4781, ZN 
                           => n4776);
   U5840 : OAI22_X1 port map( A1 => n17645, A2 => n15463, B1 => n17642, B2 => 
                           n14766, ZN => n4781);
   U5841 : AOI221_X1 port map( B1 => registers_18_27_port, B2 => n17795, C1 => 
                           registers_19_27_port, C2 => n17792, A => n4753, ZN 
                           => n4748);
   U5842 : OAI22_X1 port map( A1 => n17789, A2 => n14602, B1 => n17786, B2 => 
                           n15289, ZN => n4753);
   U5843 : AOI221_X1 port map( B1 => net227412, B2 => n17747, C1 => 
                           registers_29_28_port, C2 => n17744, A => n4632, ZN 
                           => n4627);
   U5844 : OAI22_X1 port map( A1 => n17741, A2 => n15732, B1 => n17738, B2 => 
                           n14767, ZN => n4632);
   U5845 : AOI221_X1 port map( B1 => net227415, B2 => n17699, C1 => 
                           registers_9_28_port, C2 => n17696, A => n4640, ZN =>
                           n4635);
   U5846 : OAI22_X1 port map( A1 => n17693, A2 => n15733, B1 => n17690, B2 => 
                           n12169, ZN => n4640);
   U5847 : AOI221_X1 port map( B1 => registers_41_28_port, B2 => n17651, C1 => 
                           registers_40_28_port, C2 => n17648, A => n4652, ZN 
                           => n4645);
   U5848 : OAI22_X1 port map( A1 => n17645, A2 => n15464, B1 => n17642, B2 => 
                           n14768, ZN => n4652);
   U5849 : AOI221_X1 port map( B1 => registers_18_28_port, B2 => n17795, C1 => 
                           registers_19_28_port, C2 => n17792, A => n4624, ZN 
                           => n4619);
   U5850 : OAI22_X1 port map( A1 => n17789, A2 => n14603, B1 => n17786, B2 => 
                           n15290, ZN => n4624);
   U5851 : AOI221_X1 port map( B1 => net227430, B2 => n17747, C1 => 
                           registers_29_29_port, C2 => n17744, A => n4503, ZN 
                           => n4498);
   U5852 : OAI22_X1 port map( A1 => n17741, A2 => n15734, B1 => n17738, B2 => 
                           n14769, ZN => n4503);
   U5853 : AOI221_X1 port map( B1 => net227433, B2 => n17699, C1 => 
                           registers_9_29_port, C2 => n17696, A => n4513, ZN =>
                           n4508);
   U5854 : OAI22_X1 port map( A1 => n17693, A2 => n15735, B1 => n17690, B2 => 
                           n12170, ZN => n4513);
   U5855 : AOI221_X1 port map( B1 => registers_41_29_port, B2 => n17651, C1 => 
                           registers_40_29_port, C2 => n17648, A => n4523, ZN 
                           => n4518);
   U5856 : OAI22_X1 port map( A1 => n17645, A2 => n15465, B1 => n17642, B2 => 
                           n14770, ZN => n4523);
   U5857 : AOI221_X1 port map( B1 => registers_18_29_port, B2 => n17795, C1 => 
                           registers_19_29_port, C2 => n17792, A => n4491, ZN 
                           => n4486);
   U5858 : OAI22_X1 port map( A1 => n17789, A2 => n14604, B1 => n17786, B2 => 
                           n15291, ZN => n4491);
   U5859 : AOI221_X1 port map( B1 => net227448, B2 => n17747, C1 => 
                           registers_29_30_port, C2 => n17744, A => n4163, ZN 
                           => n4138);
   U5860 : OAI22_X1 port map( A1 => n17741, A2 => n15282, B1 => n17738, B2 => 
                           n14630, ZN => n4163);
   U5861 : AOI221_X1 port map( B1 => net227451, B2 => n17699, C1 => 
                           registers_9_30_port, C2 => n17696, A => n4199, ZN =>
                           n4178);
   U5862 : OAI22_X1 port map( A1 => n17693, A2 => n15283, B1 => n17690, B2 => 
                           n12160, ZN => n4199);
   U5863 : AOI221_X1 port map( B1 => registers_41_30_port, B2 => n17651, C1 => 
                           registers_40_30_port, C2 => n17648, A => n4234, ZN 
                           => n4214);
   U5864 : OAI22_X1 port map( A1 => n17645, A2 => n15275, B1 => n17642, B2 => 
                           n14631, ZN => n4234);
   U5865 : AOI221_X1 port map( B1 => registers_18_30_port, B2 => n17795, C1 => 
                           registers_19_30_port, C2 => n17792, A => n4125, ZN 
                           => n4102);
   U5866 : OAI22_X1 port map( A1 => n17789, A2 => n14299, B1 => n17786, B2 => 
                           n15270, ZN => n4125);
   U5867 : AOI221_X1 port map( B1 => registers_47_0_port, B2 => n16289, C1 => 
                           registers_51_0_port, C2 => n16286, A => n13956, ZN 
                           => n13949);
   U5868 : OAI22_X1 port map( A1 => n16283, A2 => n15552, B1 => n16280, B2 => 
                           n14484, ZN => n13956);
   U5869 : AOI221_X1 port map( B1 => net226844, B2 => n16238, C1 => n16235, C2 
                           => datain(0), A => n13972, ZN => n13965);
   U5870 : OAI22_X1 port map( A1 => n16232, A2 => n15123, B1 => n16229, B2 => 
                           n14506, ZN => n13972);
   U5871 : AOI221_X1 port map( B1 => registers_47_1_port, B2 => n16289, C1 => 
                           registers_51_1_port, C2 => n16286, A => n13887, ZN 
                           => n13882);
   U5872 : OAI22_X1 port map( A1 => n16283, A2 => n15553, B1 => n16280, B2 => 
                           n14485, ZN => n13887);
   U5873 : AOI221_X1 port map( B1 => net226857, B2 => n16238, C1 => n16235, C2 
                           => datain(1), A => n13895, ZN => n13890);
   U5874 : OAI22_X1 port map( A1 => n16232, A2 => n15124, B1 => n16229, B2 => 
                           n14507, ZN => n13895);
   U5875 : AOI221_X1 port map( B1 => registers_47_2_port, B2 => n16289, C1 => 
                           registers_51_2_port, C2 => n16286, A => n13845, ZN 
                           => n13840);
   U5876 : OAI22_X1 port map( A1 => n16283, A2 => n15554, B1 => n16280, B2 => 
                           n14486, ZN => n13845);
   U5877 : AOI221_X1 port map( B1 => net226884, B2 => n16238, C1 => n16235, C2 
                           => datain(2), A => n13853, ZN => n13848);
   U5878 : OAI22_X1 port map( A1 => n16232, A2 => n15125, B1 => n16229, B2 => 
                           n14508, ZN => n13853);
   U5879 : AOI221_X1 port map( B1 => registers_47_3_port, B2 => n16289, C1 => 
                           registers_51_3_port, C2 => n16286, A => n13803, ZN 
                           => n13798);
   U5880 : OAI22_X1 port map( A1 => n16283, A2 => n15555, B1 => n16280, B2 => 
                           n14487, ZN => n13803);
   U5881 : AOI221_X1 port map( B1 => net226904, B2 => n16238, C1 => n16235, C2 
                           => datain(3), A => n13811, ZN => n13806);
   U5882 : OAI22_X1 port map( A1 => n16232, A2 => n14997, B1 => n16229, B2 => 
                           n14296, ZN => n13811);
   U5883 : AOI221_X1 port map( B1 => registers_47_4_port, B2 => n16289, C1 => 
                           registers_51_4_port, C2 => n16286, A => n13761, ZN 
                           => n13756);
   U5884 : OAI22_X1 port map( A1 => n16283, A2 => n15359, B1 => n16280, B2 => 
                           n14294, ZN => n13761);
   U5885 : AOI221_X1 port map( B1 => net226977, B2 => n16238, C1 => n16235, C2 
                           => datain(4), A => n13769, ZN => n13764);
   U5886 : OAI22_X1 port map( A1 => n16232, A2 => n14998, B1 => n16229, B2 => 
                           n14297, ZN => n13769);
   U5887 : AOI221_X1 port map( B1 => registers_47_5_port, B2 => n16289, C1 => 
                           registers_51_5_port, C2 => n16286, A => n13719, ZN 
                           => n13714);
   U5888 : OAI22_X1 port map( A1 => n16283, A2 => n15360, B1 => n16280, B2 => 
                           n14295, ZN => n13719);
   U5889 : AOI221_X1 port map( B1 => net226997, B2 => n16238, C1 => n16235, C2 
                           => datain(5), A => n13727, ZN => n13722);
   U5890 : OAI22_X1 port map( A1 => n16232, A2 => n14999, B1 => n16229, B2 => 
                           n14298, ZN => n13727);
   U5891 : AOI221_X1 port map( B1 => registers_47_6_port, B2 => n16289, C1 => 
                           registers_51_6_port, C2 => n16286, A => n13677, ZN 
                           => n13672);
   U5892 : OAI22_X1 port map( A1 => n16283, A2 => n15556, B1 => n16280, B2 => 
                           n14488, ZN => n13677);
   U5893 : AOI221_X1 port map( B1 => net227008, B2 => n16238, C1 => n16235, C2 
                           => datain(6), A => n13685, ZN => n13680);
   U5894 : OAI22_X1 port map( A1 => n16232, A2 => n15126, B1 => n16229, B2 => 
                           n14509, ZN => n13685);
   U5895 : AOI221_X1 port map( B1 => registers_47_7_port, B2 => n16289, C1 => 
                           registers_51_7_port, C2 => n16286, A => n13635, ZN 
                           => n13630);
   U5896 : OAI22_X1 port map( A1 => n16283, A2 => n15557, B1 => n16280, B2 => 
                           n14489, ZN => n13635);
   U5897 : AOI221_X1 port map( B1 => net227026, B2 => n16238, C1 => n16235, C2 
                           => datain(7), A => n13643, ZN => n13638);
   U5898 : OAI22_X1 port map( A1 => n16232, A2 => n15127, B1 => n16229, B2 => 
                           n14510, ZN => n13643);
   U5899 : AOI221_X1 port map( B1 => registers_47_8_port, B2 => n16289, C1 => 
                           registers_51_8_port, C2 => n16286, A => n13593, ZN 
                           => n13588);
   U5900 : OAI22_X1 port map( A1 => n16283, A2 => n15558, B1 => n16280, B2 => 
                           n14490, ZN => n13593);
   U5901 : AOI221_X1 port map( B1 => net227044, B2 => n16238, C1 => n16235, C2 
                           => datain(8), A => n13601, ZN => n13596);
   U5902 : OAI22_X1 port map( A1 => n16232, A2 => n15128, B1 => n16229, B2 => 
                           n14511, ZN => n13601);
   U5903 : AOI221_X1 port map( B1 => registers_47_9_port, B2 => n16289, C1 => 
                           registers_51_9_port, C2 => n16286, A => n13551, ZN 
                           => n13546);
   U5904 : OAI22_X1 port map( A1 => n16283, A2 => n15559, B1 => n16280, B2 => 
                           n14491, ZN => n13551);
   U5905 : AOI221_X1 port map( B1 => net227062, B2 => n16238, C1 => n16235, C2 
                           => datain(9), A => n13559, ZN => n13554);
   U5906 : OAI22_X1 port map( A1 => n16232, A2 => n15129, B1 => n16229, B2 => 
                           n14512, ZN => n13559);
   U5907 : AOI221_X1 port map( B1 => registers_47_10_port, B2 => n16289, C1 => 
                           registers_51_10_port, C2 => n16286, A => n13509, ZN 
                           => n13504);
   U5908 : OAI22_X1 port map( A1 => n16283, A2 => n15560, B1 => n16280, B2 => 
                           n14492, ZN => n13509);
   U5909 : AOI221_X1 port map( B1 => net227080, B2 => n16238, C1 => n16235, C2 
                           => datain(10), A => n13517, ZN => n13512);
   U5910 : OAI22_X1 port map( A1 => n16232, A2 => n15130, B1 => n16229, B2 => 
                           n14513, ZN => n13517);
   U5911 : AOI221_X1 port map( B1 => registers_47_11_port, B2 => n16289, C1 => 
                           registers_51_11_port, C2 => n16286, A => n13467, ZN 
                           => n13462);
   U5912 : OAI22_X1 port map( A1 => n16283, A2 => n15561, B1 => n16280, B2 => 
                           n14493, ZN => n13467);
   U5913 : AOI221_X1 port map( B1 => net227098, B2 => n16238, C1 => n16235, C2 
                           => datain(11), A => n13475, ZN => n13470);
   U5914 : OAI22_X1 port map( A1 => n16232, A2 => n15131, B1 => n16229, B2 => 
                           n14514, ZN => n13475);
   U5915 : AOI221_X1 port map( B1 => registers_47_12_port, B2 => n16290, C1 => 
                           registers_51_12_port, C2 => n16287, A => n13425, ZN 
                           => n13420);
   U5916 : OAI22_X1 port map( A1 => n16284, A2 => n15562, B1 => n16281, B2 => 
                           n14494, ZN => n13425);
   U5917 : AOI221_X1 port map( B1 => net227116, B2 => n16239, C1 => n16236, C2 
                           => datain(12), A => n13433, ZN => n13428);
   U5918 : OAI22_X1 port map( A1 => n16233, A2 => n15132, B1 => n16230, B2 => 
                           n14515, ZN => n13433);
   U5919 : AOI221_X1 port map( B1 => registers_47_13_port, B2 => n16290, C1 => 
                           registers_51_13_port, C2 => n16287, A => n13383, ZN 
                           => n13378);
   U5920 : OAI22_X1 port map( A1 => n16284, A2 => n15563, B1 => n16281, B2 => 
                           n14495, ZN => n13383);
   U5921 : AOI221_X1 port map( B1 => net227134, B2 => n16239, C1 => n16236, C2 
                           => datain(13), A => n13391, ZN => n13386);
   U5922 : OAI22_X1 port map( A1 => n16233, A2 => n15133, B1 => n16230, B2 => 
                           n14516, ZN => n13391);
   U5923 : AOI221_X1 port map( B1 => registers_47_14_port, B2 => n16290, C1 => 
                           registers_51_14_port, C2 => n16287, A => n13341, ZN 
                           => n13336);
   U5924 : OAI22_X1 port map( A1 => n16284, A2 => n15564, B1 => n16281, B2 => 
                           n14496, ZN => n13341);
   U5925 : AOI221_X1 port map( B1 => net227152, B2 => n16239, C1 => n16236, C2 
                           => datain(14), A => n13349, ZN => n13344);
   U5926 : OAI22_X1 port map( A1 => n16233, A2 => n15134, B1 => n16230, B2 => 
                           n14517, ZN => n13349);
   U5927 : AOI221_X1 port map( B1 => registers_47_15_port, B2 => n16290, C1 => 
                           registers_51_15_port, C2 => n16287, A => n13299, ZN 
                           => n13294);
   U5928 : OAI22_X1 port map( A1 => n16284, A2 => n15565, B1 => n16281, B2 => 
                           n14497, ZN => n13299);
   U5929 : AOI221_X1 port map( B1 => net227170, B2 => n16239, C1 => n16236, C2 
                           => datain(15), A => n13307, ZN => n13302);
   U5930 : OAI22_X1 port map( A1 => n16233, A2 => n15135, B1 => n16230, B2 => 
                           n14518, ZN => n13307);
   U5931 : AOI221_X1 port map( B1 => registers_47_16_port, B2 => n16290, C1 => 
                           registers_51_16_port, C2 => n16287, A => n13257, ZN 
                           => n13252);
   U5932 : OAI22_X1 port map( A1 => n16284, A2 => n15566, B1 => n16281, B2 => 
                           n14498, ZN => n13257);
   U5933 : AOI221_X1 port map( B1 => net227188, B2 => n16239, C1 => n16236, C2 
                           => datain(16), A => n13265, ZN => n13260);
   U5934 : OAI22_X1 port map( A1 => n16233, A2 => n15136, B1 => n16230, B2 => 
                           n14519, ZN => n13265);
   U5935 : AOI221_X1 port map( B1 => registers_47_17_port, B2 => n16290, C1 => 
                           registers_51_17_port, C2 => n16287, A => n13215, ZN 
                           => n13210);
   U5936 : OAI22_X1 port map( A1 => n16284, A2 => n15567, B1 => n16281, B2 => 
                           n14499, ZN => n13215);
   U5937 : AOI221_X1 port map( B1 => net227206, B2 => n16239, C1 => n16236, C2 
                           => datain(17), A => n13223, ZN => n13218);
   U5938 : OAI22_X1 port map( A1 => n16233, A2 => n15137, B1 => n16230, B2 => 
                           n14520, ZN => n13223);
   U5939 : AOI221_X1 port map( B1 => registers_47_18_port, B2 => n16290, C1 => 
                           registers_51_18_port, C2 => n16287, A => n13173, ZN 
                           => n13168);
   U5940 : OAI22_X1 port map( A1 => n16284, A2 => n15568, B1 => n16281, B2 => 
                           n14500, ZN => n13173);
   U5941 : AOI221_X1 port map( B1 => net227224, B2 => n16239, C1 => n16236, C2 
                           => datain(18), A => n13181, ZN => n13176);
   U5942 : OAI22_X1 port map( A1 => n16233, A2 => n15138, B1 => n16230, B2 => 
                           n14521, ZN => n13181);
   U5943 : AOI221_X1 port map( B1 => registers_47_19_port, B2 => n16290, C1 => 
                           registers_51_19_port, C2 => n16287, A => n13131, ZN 
                           => n13126);
   U5944 : OAI22_X1 port map( A1 => n16284, A2 => n15569, B1 => n16281, B2 => 
                           n14501, ZN => n13131);
   U5945 : AOI221_X1 port map( B1 => net227242, B2 => n16239, C1 => n16236, C2 
                           => datain(19), A => n13139, ZN => n13134);
   U5946 : OAI22_X1 port map( A1 => n16233, A2 => n15139, B1 => n16230, B2 => 
                           n14522, ZN => n13139);
   U5947 : AOI221_X1 port map( B1 => registers_47_20_port, B2 => n16290, C1 => 
                           registers_51_20_port, C2 => n16287, A => n13089, ZN 
                           => n13084);
   U5948 : OAI22_X1 port map( A1 => n16284, A2 => n15570, B1 => n16281, B2 => 
                           n14502, ZN => n13089);
   U5949 : AOI221_X1 port map( B1 => net227260, B2 => n16239, C1 => n16236, C2 
                           => datain(20), A => n13097, ZN => n13092);
   U5950 : OAI22_X1 port map( A1 => n16233, A2 => n15140, B1 => n16230, B2 => 
                           n14523, ZN => n13097);
   U5951 : AOI221_X1 port map( B1 => registers_47_21_port, B2 => n16290, C1 => 
                           registers_51_21_port, C2 => n16287, A => n13047, ZN 
                           => n13042);
   U5952 : OAI22_X1 port map( A1 => n16284, A2 => n15571, B1 => n16281, B2 => 
                           n14503, ZN => n13047);
   U5953 : AOI221_X1 port map( B1 => net227278, B2 => n16239, C1 => n16236, C2 
                           => datain(21), A => n13055, ZN => n13050);
   U5954 : OAI22_X1 port map( A1 => n16233, A2 => n15141, B1 => n16230, B2 => 
                           n14524, ZN => n13055);
   U5955 : AOI221_X1 port map( B1 => registers_47_22_port, B2 => n16290, C1 => 
                           registers_51_22_port, C2 => n16287, A => n13005, ZN 
                           => n13000);
   U5956 : OAI22_X1 port map( A1 => n16284, A2 => n15572, B1 => n16281, B2 => 
                           n14504, ZN => n13005);
   U5957 : AOI221_X1 port map( B1 => net227296, B2 => n16239, C1 => n16236, C2 
                           => datain(22), A => n13013, ZN => n13008);
   U5958 : OAI22_X1 port map( A1 => n16233, A2 => n15142, B1 => n16230, B2 => 
                           n14525, ZN => n13013);
   U5959 : AOI221_X1 port map( B1 => registers_47_23_port, B2 => n16290, C1 => 
                           registers_51_23_port, C2 => n16287, A => n12963, ZN 
                           => n12958);
   U5960 : OAI22_X1 port map( A1 => n16284, A2 => n15573, B1 => n16281, B2 => 
                           n14505, ZN => n12963);
   U5961 : AOI221_X1 port map( B1 => net227314, B2 => n16239, C1 => n16236, C2 
                           => datain(23), A => n12971, ZN => n12966);
   U5962 : OAI22_X1 port map( A1 => n16233, A2 => n15143, B1 => n16230, B2 => 
                           n14526, ZN => n12971);
   U5963 : AOI221_X1 port map( B1 => net226844, B2 => n16490, C1 => datain(0), 
                           C2 => n16487, A => n12491, ZN => n12484);
   U5964 : OAI22_X1 port map( A1 => n16484, A2 => n15123, B1 => n16481, B2 => 
                           n14506, ZN => n12491);
   U5965 : AOI221_X1 port map( B1 => net226857, B2 => n16490, C1 => datain(1), 
                           C2 => n16487, A => n12299, ZN => n12294);
   U5966 : OAI22_X1 port map( A1 => n16484, A2 => n15124, B1 => n16481, B2 => 
                           n14507, ZN => n12299);
   U5967 : AOI221_X1 port map( B1 => net226884, B2 => n16490, C1 => datain(2), 
                           C2 => n16487, A => n12146, ZN => n12141);
   U5968 : OAI22_X1 port map( A1 => n16484, A2 => n15125, B1 => n16481, B2 => 
                           n14508, ZN => n12146);
   U5969 : AOI221_X1 port map( B1 => net226904, B2 => n16490, C1 => datain(3), 
                           C2 => n16487, A => n11993, ZN => n11988);
   U5970 : OAI22_X1 port map( A1 => n16484, A2 => n14997, B1 => n16481, B2 => 
                           n14296, ZN => n11993);
   U5971 : AOI221_X1 port map( B1 => net226977, B2 => n16490, C1 => n16487, C2 
                           => datain(4), A => n11840, ZN => n11835);
   U5972 : OAI22_X1 port map( A1 => n16484, A2 => n14998, B1 => n16481, B2 => 
                           n14297, ZN => n11840);
   U5973 : AOI221_X1 port map( B1 => net226997, B2 => n16490, C1 => n16487, C2 
                           => datain(5), A => n11797, ZN => n11792);
   U5974 : OAI22_X1 port map( A1 => n16484, A2 => n14999, B1 => n16481, B2 => 
                           n14298, ZN => n11797);
   U5975 : AOI221_X1 port map( B1 => net227008, B2 => n16490, C1 => n16487, C2 
                           => datain(6), A => n11754, ZN => n11749);
   U5976 : OAI22_X1 port map( A1 => n16484, A2 => n15126, B1 => n16481, B2 => 
                           n14509, ZN => n11754);
   U5977 : AOI221_X1 port map( B1 => net227026, B2 => n16490, C1 => n16487, C2 
                           => datain(7), A => n11711, ZN => n11706);
   U5978 : OAI22_X1 port map( A1 => n16484, A2 => n15127, B1 => n16481, B2 => 
                           n14510, ZN => n11711);
   U5979 : AOI221_X1 port map( B1 => net227044, B2 => n16490, C1 => n16487, C2 
                           => datain(8), A => n11668, ZN => n11663);
   U5980 : OAI22_X1 port map( A1 => n16484, A2 => n15128, B1 => n16481, B2 => 
                           n14511, ZN => n11668);
   U5981 : AOI221_X1 port map( B1 => net227062, B2 => n16490, C1 => n16487, C2 
                           => datain(9), A => n11625, ZN => n11620);
   U5982 : OAI22_X1 port map( A1 => n16484, A2 => n15129, B1 => n16481, B2 => 
                           n14512, ZN => n11625);
   U5983 : AOI221_X1 port map( B1 => net227080, B2 => n16490, C1 => n16487, C2 
                           => datain(10), A => n11582, ZN => n11577);
   U5984 : OAI22_X1 port map( A1 => n16484, A2 => n15130, B1 => n16481, B2 => 
                           n14513, ZN => n11582);
   U5985 : AOI221_X1 port map( B1 => net227098, B2 => n16490, C1 => n16487, C2 
                           => datain(11), A => n11539, ZN => n11534);
   U5986 : OAI22_X1 port map( A1 => n16484, A2 => n15131, B1 => n16481, B2 => 
                           n14514, ZN => n11539);
   U5987 : AOI221_X1 port map( B1 => net227116, B2 => n16491, C1 => n16487, C2 
                           => datain(12), A => n11496, ZN => n11491);
   U5988 : OAI22_X1 port map( A1 => n16485, A2 => n15132, B1 => n16482, B2 => 
                           n14515, ZN => n11496);
   U5989 : AOI221_X1 port map( B1 => net227134, B2 => n16491, C1 => n16488, C2 
                           => datain(13), A => n11452, ZN => n11447);
   U5990 : OAI22_X1 port map( A1 => n16485, A2 => n15133, B1 => n16482, B2 => 
                           n14516, ZN => n11452);
   U5991 : AOI221_X1 port map( B1 => net227152, B2 => n16491, C1 => n16488, C2 
                           => datain(14), A => n11409, ZN => n11404);
   U5992 : OAI22_X1 port map( A1 => n16485, A2 => n15134, B1 => n16482, B2 => 
                           n14517, ZN => n11409);
   U5993 : AOI221_X1 port map( B1 => net227170, B2 => n16491, C1 => n16488, C2 
                           => datain(15), A => n11366, ZN => n11361);
   U5994 : OAI22_X1 port map( A1 => n16485, A2 => n15135, B1 => n16482, B2 => 
                           n14518, ZN => n11366);
   U5995 : AOI221_X1 port map( B1 => net227188, B2 => n16491, C1 => n16488, C2 
                           => datain(16), A => n11323, ZN => n11318);
   U5996 : OAI22_X1 port map( A1 => n16485, A2 => n15136, B1 => n16482, B2 => 
                           n14519, ZN => n11323);
   U5997 : AOI221_X1 port map( B1 => net227206, B2 => n16491, C1 => n16488, C2 
                           => datain(17), A => n11280, ZN => n11275);
   U5998 : OAI22_X1 port map( A1 => n16485, A2 => n15137, B1 => n16482, B2 => 
                           n14520, ZN => n11280);
   U5999 : AOI221_X1 port map( B1 => net227224, B2 => n16491, C1 => n16488, C2 
                           => datain(18), A => n11237, ZN => n11232);
   U6000 : OAI22_X1 port map( A1 => n16485, A2 => n15138, B1 => n16482, B2 => 
                           n14521, ZN => n11237);
   U6001 : AOI221_X1 port map( B1 => net227242, B2 => n16491, C1 => n16488, C2 
                           => datain(19), A => n11194, ZN => n11189);
   U6002 : OAI22_X1 port map( A1 => n16485, A2 => n15139, B1 => n16482, B2 => 
                           n14522, ZN => n11194);
   U6003 : AOI221_X1 port map( B1 => net227260, B2 => n16491, C1 => n16488, C2 
                           => datain(20), A => n11151, ZN => n11146);
   U6004 : OAI22_X1 port map( A1 => n16485, A2 => n15140, B1 => n16482, B2 => 
                           n14523, ZN => n11151);
   U6005 : AOI221_X1 port map( B1 => net227278, B2 => n16491, C1 => n16488, C2 
                           => datain(21), A => n11108, ZN => n11103);
   U6006 : OAI22_X1 port map( A1 => n16485, A2 => n15141, B1 => n16482, B2 => 
                           n14524, ZN => n11108);
   U6007 : AOI221_X1 port map( B1 => net227296, B2 => n16491, C1 => n16488, C2 
                           => datain(22), A => n11065, ZN => n11060);
   U6008 : OAI22_X1 port map( A1 => n16485, A2 => n15142, B1 => n16482, B2 => 
                           n14525, ZN => n11065);
   U6009 : AOI221_X1 port map( B1 => net227314, B2 => n16491, C1 => n16488, C2 
                           => datain(23), A => n11022, ZN => n11017);
   U6010 : OAI22_X1 port map( A1 => n16485, A2 => n15143, B1 => n16482, B2 => 
                           n14526, ZN => n11022);
   U6011 : AOI221_X1 port map( B1 => net226839, B2 => n17745, C1 => 
                           registers_29_0_port, C2 => n17742, A => n12389, ZN 
                           => n12384);
   U6012 : OAI22_X1 port map( A1 => n17739, A2 => n15736, B1 => n17736, B2 => 
                           n14771, ZN => n12389);
   U6013 : AOI221_X1 port map( B1 => registers_41_0_port, B2 => n17649, C1 => 
                           registers_40_0_port, C2 => n17646, A => n12405, ZN 
                           => n12400);
   U6014 : OAI22_X1 port map( A1 => n17643, A2 => n15466, B1 => n17640, B2 => 
                           n14772, ZN => n12405);
   U6015 : AOI221_X1 port map( B1 => registers_18_0_port, B2 => n17793, C1 => 
                           registers_19_0_port, C2 => n17790, A => n12381, ZN 
                           => n12376);
   U6016 : OAI22_X1 port map( A1 => n17787, A2 => n14605, B1 => n17784, B2 => 
                           n15292, ZN => n12381);
   U6017 : AOI221_X1 port map( B1 => net226861, B2 => n17745, C1 => 
                           registers_29_1_port, C2 => n17742, A => n12235, ZN 
                           => n12230);
   U6018 : OAI22_X1 port map( A1 => n17739, A2 => n15737, B1 => n17736, B2 => 
                           n14773, ZN => n12235);
   U6019 : AOI221_X1 port map( B1 => registers_41_1_port, B2 => n17649, C1 => 
                           registers_40_1_port, C2 => n17646, A => n12251, ZN 
                           => n12246);
   U6020 : OAI22_X1 port map( A1 => n17643, A2 => n15467, B1 => n17640, B2 => 
                           n14774, ZN => n12251);
   U6021 : AOI221_X1 port map( B1 => registers_18_1_port, B2 => n17793, C1 => 
                           registers_19_1_port, C2 => n17790, A => n12227, ZN 
                           => n12222);
   U6022 : OAI22_X1 port map( A1 => n17787, A2 => n14606, B1 => n17784, B2 => 
                           n15293, ZN => n12227);
   U6023 : AOI221_X1 port map( B1 => net226889, B2 => n17745, C1 => 
                           registers_29_2_port, C2 => n17742, A => n12080, ZN 
                           => n12075);
   U6024 : OAI22_X1 port map( A1 => n17739, A2 => n15738, B1 => n17736, B2 => 
                           n14775, ZN => n12080);
   U6025 : AOI221_X1 port map( B1 => registers_41_2_port, B2 => n17649, C1 => 
                           registers_40_2_port, C2 => n17646, A => n12096, ZN 
                           => n12091);
   U6026 : OAI22_X1 port map( A1 => n17643, A2 => n15468, B1 => n17640, B2 => 
                           n14776, ZN => n12096);
   U6027 : AOI221_X1 port map( B1 => registers_18_2_port, B2 => n17793, C1 => 
                           registers_19_2_port, C2 => n17790, A => n12072, ZN 
                           => n12067);
   U6028 : OAI22_X1 port map( A1 => n17787, A2 => n14607, B1 => n17784, B2 => 
                           n15294, ZN => n12072);
   U6029 : AOI221_X1 port map( B1 => net226909, B2 => n17745, C1 => 
                           registers_29_3_port, C2 => n17742, A => n11927, ZN 
                           => n11922);
   U6030 : OAI22_X1 port map( A1 => n17739, A2 => n15367, B1 => n17736, B2 => 
                           n14777, ZN => n11927);
   U6031 : AOI221_X1 port map( B1 => registers_41_3_port, B2 => n17649, C1 => 
                           registers_40_3_port, C2 => n17646, A => n11943, ZN 
                           => n11938);
   U6032 : OAI22_X1 port map( A1 => n17643, A2 => n15356, B1 => n17640, B2 => 
                           n14641, ZN => n11943);
   U6033 : AOI221_X1 port map( B1 => registers_18_3_port, B2 => n17793, C1 => 
                           registers_19_3_port, C2 => n17790, A => n11919, ZN 
                           => n11914);
   U6034 : OAI22_X1 port map( A1 => n17787, A2 => n14608, B1 => n17784, B2 => 
                           n15284, ZN => n11919);
   U6035 : AOI221_X1 port map( B1 => net226983, B2 => n17745, C1 => 
                           registers_29_4_port, C2 => n17742, A => n10484, ZN 
                           => n10479);
   U6036 : OAI22_X1 port map( A1 => n17739, A2 => n15368, B1 => n17736, B2 => 
                           n14778, ZN => n10484);
   U6037 : AOI221_X1 port map( B1 => registers_41_4_port, B2 => n17649, C1 => 
                           registers_40_4_port, C2 => n17646, A => n10500, ZN 
                           => n10495);
   U6038 : OAI22_X1 port map( A1 => n17643, A2 => n15469, B1 => n17640, B2 => 
                           n14779, ZN => n10500);
   U6039 : AOI221_X1 port map( B1 => registers_18_4_port, B2 => n17793, C1 => 
                           registers_19_4_port, C2 => n17790, A => n10476, ZN 
                           => n10471);
   U6040 : OAI22_X1 port map( A1 => n17787, A2 => n14569, B1 => n17784, B2 => 
                           n15295, ZN => n10476);
   U6041 : AOI221_X1 port map( B1 => net226992, B2 => n17745, C1 => 
                           registers_29_5_port, C2 => n17742, A => n10374, ZN 
                           => n10369);
   U6042 : OAI22_X1 port map( A1 => n17739, A2 => n15739, B1 => n17736, B2 => 
                           n14780, ZN => n10374);
   U6043 : AOI221_X1 port map( B1 => registers_41_5_port, B2 => n17649, C1 => 
                           registers_40_5_port, C2 => n17646, A => n10390, ZN 
                           => n10385);
   U6044 : OAI22_X1 port map( A1 => n17643, A2 => n15357, B1 => n17640, B2 => 
                           n14642, ZN => n10390);
   U6045 : AOI221_X1 port map( B1 => registers_18_5_port, B2 => n17793, C1 => 
                           registers_19_5_port, C2 => n17790, A => n10366, ZN 
                           => n10361);
   U6046 : OAI22_X1 port map( A1 => n17787, A2 => n14609, B1 => n17784, B2 => 
                           n15296, ZN => n10366);
   U6047 : AOI221_X1 port map( B1 => net227016, B2 => n17745, C1 => 
                           registers_29_6_port, C2 => n17742, A => n10262, ZN 
                           => n10257);
   U6048 : OAI22_X1 port map( A1 => n17739, A2 => n15740, B1 => n17736, B2 => 
                           n14781, ZN => n10262);
   U6049 : AOI221_X1 port map( B1 => registers_41_6_port, B2 => n17649, C1 => 
                           registers_40_6_port, C2 => n17646, A => n10278, ZN 
                           => n10273);
   U6050 : OAI22_X1 port map( A1 => n17643, A2 => n15470, B1 => n17640, B2 => 
                           n14782, ZN => n10278);
   U6051 : AOI221_X1 port map( B1 => registers_18_6_port, B2 => n17793, C1 => 
                           registers_19_6_port, C2 => n17790, A => n10254, ZN 
                           => n10249);
   U6052 : OAI22_X1 port map( A1 => n17787, A2 => n14610, B1 => n17784, B2 => 
                           n15297, ZN => n10254);
   U6053 : AOI221_X1 port map( B1 => net227034, B2 => n17745, C1 => 
                           registers_29_7_port, C2 => n17742, A => n7626, ZN =>
                           n7621);
   U6054 : OAI22_X1 port map( A1 => n17739, A2 => n15741, B1 => n17736, B2 => 
                           n14783, ZN => n7626);
   U6055 : AOI221_X1 port map( B1 => registers_41_7_port, B2 => n17649, C1 => 
                           registers_40_7_port, C2 => n17646, A => n7642, ZN =>
                           n7637);
   U6056 : OAI22_X1 port map( A1 => n17643, A2 => n15471, B1 => n17640, B2 => 
                           n14784, ZN => n7642);
   U6057 : AOI221_X1 port map( B1 => registers_18_7_port, B2 => n17793, C1 => 
                           registers_19_7_port, C2 => n17790, A => n7618, ZN =>
                           n7613);
   U6058 : OAI22_X1 port map( A1 => n17787, A2 => n14611, B1 => n17784, B2 => 
                           n15298, ZN => n7618);
   U6059 : AOI221_X1 port map( B1 => net227052, B2 => n17745, C1 => 
                           registers_29_8_port, C2 => n17742, A => n7511, ZN =>
                           n7506);
   U6060 : OAI22_X1 port map( A1 => n17739, A2 => n15742, B1 => n17736, B2 => 
                           n14785, ZN => n7511);
   U6061 : AOI221_X1 port map( B1 => registers_41_8_port, B2 => n17649, C1 => 
                           registers_40_8_port, C2 => n17646, A => n7527, ZN =>
                           n7522);
   U6062 : OAI22_X1 port map( A1 => n17643, A2 => n15472, B1 => n17640, B2 => 
                           n14786, ZN => n7527);
   U6063 : AOI221_X1 port map( B1 => registers_18_8_port, B2 => n17793, C1 => 
                           registers_19_8_port, C2 => n17790, A => n7503, ZN =>
                           n7498);
   U6064 : OAI22_X1 port map( A1 => n17787, A2 => n14612, B1 => n17784, B2 => 
                           n15299, ZN => n7503);
   U6065 : AOI221_X1 port map( B1 => net227070, B2 => n17745, C1 => 
                           registers_29_9_port, C2 => n17742, A => n7402, ZN =>
                           n7397);
   U6066 : OAI22_X1 port map( A1 => n17739, A2 => n15743, B1 => n17736, B2 => 
                           n14787, ZN => n7402);
   U6067 : AOI221_X1 port map( B1 => registers_41_9_port, B2 => n17649, C1 => 
                           registers_40_9_port, C2 => n17646, A => n7418, ZN =>
                           n7413);
   U6068 : OAI22_X1 port map( A1 => n17643, A2 => n15473, B1 => n17640, B2 => 
                           n14788, ZN => n7418);
   U6069 : AOI221_X1 port map( B1 => registers_18_9_port, B2 => n17793, C1 => 
                           registers_19_9_port, C2 => n17790, A => n7394, ZN =>
                           n7389);
   U6070 : OAI22_X1 port map( A1 => n17787, A2 => n14613, B1 => n17784, B2 => 
                           n15300, ZN => n7394);
   U6071 : AOI221_X1 port map( B1 => net227088, B2 => n17745, C1 => 
                           registers_29_10_port, C2 => n17742, A => n7293, ZN 
                           => n7288);
   U6072 : OAI22_X1 port map( A1 => n17739, A2 => n15744, B1 => n17736, B2 => 
                           n14789, ZN => n7293);
   U6073 : AOI221_X1 port map( B1 => registers_41_10_port, B2 => n17649, C1 => 
                           registers_40_10_port, C2 => n17646, A => n7309, ZN 
                           => n7304);
   U6074 : OAI22_X1 port map( A1 => n17643, A2 => n15474, B1 => n17640, B2 => 
                           n14790, ZN => n7309);
   U6075 : AOI221_X1 port map( B1 => registers_18_10_port, B2 => n17793, C1 => 
                           registers_19_10_port, C2 => n17790, A => n7285, ZN 
                           => n7280);
   U6076 : OAI22_X1 port map( A1 => n17787, A2 => n14614, B1 => n17784, B2 => 
                           n15301, ZN => n7285);
   U6077 : AOI221_X1 port map( B1 => net227106, B2 => n17746, C1 => 
                           registers_29_11_port, C2 => n17743, A => n7179, ZN 
                           => n7174);
   U6078 : OAI22_X1 port map( A1 => n17740, A2 => n15745, B1 => n17737, B2 => 
                           n14791, ZN => n7179);
   U6079 : AOI221_X1 port map( B1 => registers_41_11_port, B2 => n17650, C1 => 
                           registers_40_11_port, C2 => n17647, A => n7195, ZN 
                           => n7190);
   U6080 : OAI22_X1 port map( A1 => n17644, A2 => n15475, B1 => n17641, B2 => 
                           n14792, ZN => n7195);
   U6081 : AOI221_X1 port map( B1 => registers_18_11_port, B2 => n17794, C1 => 
                           registers_19_11_port, C2 => n17791, A => n7171, ZN 
                           => n7166);
   U6082 : OAI22_X1 port map( A1 => n17788, A2 => n14615, B1 => n17785, B2 => 
                           n15302, ZN => n7171);
   U6083 : AOI221_X1 port map( B1 => net227124, B2 => n17746, C1 => 
                           registers_29_12_port, C2 => n17743, A => n7070, ZN 
                           => n7065);
   U6084 : OAI22_X1 port map( A1 => n17740, A2 => n15746, B1 => n17737, B2 => 
                           n14793, ZN => n7070);
   U6085 : AOI221_X1 port map( B1 => registers_41_12_port, B2 => n17650, C1 => 
                           registers_40_12_port, C2 => n17647, A => n7086, ZN 
                           => n7081);
   U6086 : OAI22_X1 port map( A1 => n17644, A2 => n15476, B1 => n17641, B2 => 
                           n14794, ZN => n7086);
   U6087 : AOI221_X1 port map( B1 => registers_18_12_port, B2 => n17794, C1 => 
                           registers_19_12_port, C2 => n17791, A => n7062, ZN 
                           => n7057);
   U6088 : OAI22_X1 port map( A1 => n17788, A2 => n14616, B1 => n17785, B2 => 
                           n15303, ZN => n7062);
   U6089 : AOI221_X1 port map( B1 => net227142, B2 => n17746, C1 => 
                           registers_29_13_port, C2 => n17743, A => n6961, ZN 
                           => n6956);
   U6090 : OAI22_X1 port map( A1 => n17740, A2 => n15747, B1 => n17737, B2 => 
                           n14795, ZN => n6961);
   U6091 : AOI221_X1 port map( B1 => registers_41_13_port, B2 => n17650, C1 => 
                           registers_40_13_port, C2 => n17647, A => n6977, ZN 
                           => n6972);
   U6092 : OAI22_X1 port map( A1 => n17644, A2 => n15477, B1 => n17641, B2 => 
                           n14796, ZN => n6977);
   U6093 : AOI221_X1 port map( B1 => registers_18_13_port, B2 => n17794, C1 => 
                           registers_19_13_port, C2 => n17791, A => n6953, ZN 
                           => n6948);
   U6094 : OAI22_X1 port map( A1 => n17788, A2 => n14617, B1 => n17785, B2 => 
                           n15304, ZN => n6953);
   U6095 : AOI221_X1 port map( B1 => net227160, B2 => n17746, C1 => 
                           registers_29_14_port, C2 => n17743, A => n6852, ZN 
                           => n6847);
   U6096 : OAI22_X1 port map( A1 => n17740, A2 => n15748, B1 => n17737, B2 => 
                           n14797, ZN => n6852);
   U6097 : AOI221_X1 port map( B1 => registers_41_14_port, B2 => n17650, C1 => 
                           registers_40_14_port, C2 => n17647, A => n6868, ZN 
                           => n6863);
   U6098 : OAI22_X1 port map( A1 => n17644, A2 => n15478, B1 => n17641, B2 => 
                           n14798, ZN => n6868);
   U6099 : AOI221_X1 port map( B1 => registers_18_14_port, B2 => n17794, C1 => 
                           registers_19_14_port, C2 => n17791, A => n6844, ZN 
                           => n6839);
   U6100 : OAI22_X1 port map( A1 => n17788, A2 => n14618, B1 => n17785, B2 => 
                           n15305, ZN => n6844);
   U6101 : AOI221_X1 port map( B1 => net227178, B2 => n17746, C1 => 
                           registers_29_15_port, C2 => n17743, A => n6743, ZN 
                           => n6738);
   U6102 : OAI22_X1 port map( A1 => n17740, A2 => n15749, B1 => n17737, B2 => 
                           n14799, ZN => n6743);
   U6103 : AOI221_X1 port map( B1 => registers_41_15_port, B2 => n17650, C1 => 
                           registers_40_15_port, C2 => n17647, A => n6759, ZN 
                           => n6754);
   U6104 : OAI22_X1 port map( A1 => n17644, A2 => n15479, B1 => n17641, B2 => 
                           n14800, ZN => n6759);
   U6105 : AOI221_X1 port map( B1 => registers_18_15_port, B2 => n17794, C1 => 
                           registers_19_15_port, C2 => n17791, A => n6735, ZN 
                           => n6730);
   U6106 : OAI22_X1 port map( A1 => n17788, A2 => n14619, B1 => n17785, B2 => 
                           n15306, ZN => n6735);
   U6107 : AOI221_X1 port map( B1 => net227196, B2 => n17746, C1 => 
                           registers_29_16_port, C2 => n17743, A => n6600, ZN 
                           => n6580);
   U6108 : OAI22_X1 port map( A1 => n17740, A2 => n15750, B1 => n17737, B2 => 
                           n14801, ZN => n6600);
   U6109 : AOI221_X1 port map( B1 => registers_41_16_port, B2 => n17650, C1 => 
                           registers_40_16_port, C2 => n17647, A => n6619, ZN 
                           => n6614);
   U6110 : OAI22_X1 port map( A1 => n17644, A2 => n15480, B1 => n17641, B2 => 
                           n14802, ZN => n6619);
   U6111 : AOI221_X1 port map( B1 => registers_18_16_port, B2 => n17794, C1 => 
                           registers_19_16_port, C2 => n17791, A => n6575, ZN 
                           => n6568);
   U6112 : OAI22_X1 port map( A1 => n17788, A2 => n14620, B1 => n17785, B2 => 
                           n15307, ZN => n6575);
   U6113 : AOI221_X1 port map( B1 => net227214, B2 => n17746, C1 => 
                           registers_29_17_port, C2 => n17743, A => n6413, ZN 
                           => n6393);
   U6114 : OAI22_X1 port map( A1 => n17740, A2 => n15751, B1 => n17737, B2 => 
                           n14803, ZN => n6413);
   U6115 : AOI221_X1 port map( B1 => registers_41_17_port, B2 => n17650, C1 => 
                           registers_40_17_port, C2 => n17647, A => n6434, ZN 
                           => n6427);
   U6116 : OAI22_X1 port map( A1 => n17644, A2 => n15481, B1 => n17641, B2 => 
                           n14804, ZN => n6434);
   U6117 : AOI221_X1 port map( B1 => registers_18_17_port, B2 => n17794, C1 => 
                           registers_19_17_port, C2 => n17791, A => n6388, ZN 
                           => n6383);
   U6118 : OAI22_X1 port map( A1 => n17788, A2 => n14621, B1 => n17785, B2 => 
                           n15308, ZN => n6388);
   U6119 : AOI221_X1 port map( B1 => net227232, B2 => n17746, C1 => 
                           registers_29_18_port, C2 => n17743, A => n6226, ZN 
                           => n6221);
   U6120 : OAI22_X1 port map( A1 => n17740, A2 => n15752, B1 => n17737, B2 => 
                           n14805, ZN => n6226);
   U6121 : AOI221_X1 port map( B1 => registers_41_18_port, B2 => n17650, C1 => 
                           registers_40_18_port, C2 => n17647, A => n6248, ZN 
                           => n6240);
   U6122 : OAI22_X1 port map( A1 => n17644, A2 => n15482, B1 => n17641, B2 => 
                           n14806, ZN => n6248);
   U6123 : AOI221_X1 port map( B1 => registers_18_18_port, B2 => n17794, C1 => 
                           registers_19_18_port, C2 => n17791, A => n6203, ZN 
                           => n6196);
   U6124 : OAI22_X1 port map( A1 => n17788, A2 => n14622, B1 => n17785, B2 => 
                           n15309, ZN => n6203);
   U6125 : AOI221_X1 port map( B1 => net227250, B2 => n17746, C1 => 
                           registers_29_19_port, C2 => n17743, A => n6039, ZN 
                           => n6034);
   U6126 : OAI22_X1 port map( A1 => n17740, A2 => n15753, B1 => n17737, B2 => 
                           n14807, ZN => n6039);
   U6127 : AOI221_X1 port map( B1 => registers_41_19_port, B2 => n17650, C1 => 
                           registers_40_19_port, C2 => n17647, A => n6061, ZN 
                           => n6055);
   U6128 : OAI22_X1 port map( A1 => n17644, A2 => n15483, B1 => n17641, B2 => 
                           n14808, ZN => n6061);
   U6129 : AOI221_X1 port map( B1 => registers_18_19_port, B2 => n17794, C1 => 
                           registers_19_19_port, C2 => n17791, A => n6031, ZN 
                           => n6009);
   U6130 : OAI22_X1 port map( A1 => n17788, A2 => n14623, B1 => n17785, B2 => 
                           n15310, ZN => n6031);
   U6131 : AOI221_X1 port map( B1 => net227268, B2 => n17746, C1 => 
                           registers_29_20_port, C2 => n17743, A => n5853, ZN 
                           => n5847);
   U6132 : OAI22_X1 port map( A1 => n17740, A2 => n15754, B1 => n17737, B2 => 
                           n14809, ZN => n5853);
   U6133 : AOI221_X1 port map( B1 => registers_41_20_port, B2 => n17650, C1 => 
                           registers_40_20_port, C2 => n17647, A => n5875, ZN 
                           => n5869);
   U6134 : OAI22_X1 port map( A1 => n17644, A2 => n15484, B1 => n17641, B2 => 
                           n14810, ZN => n5875);
   U6135 : AOI221_X1 port map( B1 => registers_18_20_port, B2 => n17794, C1 => 
                           registers_19_20_port, C2 => n17791, A => n5844, ZN 
                           => n5824);
   U6136 : OAI22_X1 port map( A1 => n17788, A2 => n14624, B1 => n17785, B2 => 
                           n15311, ZN => n5844);
   U6137 : AOI221_X1 port map( B1 => net227286, B2 => n17746, C1 => 
                           registers_29_21_port, C2 => n17743, A => n5667, ZN 
                           => n5660);
   U6138 : OAI22_X1 port map( A1 => n17740, A2 => n15755, B1 => n17737, B2 => 
                           n14811, ZN => n5667);
   U6139 : AOI221_X1 port map( B1 => registers_41_21_port, B2 => n17650, C1 => 
                           registers_40_21_port, C2 => n17647, A => n5690, ZN 
                           => n5682);
   U6140 : OAI22_X1 port map( A1 => n17644, A2 => n15485, B1 => n17641, B2 => 
                           n14812, ZN => n5690);
   U6141 : AOI221_X1 port map( B1 => registers_18_21_port, B2 => n17794, C1 => 
                           registers_19_21_port, C2 => n17791, A => n5657, ZN 
                           => n5637);
   U6142 : OAI22_X1 port map( A1 => n17788, A2 => n14625, B1 => n17785, B2 => 
                           n15312, ZN => n5657);
   U6143 : AOI221_X1 port map( B1 => net227304, B2 => n17746, C1 => 
                           registers_29_22_port, C2 => n17743, A => n5481, ZN 
                           => n5473);
   U6144 : OAI22_X1 port map( A1 => n17740, A2 => n15756, B1 => n17737, B2 => 
                           n14813, ZN => n5481);
   U6145 : AOI221_X1 port map( B1 => registers_41_22_port, B2 => n17650, C1 => 
                           registers_40_22_port, C2 => n17647, A => n5503, ZN 
                           => n5495);
   U6146 : OAI22_X1 port map( A1 => n17644, A2 => n15486, B1 => n17641, B2 => 
                           n14814, ZN => n5503);
   U6147 : AOI221_X1 port map( B1 => registers_18_22_port, B2 => n17794, C1 => 
                           registers_19_22_port, C2 => n17791, A => n5470, ZN 
                           => n5465);
   U6148 : OAI22_X1 port map( A1 => n17788, A2 => n14626, B1 => n17785, B2 => 
                           n15313, ZN => n5470);
   U6149 : AOI221_X1 port map( B1 => net227466, B2 => n17745, C1 => 
                           registers_29_31_port, C2 => n17742, A => n14139, ZN 
                           => n14110);
   U6150 : OAI22_X1 port map( A1 => n17739, A2 => n15757, B1 => n17736, B2 => 
                           n14815, ZN => n14139);
   U6151 : AOI221_X1 port map( B1 => registers_41_31_port, B2 => n17649, C1 => 
                           registers_40_31_port, C2 => n17646, A => n14203, ZN 
                           => n14188);
   U6152 : OAI22_X1 port map( A1 => n17643, A2 => n15487, B1 => n17640, B2 => 
                           n14816, ZN => n14203);
   U6153 : AOI221_X1 port map( B1 => registers_18_31_port, B2 => n17793, C1 => 
                           registers_19_31_port, C2 => n17790, A => n14102, ZN 
                           => n14081);
   U6154 : OAI22_X1 port map( A1 => n17787, A2 => n14627, B1 => n17784, B2 => 
                           n15314, ZN => n14102);
   U6155 : AOI221_X1 port map( B1 => registers_50_24_port, B2 => n16279, C1 => 
                           net227335, C2 => n16276, A => n12922, ZN => n12915);
   U6156 : OAI22_X1 port map( A1 => n16273, A2 => n12349, B1 => n16270, B2 => 
                           n14931, ZN => n12922);
   U6157 : AOI221_X1 port map( B1 => registers_50_25_port, B2 => n16279, C1 => 
                           net227353, C2 => n16276, A => n12880, ZN => n12873);
   U6158 : OAI22_X1 port map( A1 => n16273, A2 => n12350, B1 => n16270, B2 => 
                           n14932, ZN => n12880);
   U6159 : AOI221_X1 port map( B1 => registers_50_26_port, B2 => n16279, C1 => 
                           net227371, C2 => n16276, A => n12838, ZN => n12831);
   U6160 : OAI22_X1 port map( A1 => n16273, A2 => n12351, B1 => n16270, B2 => 
                           n14933, ZN => n12838);
   U6161 : AOI221_X1 port map( B1 => registers_50_27_port, B2 => n16279, C1 => 
                           net227389, C2 => n16276, A => n12796, ZN => n12789);
   U6162 : OAI22_X1 port map( A1 => n16273, A2 => n12352, B1 => n16270, B2 => 
                           n14934, ZN => n12796);
   U6163 : AOI221_X1 port map( B1 => registers_50_28_port, B2 => n16279, C1 => 
                           net227407, C2 => n16276, A => n12754, ZN => n12747);
   U6164 : OAI22_X1 port map( A1 => n16273, A2 => n12353, B1 => n16270, B2 => 
                           n14935, ZN => n12754);
   U6165 : AOI221_X1 port map( B1 => registers_50_29_port, B2 => n16279, C1 => 
                           net227425, C2 => n16276, A => n12712, ZN => n12705);
   U6166 : OAI22_X1 port map( A1 => n16273, A2 => n12354, B1 => n16270, B2 => 
                           n14936, ZN => n12712);
   U6167 : AOI221_X1 port map( B1 => registers_50_30_port, B2 => n16279, C1 => 
                           net227443, C2 => n16276, A => n12670, ZN => n12662);
   U6168 : OAI22_X1 port map( A1 => n16273, A2 => n12197, B1 => n16270, B2 => 
                           n14855, ZN => n12670);
   U6169 : AOI221_X1 port map( B1 => registers_50_31_port, B2 => n16279, C1 => 
                           net227461, C2 => n16276, A => n12605, ZN => n12582);
   U6170 : OAI22_X1 port map( A1 => n16273, A2 => n12355, B1 => n16270, B2 => 
                           n14937, ZN => n12605);
   U6171 : AOI221_X1 port map( B1 => registers_50_24_port, B2 => n16531, C1 => 
                           net227335, C2 => n16528, A => n10972, ZN => n10965);
   U6172 : OAI22_X1 port map( A1 => n16525, A2 => n12349, B1 => n16522, B2 => 
                           n14931, ZN => n10972);
   U6173 : AOI221_X1 port map( B1 => registers_7_24_port, B2 => n16480, C1 => 
                           registers_42_24_port, C2 => n16477, A => n10980, ZN 
                           => n10973);
   U6174 : OAI22_X1 port map( A1 => n16474, A2 => n15233, B1 => n16471, B2 => 
                           n14352, ZN => n10980);
   U6175 : AOI221_X1 port map( B1 => registers_50_25_port, B2 => n16531, C1 => 
                           net227353, C2 => n16528, A => n10929, ZN => n10922);
   U6176 : OAI22_X1 port map( A1 => n16525, A2 => n12350, B1 => n16522, B2 => 
                           n14932, ZN => n10929);
   U6177 : AOI221_X1 port map( B1 => registers_7_25_port, B2 => n16480, C1 => 
                           registers_42_25_port, C2 => n16477, A => n10937, ZN 
                           => n10930);
   U6178 : OAI22_X1 port map( A1 => n16474, A2 => n15234, B1 => n16471, B2 => 
                           n14353, ZN => n10937);
   U6179 : AOI221_X1 port map( B1 => registers_50_26_port, B2 => n16531, C1 => 
                           net227371, C2 => n16528, A => n10886, ZN => n10879);
   U6180 : OAI22_X1 port map( A1 => n16525, A2 => n12351, B1 => n16522, B2 => 
                           n14933, ZN => n10886);
   U6181 : AOI221_X1 port map( B1 => registers_7_26_port, B2 => n16480, C1 => 
                           registers_42_26_port, C2 => n16477, A => n10894, ZN 
                           => n10887);
   U6182 : OAI22_X1 port map( A1 => n16474, A2 => n15235, B1 => n16471, B2 => 
                           n14354, ZN => n10894);
   U6183 : AOI221_X1 port map( B1 => registers_50_27_port, B2 => n16531, C1 => 
                           net227389, C2 => n16528, A => n10843, ZN => n10836);
   U6184 : OAI22_X1 port map( A1 => n16525, A2 => n12352, B1 => n16522, B2 => 
                           n14934, ZN => n10843);
   U6185 : AOI221_X1 port map( B1 => registers_7_27_port, B2 => n16480, C1 => 
                           registers_42_27_port, C2 => n16477, A => n10851, ZN 
                           => n10844);
   U6186 : OAI22_X1 port map( A1 => n16474, A2 => n15236, B1 => n16471, B2 => 
                           n14355, ZN => n10851);
   U6187 : AOI221_X1 port map( B1 => registers_50_28_port, B2 => n16531, C1 => 
                           net227407, C2 => n16528, A => n10800, ZN => n10793);
   U6188 : OAI22_X1 port map( A1 => n16525, A2 => n12353, B1 => n16522, B2 => 
                           n14935, ZN => n10800);
   U6189 : AOI221_X1 port map( B1 => registers_7_28_port, B2 => n16480, C1 => 
                           registers_42_28_port, C2 => n16477, A => n10808, ZN 
                           => n10801);
   U6190 : OAI22_X1 port map( A1 => n16474, A2 => n15237, B1 => n16471, B2 => 
                           n14356, ZN => n10808);
   U6191 : AOI221_X1 port map( B1 => registers_50_29_port, B2 => n16531, C1 => 
                           net227425, C2 => n16528, A => n10757, ZN => n10750);
   U6192 : OAI22_X1 port map( A1 => n16525, A2 => n12354, B1 => n16522, B2 => 
                           n14936, ZN => n10757);
   U6193 : AOI221_X1 port map( B1 => registers_7_29_port, B2 => n16480, C1 => 
                           registers_42_29_port, C2 => n16477, A => n10765, ZN 
                           => n10758);
   U6194 : OAI22_X1 port map( A1 => n16474, A2 => n15238, B1 => n16471, B2 => 
                           n14357, ZN => n10765);
   U6195 : AOI221_X1 port map( B1 => registers_50_30_port, B2 => n16531, C1 => 
                           net227443, C2 => n16528, A => n10711, ZN => n10700);
   U6196 : OAI22_X1 port map( A1 => n16525, A2 => n12197, B1 => n16522, B2 => 
                           n14855, ZN => n10711);
   U6197 : AOI221_X1 port map( B1 => registers_7_30_port, B2 => n16480, C1 => 
                           registers_42_30_port, C2 => n16477, A => n10720, ZN 
                           => n10713);
   U6198 : OAI22_X1 port map( A1 => n16474, A2 => n14874, B1 => n16471, B2 => 
                           n14055, ZN => n10720);
   U6199 : AOI221_X1 port map( B1 => registers_50_31_port, B2 => n16531, C1 => 
                           net227461, C2 => n16528, A => n10623, ZN => n10596);
   U6200 : OAI22_X1 port map( A1 => n16525, A2 => n12355, B1 => n16522, B2 => 
                           n14937, ZN => n10623);
   U6201 : AOI221_X1 port map( B1 => registers_7_31_port, B2 => n16480, C1 => 
                           registers_42_31_port, C2 => n16477, A => n10657, ZN 
                           => n10628);
   U6202 : OAI22_X1 port map( A1 => n16474, A2 => n15239, B1 => n16471, B2 => 
                           n14358, ZN => n10657);
   U6203 : AOI221_X1 port map( B1 => registers_48_23_port, B2 => n17639, C1 => 
                           registers_4_23_port, C2 => n17636, A => n5319, ZN =>
                           n5309);
   U6204 : OAI22_X1 port map( A1 => n17633, A2 => n15488, B1 => n17630, B2 => 
                           n14671, ZN => n5319);
   U6205 : AOI221_X1 port map( B1 => registers_23_23_port, B2 => n17783, C1 => 
                           registers_22_23_port, C2 => n17780, A => n5285, ZN 
                           => n5277);
   U6206 : OAI22_X1 port map( A1 => n17777, A2 => n12198, B1 => n17774, B2 => 
                           n14824, ZN => n5285);
   U6207 : AOI221_X1 port map( B1 => registers_48_24_port, B2 => n17639, C1 => 
                           registers_4_24_port, C2 => n17636, A => n5147, ZN =>
                           n5138);
   U6208 : OAI22_X1 port map( A1 => n17633, A2 => n15489, B1 => n17630, B2 => 
                           n14672, ZN => n5147);
   U6209 : AOI221_X1 port map( B1 => registers_23_24_port, B2 => n17783, C1 => 
                           registers_22_24_port, C2 => n17780, A => n5119, ZN 
                           => n5111);
   U6210 : OAI22_X1 port map( A1 => n17777, A2 => n12199, B1 => n17774, B2 => 
                           n14825, ZN => n5119);
   U6211 : AOI221_X1 port map( B1 => registers_48_25_port, B2 => n17639, C1 => 
                           registers_4_25_port, C2 => n17636, A => n5031, ZN =>
                           n5024);
   U6212 : OAI22_X1 port map( A1 => n17633, A2 => n15490, B1 => n17630, B2 => 
                           n14673, ZN => n5031);
   U6213 : AOI221_X1 port map( B1 => registers_23_25_port, B2 => n17783, C1 => 
                           registers_22_25_port, C2 => n17780, A => n5005, ZN 
                           => n4998);
   U6214 : OAI22_X1 port map( A1 => n17777, A2 => n12200, B1 => n17774, B2 => 
                           n14826, ZN => n5005);
   U6215 : AOI221_X1 port map( B1 => registers_48_26_port, B2 => n17639, C1 => 
                           registers_4_26_port, C2 => n17636, A => n4913, ZN =>
                           n4906);
   U6216 : OAI22_X1 port map( A1 => n17633, A2 => n15491, B1 => n17630, B2 => 
                           n14674, ZN => n4913);
   U6217 : AOI221_X1 port map( B1 => registers_23_26_port, B2 => n17783, C1 => 
                           registers_22_26_port, C2 => n17780, A => n4883, ZN 
                           => n4876);
   U6218 : OAI22_X1 port map( A1 => n17777, A2 => n12201, B1 => n17774, B2 => 
                           n14827, ZN => n4883);
   U6219 : AOI221_X1 port map( B1 => registers_48_27_port, B2 => n17639, C1 => 
                           registers_4_27_port, C2 => n17636, A => n4782, ZN =>
                           n4775);
   U6220 : OAI22_X1 port map( A1 => n17633, A2 => n15492, B1 => n17630, B2 => 
                           n14675, ZN => n4782);
   U6221 : AOI221_X1 port map( B1 => registers_23_27_port, B2 => n17783, C1 => 
                           registers_22_27_port, C2 => n17780, A => n4756, ZN 
                           => n4745);
   U6222 : OAI22_X1 port map( A1 => n17777, A2 => n12202, B1 => n17774, B2 => 
                           n14828, ZN => n4756);
   U6223 : AOI221_X1 port map( B1 => registers_48_28_port, B2 => n17639, C1 => 
                           registers_4_28_port, C2 => n17636, A => n4653, ZN =>
                           n4642);
   U6224 : OAI22_X1 port map( A1 => n17633, A2 => n15493, B1 => n17630, B2 => 
                           n14676, ZN => n4653);
   U6225 : AOI221_X1 port map( B1 => registers_23_28_port, B2 => n17783, C1 => 
                           registers_22_28_port, C2 => n17780, A => n4625, ZN 
                           => n4618);
   U6226 : OAI22_X1 port map( A1 => n17777, A2 => n12203, B1 => n17774, B2 => 
                           n14829, ZN => n4625);
   U6227 : AOI221_X1 port map( B1 => registers_48_29_port, B2 => n17639, C1 => 
                           registers_4_29_port, C2 => n17636, A => n4524, ZN =>
                           n4517);
   U6228 : OAI22_X1 port map( A1 => n17633, A2 => n15494, B1 => n17630, B2 => 
                           n14677, ZN => n4524);
   U6229 : AOI221_X1 port map( B1 => registers_23_29_port, B2 => n17783, C1 => 
                           registers_22_29_port, C2 => n17780, A => n4492, ZN 
                           => n4485);
   U6230 : OAI22_X1 port map( A1 => n17777, A2 => n12204, B1 => n17774, B2 => 
                           n14830, ZN => n4492);
   U6231 : AOI221_X1 port map( B1 => registers_48_30_port, B2 => n17639, C1 => 
                           registers_4_30_port, C2 => n17636, A => n4241, ZN =>
                           n4213);
   U6232 : OAI22_X1 port map( A1 => n17633, A2 => n15276, B1 => n17630, B2 => 
                           n14628, ZN => n4241);
   U6233 : AOI221_X1 port map( B1 => registers_23_30_port, B2 => n17783, C1 => 
                           registers_22_30_port, C2 => n17780, A => n4132, ZN 
                           => n4101);
   U6234 : OAI22_X1 port map( A1 => n17777, A2 => n12161, B1 => n17774, B2 => 
                           n14822, ZN => n4132);
   U6235 : AOI221_X1 port map( B1 => registers_7_0_port, B2 => n16226, C1 => 
                           registers_42_0_port, C2 => n16223, A => n13977, ZN 
                           => n13964);
   U6236 : OAI22_X1 port map( A1 => n16220, A2 => n15210, B1 => n16217, B2 => 
                           n14329, ZN => n13977);
   U6237 : AOI221_X1 port map( B1 => registers_7_1_port, B2 => n16226, C1 => 
                           registers_42_1_port, C2 => n16223, A => n13896, ZN 
                           => n13889);
   U6238 : OAI22_X1 port map( A1 => n16220, A2 => n15211, B1 => n16217, B2 => 
                           n14330, ZN => n13896);
   U6239 : AOI221_X1 port map( B1 => registers_7_2_port, B2 => n16226, C1 => 
                           registers_42_2_port, C2 => n16223, A => n13854, ZN 
                           => n13847);
   U6240 : OAI22_X1 port map( A1 => n16220, A2 => n15212, B1 => n16217, B2 => 
                           n14331, ZN => n13854);
   U6241 : AOI221_X1 port map( B1 => registers_7_3_port, B2 => n16226, C1 => 
                           registers_42_3_port, C2 => n16223, A => n13812, ZN 
                           => n13805);
   U6242 : OAI22_X1 port map( A1 => n16220, A2 => n15003, B1 => n16217, B2 => 
                           n14288, ZN => n13812);
   U6243 : AOI221_X1 port map( B1 => registers_7_4_port, B2 => n16226, C1 => 
                           registers_42_4_port, C2 => n16223, A => n13770, ZN 
                           => n13763);
   U6244 : OAI22_X1 port map( A1 => n16220, A2 => n15213, B1 => n16217, B2 => 
                           n14332, ZN => n13770);
   U6245 : AOI221_X1 port map( B1 => registers_7_5_port, B2 => n16226, C1 => 
                           registers_42_5_port, C2 => n16223, A => n13728, ZN 
                           => n13721);
   U6246 : OAI22_X1 port map( A1 => n16220, A2 => n15214, B1 => n16217, B2 => 
                           n14333, ZN => n13728);
   U6247 : AOI221_X1 port map( B1 => registers_7_6_port, B2 => n16226, C1 => 
                           registers_42_6_port, C2 => n16223, A => n13686, ZN 
                           => n13679);
   U6248 : OAI22_X1 port map( A1 => n16220, A2 => n15215, B1 => n16217, B2 => 
                           n14334, ZN => n13686);
   U6249 : AOI221_X1 port map( B1 => registers_7_7_port, B2 => n16226, C1 => 
                           registers_42_7_port, C2 => n16223, A => n13644, ZN 
                           => n13637);
   U6250 : OAI22_X1 port map( A1 => n16220, A2 => n15216, B1 => n16217, B2 => 
                           n14335, ZN => n13644);
   U6251 : AOI221_X1 port map( B1 => registers_7_8_port, B2 => n16226, C1 => 
                           registers_42_8_port, C2 => n16223, A => n13602, ZN 
                           => n13595);
   U6252 : OAI22_X1 port map( A1 => n16220, A2 => n15217, B1 => n16217, B2 => 
                           n14336, ZN => n13602);
   U6253 : AOI221_X1 port map( B1 => registers_7_9_port, B2 => n16226, C1 => 
                           registers_42_9_port, C2 => n16223, A => n13560, ZN 
                           => n13553);
   U6254 : OAI22_X1 port map( A1 => n16220, A2 => n15218, B1 => n16217, B2 => 
                           n14337, ZN => n13560);
   U6255 : AOI221_X1 port map( B1 => registers_7_10_port, B2 => n16226, C1 => 
                           registers_42_10_port, C2 => n16223, A => n13518, ZN 
                           => n13511);
   U6256 : OAI22_X1 port map( A1 => n16220, A2 => n15219, B1 => n16217, B2 => 
                           n14338, ZN => n13518);
   U6257 : AOI221_X1 port map( B1 => registers_7_11_port, B2 => n16226, C1 => 
                           registers_42_11_port, C2 => n16223, A => n13476, ZN 
                           => n13469);
   U6258 : OAI22_X1 port map( A1 => n16220, A2 => n15220, B1 => n16217, B2 => 
                           n14339, ZN => n13476);
   U6259 : AOI221_X1 port map( B1 => registers_7_12_port, B2 => n16227, C1 => 
                           registers_42_12_port, C2 => n16224, A => n13434, ZN 
                           => n13427);
   U6260 : OAI22_X1 port map( A1 => n16221, A2 => n15221, B1 => n16218, B2 => 
                           n14340, ZN => n13434);
   U6261 : AOI221_X1 port map( B1 => registers_7_13_port, B2 => n16227, C1 => 
                           registers_42_13_port, C2 => n16224, A => n13392, ZN 
                           => n13385);
   U6262 : OAI22_X1 port map( A1 => n16221, A2 => n15222, B1 => n16218, B2 => 
                           n14341, ZN => n13392);
   U6263 : AOI221_X1 port map( B1 => registers_7_14_port, B2 => n16227, C1 => 
                           registers_42_14_port, C2 => n16224, A => n13350, ZN 
                           => n13343);
   U6264 : OAI22_X1 port map( A1 => n16221, A2 => n15223, B1 => n16218, B2 => 
                           n14342, ZN => n13350);
   U6265 : AOI221_X1 port map( B1 => registers_7_15_port, B2 => n16227, C1 => 
                           registers_42_15_port, C2 => n16224, A => n13308, ZN 
                           => n13301);
   U6266 : OAI22_X1 port map( A1 => n16221, A2 => n15224, B1 => n16218, B2 => 
                           n14343, ZN => n13308);
   U6267 : AOI221_X1 port map( B1 => registers_7_16_port, B2 => n16227, C1 => 
                           registers_42_16_port, C2 => n16224, A => n13266, ZN 
                           => n13259);
   U6268 : OAI22_X1 port map( A1 => n16221, A2 => n15225, B1 => n16218, B2 => 
                           n14344, ZN => n13266);
   U6269 : AOI221_X1 port map( B1 => registers_7_17_port, B2 => n16227, C1 => 
                           registers_42_17_port, C2 => n16224, A => n13224, ZN 
                           => n13217);
   U6270 : OAI22_X1 port map( A1 => n16221, A2 => n15226, B1 => n16218, B2 => 
                           n14345, ZN => n13224);
   U6271 : AOI221_X1 port map( B1 => registers_7_18_port, B2 => n16227, C1 => 
                           registers_42_18_port, C2 => n16224, A => n13182, ZN 
                           => n13175);
   U6272 : OAI22_X1 port map( A1 => n16221, A2 => n15227, B1 => n16218, B2 => 
                           n14346, ZN => n13182);
   U6273 : AOI221_X1 port map( B1 => registers_7_19_port, B2 => n16227, C1 => 
                           registers_42_19_port, C2 => n16224, A => n13140, ZN 
                           => n13133);
   U6274 : OAI22_X1 port map( A1 => n16221, A2 => n15228, B1 => n16218, B2 => 
                           n14347, ZN => n13140);
   U6275 : AOI221_X1 port map( B1 => registers_7_20_port, B2 => n16227, C1 => 
                           registers_42_20_port, C2 => n16224, A => n13098, ZN 
                           => n13091);
   U6276 : OAI22_X1 port map( A1 => n16221, A2 => n15229, B1 => n16218, B2 => 
                           n14348, ZN => n13098);
   U6277 : AOI221_X1 port map( B1 => registers_7_21_port, B2 => n16227, C1 => 
                           registers_42_21_port, C2 => n16224, A => n13056, ZN 
                           => n13049);
   U6278 : OAI22_X1 port map( A1 => n16221, A2 => n15230, B1 => n16218, B2 => 
                           n14349, ZN => n13056);
   U6279 : AOI221_X1 port map( B1 => registers_7_22_port, B2 => n16227, C1 => 
                           registers_42_22_port, C2 => n16224, A => n13014, ZN 
                           => n13007);
   U6280 : OAI22_X1 port map( A1 => n16221, A2 => n15231, B1 => n16218, B2 => 
                           n14350, ZN => n13014);
   U6281 : AOI221_X1 port map( B1 => registers_7_23_port, B2 => n16227, C1 => 
                           registers_42_23_port, C2 => n16224, A => n12972, ZN 
                           => n12965);
   U6282 : OAI22_X1 port map( A1 => n16221, A2 => n15232, B1 => n16218, B2 => 
                           n14351, ZN => n12972);
   U6283 : AOI221_X1 port map( B1 => registers_50_0_port, B2 => n16529, C1 => 
                           net226846, C2 => n16526, A => n12478, ZN => n12467);
   U6284 : OAI22_X1 port map( A1 => n16523, A2 => n12356, B1 => n16520, B2 => 
                           n14938, ZN => n12478);
   U6285 : AOI221_X1 port map( B1 => registers_7_0_port, B2 => n16478, C1 => 
                           registers_42_0_port, C2 => n16475, A => n12496, ZN 
                           => n12483);
   U6286 : OAI22_X1 port map( A1 => n16472, A2 => n15210, B1 => n16469, B2 => 
                           n14329, ZN => n12496);
   U6287 : AOI221_X1 port map( B1 => registers_50_1_port, B2 => n16529, C1 => 
                           net226859, C2 => n16526, A => n12292, ZN => n12285);
   U6288 : OAI22_X1 port map( A1 => n16523, A2 => n12358, B1 => n16520, B2 => 
                           n14939, ZN => n12292);
   U6289 : AOI221_X1 port map( B1 => registers_7_1_port, B2 => n16478, C1 => 
                           registers_42_1_port, C2 => n16475, A => n12300, ZN 
                           => n12293);
   U6290 : OAI22_X1 port map( A1 => n16472, A2 => n15211, B1 => n16469, B2 => 
                           n14330, ZN => n12300);
   U6291 : AOI221_X1 port map( B1 => registers_50_2_port, B2 => n16529, C1 => 
                           net226885, C2 => n16526, A => n12139, ZN => n12132);
   U6292 : OAI22_X1 port map( A1 => n16523, A2 => n12360, B1 => n16520, B2 => 
                           n14940, ZN => n12139);
   U6293 : AOI221_X1 port map( B1 => registers_7_2_port, B2 => n16478, C1 => 
                           registers_42_2_port, C2 => n16475, A => n12147, ZN 
                           => n12140);
   U6294 : OAI22_X1 port map( A1 => n16472, A2 => n15212, B1 => n16469, B2 => 
                           n14331, ZN => n12147);
   U6295 : AOI221_X1 port map( B1 => registers_50_3_port, B2 => n16529, C1 => 
                           net226898, C2 => n16526, A => n11986, ZN => n11979);
   U6296 : OAI22_X1 port map( A1 => n16523, A2 => n12340, B1 => n16520, B2 => 
                           n14941, ZN => n11986);
   U6297 : AOI221_X1 port map( B1 => registers_7_3_port, B2 => n16478, C1 => 
                           registers_42_3_port, C2 => n16475, A => n11994, ZN 
                           => n11987);
   U6298 : OAI22_X1 port map( A1 => n16472, A2 => n15003, B1 => n16469, B2 => 
                           n14288, ZN => n11994);
   U6299 : AOI221_X1 port map( B1 => registers_50_4_port, B2 => n16529, C1 => 
                           net226980, C2 => n16526, A => n11833, ZN => n11826);
   U6300 : OAI22_X1 port map( A1 => n16523, A2 => n12341, B1 => n16520, B2 => 
                           n14866, ZN => n11833);
   U6301 : AOI221_X1 port map( B1 => registers_7_4_port, B2 => n16478, C1 => 
                           registers_42_4_port, C2 => n16475, A => n11841, ZN 
                           => n11834);
   U6302 : OAI22_X1 port map( A1 => n16472, A2 => n15213, B1 => n16469, B2 => 
                           n14332, ZN => n11841);
   U6303 : AOI221_X1 port map( B1 => registers_50_5_port, B2 => n16529, C1 => 
                           net227000, C2 => n16526, A => n11790, ZN => n11783);
   U6304 : OAI22_X1 port map( A1 => n16523, A2 => n12364, B1 => n16520, B2 => 
                           n14867, ZN => n11790);
   U6305 : AOI221_X1 port map( B1 => registers_7_5_port, B2 => n16478, C1 => 
                           registers_42_5_port, C2 => n16475, A => n11798, ZN 
                           => n11791);
   U6306 : OAI22_X1 port map( A1 => n16472, A2 => n15214, B1 => n16469, B2 => 
                           n14333, ZN => n11798);
   U6307 : AOI221_X1 port map( B1 => registers_50_6_port, B2 => n16529, C1 => 
                           net227011, C2 => n16526, A => n11747, ZN => n11740);
   U6308 : OAI22_X1 port map( A1 => n16523, A2 => n12366, B1 => n16520, B2 => 
                           n14942, ZN => n11747);
   U6309 : AOI221_X1 port map( B1 => registers_7_6_port, B2 => n16478, C1 => 
                           registers_42_6_port, C2 => n16475, A => n11755, ZN 
                           => n11748);
   U6310 : OAI22_X1 port map( A1 => n16472, A2 => n15215, B1 => n16469, B2 => 
                           n14334, ZN => n11755);
   U6311 : AOI221_X1 port map( B1 => registers_50_7_port, B2 => n16529, C1 => 
                           net227029, C2 => n16526, A => n11704, ZN => n11697);
   U6312 : OAI22_X1 port map( A1 => n16523, A2 => n12368, B1 => n16520, B2 => 
                           n14943, ZN => n11704);
   U6313 : AOI221_X1 port map( B1 => registers_7_7_port, B2 => n16478, C1 => 
                           registers_42_7_port, C2 => n16475, A => n11712, ZN 
                           => n11705);
   U6314 : OAI22_X1 port map( A1 => n16472, A2 => n15216, B1 => n16469, B2 => 
                           n14335, ZN => n11712);
   U6315 : AOI221_X1 port map( B1 => registers_50_8_port, B2 => n16529, C1 => 
                           net227047, C2 => n16526, A => n11661, ZN => n11654);
   U6316 : OAI22_X1 port map( A1 => n16523, A2 => n12407, B1 => n16520, B2 => 
                           n14944, ZN => n11661);
   U6317 : AOI221_X1 port map( B1 => registers_7_8_port, B2 => n16478, C1 => 
                           registers_42_8_port, C2 => n16475, A => n11669, ZN 
                           => n11662);
   U6318 : OAI22_X1 port map( A1 => n16472, A2 => n15217, B1 => n16469, B2 => 
                           n14336, ZN => n11669);
   U6319 : AOI221_X1 port map( B1 => registers_50_9_port, B2 => n16529, C1 => 
                           net227065, C2 => n16526, A => n11618, ZN => n11611);
   U6320 : OAI22_X1 port map( A1 => n16523, A2 => n12409, B1 => n16520, B2 => 
                           n14945, ZN => n11618);
   U6321 : AOI221_X1 port map( B1 => registers_7_9_port, B2 => n16478, C1 => 
                           registers_42_9_port, C2 => n16475, A => n11626, ZN 
                           => n11619);
   U6322 : OAI22_X1 port map( A1 => n16472, A2 => n15218, B1 => n16469, B2 => 
                           n14337, ZN => n11626);
   U6323 : AOI221_X1 port map( B1 => registers_50_10_port, B2 => n16529, C1 => 
                           net227083, C2 => n16526, A => n11575, ZN => n11568);
   U6324 : OAI22_X1 port map( A1 => n16523, A2 => n12411, B1 => n16520, B2 => 
                           n14946, ZN => n11575);
   U6325 : AOI221_X1 port map( B1 => registers_7_10_port, B2 => n16478, C1 => 
                           registers_42_10_port, C2 => n16475, A => n11583, ZN 
                           => n11576);
   U6326 : OAI22_X1 port map( A1 => n16472, A2 => n15219, B1 => n16469, B2 => 
                           n14338, ZN => n11583);
   U6327 : AOI221_X1 port map( B1 => registers_50_11_port, B2 => n16529, C1 => 
                           net227101, C2 => n16526, A => n11532, ZN => n11525);
   U6328 : OAI22_X1 port map( A1 => n16523, A2 => n12600, B1 => n16520, B2 => 
                           n14947, ZN => n11532);
   U6329 : AOI221_X1 port map( B1 => registers_7_11_port, B2 => n16478, C1 => 
                           registers_42_11_port, C2 => n16475, A => n11540, ZN 
                           => n11533);
   U6330 : OAI22_X1 port map( A1 => n16472, A2 => n15220, B1 => n16469, B2 => 
                           n14339, ZN => n11540);
   U6331 : AOI221_X1 port map( B1 => registers_50_12_port, B2 => n16530, C1 => 
                           net227119, C2 => n16527, A => n11489, ZN => n11482);
   U6332 : OAI22_X1 port map( A1 => n16524, A2 => n12652, B1 => n16521, B2 => 
                           n14948, ZN => n11489);
   U6333 : AOI221_X1 port map( B1 => registers_7_12_port, B2 => n16479, C1 => 
                           registers_42_12_port, C2 => n16476, A => n11497, ZN 
                           => n11490);
   U6334 : OAI22_X1 port map( A1 => n16473, A2 => n15221, B1 => n16470, B2 => 
                           n14340, ZN => n11497);
   U6335 : AOI221_X1 port map( B1 => registers_50_13_port, B2 => n16530, C1 => 
                           net227137, C2 => n16527, A => n11445, ZN => n11438);
   U6336 : OAI22_X1 port map( A1 => n16524, A2 => n13996, B1 => n16521, B2 => 
                           n14949, ZN => n11445);
   U6337 : AOI221_X1 port map( B1 => registers_7_13_port, B2 => n16479, C1 => 
                           registers_42_13_port, C2 => n16476, A => n11453, ZN 
                           => n11446);
   U6338 : OAI22_X1 port map( A1 => n16473, A2 => n15222, B1 => n16470, B2 => 
                           n14341, ZN => n11453);
   U6339 : AOI221_X1 port map( B1 => registers_50_14_port, B2 => n16530, C1 => 
                           net227155, C2 => n16527, A => n11402, ZN => n11395);
   U6340 : OAI22_X1 port map( A1 => n16524, A2 => n14008, B1 => n16521, B2 => 
                           n14950, ZN => n11402);
   U6341 : AOI221_X1 port map( B1 => registers_7_14_port, B2 => n16479, C1 => 
                           registers_42_14_port, C2 => n16476, A => n11410, ZN 
                           => n11403);
   U6342 : OAI22_X1 port map( A1 => n16473, A2 => n15223, B1 => n16470, B2 => 
                           n14342, ZN => n11410);
   U6343 : AOI221_X1 port map( B1 => registers_50_15_port, B2 => n16530, C1 => 
                           net227173, C2 => n16527, A => n11359, ZN => n11352);
   U6344 : OAI22_X1 port map( A1 => n16524, A2 => n14015, B1 => n16521, B2 => 
                           n14951, ZN => n11359);
   U6345 : AOI221_X1 port map( B1 => registers_7_15_port, B2 => n16479, C1 => 
                           registers_42_15_port, C2 => n16476, A => n11367, ZN 
                           => n11360);
   U6346 : OAI22_X1 port map( A1 => n16473, A2 => n15224, B1 => n16470, B2 => 
                           n14343, ZN => n11367);
   U6347 : AOI221_X1 port map( B1 => registers_50_16_port, B2 => n16530, C1 => 
                           net227191, C2 => n16527, A => n11316, ZN => n11309);
   U6348 : OAI22_X1 port map( A1 => n16524, A2 => n14035, B1 => n16521, B2 => 
                           n14952, ZN => n11316);
   U6349 : AOI221_X1 port map( B1 => registers_7_16_port, B2 => n16479, C1 => 
                           registers_42_16_port, C2 => n16476, A => n11324, ZN 
                           => n11317);
   U6350 : OAI22_X1 port map( A1 => n16473, A2 => n15225, B1 => n16470, B2 => 
                           n14344, ZN => n11324);
   U6351 : AOI221_X1 port map( B1 => registers_50_17_port, B2 => n16530, C1 => 
                           net227209, C2 => n16527, A => n11273, ZN => n11266);
   U6352 : OAI22_X1 port map( A1 => n16524, A2 => n14037, B1 => n16521, B2 => 
                           n14953, ZN => n11273);
   U6353 : AOI221_X1 port map( B1 => registers_7_17_port, B2 => n16479, C1 => 
                           registers_42_17_port, C2 => n16476, A => n11281, ZN 
                           => n11274);
   U6354 : OAI22_X1 port map( A1 => n16473, A2 => n15226, B1 => n16470, B2 => 
                           n14345, ZN => n11281);
   U6355 : AOI221_X1 port map( B1 => registers_50_18_port, B2 => n16530, C1 => 
                           net227227, C2 => n16527, A => n11230, ZN => n11223);
   U6356 : OAI22_X1 port map( A1 => n16524, A2 => n14039, B1 => n16521, B2 => 
                           n14954, ZN => n11230);
   U6357 : AOI221_X1 port map( B1 => registers_7_18_port, B2 => n16479, C1 => 
                           registers_42_18_port, C2 => n16476, A => n11238, ZN 
                           => n11231);
   U6358 : OAI22_X1 port map( A1 => n16473, A2 => n15227, B1 => n16470, B2 => 
                           n14346, ZN => n11238);
   U6359 : AOI221_X1 port map( B1 => registers_50_19_port, B2 => n16530, C1 => 
                           net227245, C2 => n16527, A => n11187, ZN => n11180);
   U6360 : OAI22_X1 port map( A1 => n16524, A2 => n14041, B1 => n16521, B2 => 
                           n14955, ZN => n11187);
   U6361 : AOI221_X1 port map( B1 => registers_7_19_port, B2 => n16479, C1 => 
                           registers_42_19_port, C2 => n16476, A => n11195, ZN 
                           => n11188);
   U6362 : OAI22_X1 port map( A1 => n16473, A2 => n15228, B1 => n16470, B2 => 
                           n14347, ZN => n11195);
   U6363 : AOI221_X1 port map( B1 => registers_50_20_port, B2 => n16530, C1 => 
                           net227263, C2 => n16527, A => n11144, ZN => n11137);
   U6364 : OAI22_X1 port map( A1 => n16524, A2 => n14043, B1 => n16521, B2 => 
                           n14956, ZN => n11144);
   U6365 : AOI221_X1 port map( B1 => registers_7_20_port, B2 => n16479, C1 => 
                           registers_42_20_port, C2 => n16476, A => n11152, ZN 
                           => n11145);
   U6366 : OAI22_X1 port map( A1 => n16473, A2 => n15229, B1 => n16470, B2 => 
                           n14348, ZN => n11152);
   U6367 : AOI221_X1 port map( B1 => registers_50_21_port, B2 => n16530, C1 => 
                           net227281, C2 => n16527, A => n11101, ZN => n11094);
   U6368 : OAI22_X1 port map( A1 => n16524, A2 => n14045, B1 => n16521, B2 => 
                           n14957, ZN => n11101);
   U6369 : AOI221_X1 port map( B1 => registers_7_21_port, B2 => n16479, C1 => 
                           registers_42_21_port, C2 => n16476, A => n11109, ZN 
                           => n11102);
   U6370 : OAI22_X1 port map( A1 => n16473, A2 => n15230, B1 => n16470, B2 => 
                           n14349, ZN => n11109);
   U6371 : AOI221_X1 port map( B1 => registers_50_22_port, B2 => n16530, C1 => 
                           net227299, C2 => n16527, A => n11058, ZN => n11051);
   U6372 : OAI22_X1 port map( A1 => n16524, A2 => n14047, B1 => n16521, B2 => 
                           n14958, ZN => n11058);
   U6373 : AOI221_X1 port map( B1 => registers_7_22_port, B2 => n16479, C1 => 
                           registers_42_22_port, C2 => n16476, A => n11066, ZN 
                           => n11059);
   U6374 : OAI22_X1 port map( A1 => n16473, A2 => n15231, B1 => n16470, B2 => 
                           n14350, ZN => n11066);
   U6375 : AOI221_X1 port map( B1 => registers_50_23_port, B2 => n16530, C1 => 
                           net227317, C2 => n16527, A => n11015, ZN => n11008);
   U6376 : OAI22_X1 port map( A1 => n16524, A2 => n14049, B1 => n16521, B2 => 
                           n14959, ZN => n11015);
   U6377 : AOI221_X1 port map( B1 => registers_7_23_port, B2 => n16479, C1 => 
                           registers_42_23_port, C2 => n16476, A => n11023, ZN 
                           => n11016);
   U6378 : OAI22_X1 port map( A1 => n16473, A2 => n15232, B1 => n16470, B2 => 
                           n14351, ZN => n11023);
   U6379 : AOI221_X1 port map( B1 => registers_48_0_port, B2 => n17637, C1 => 
                           registers_4_0_port, C2 => n17634, A => n12406, ZN =>
                           n12399);
   U6380 : OAI22_X1 port map( A1 => n17631, A2 => n15495, B1 => n17628, B2 => 
                           n14678, ZN => n12406);
   U6381 : AOI221_X1 port map( B1 => registers_23_0_port, B2 => n17781, C1 => 
                           registers_22_0_port, C2 => n17778, A => n12382, ZN 
                           => n12375);
   U6382 : OAI22_X1 port map( A1 => n17775, A2 => n12205, B1 => n17772, B2 => 
                           n14831, ZN => n12382);
   U6383 : AOI221_X1 port map( B1 => registers_48_1_port, B2 => n17637, C1 => 
                           registers_4_1_port, C2 => n17634, A => n12252, ZN =>
                           n12245);
   U6384 : OAI22_X1 port map( A1 => n17631, A2 => n15496, B1 => n17628, B2 => 
                           n14679, ZN => n12252);
   U6385 : AOI221_X1 port map( B1 => registers_23_1_port, B2 => n17781, C1 => 
                           registers_22_1_port, C2 => n17778, A => n12228, ZN 
                           => n12221);
   U6386 : OAI22_X1 port map( A1 => n17775, A2 => n12206, B1 => n17772, B2 => 
                           n14832, ZN => n12228);
   U6387 : AOI221_X1 port map( B1 => registers_48_2_port, B2 => n17637, C1 => 
                           registers_4_2_port, C2 => n17634, A => n12097, ZN =>
                           n12090);
   U6388 : OAI22_X1 port map( A1 => n17631, A2 => n15497, B1 => n17628, B2 => 
                           n14680, ZN => n12097);
   U6389 : AOI221_X1 port map( B1 => registers_23_2_port, B2 => n17781, C1 => 
                           registers_22_2_port, C2 => n17778, A => n12073, ZN 
                           => n12066);
   U6390 : OAI22_X1 port map( A1 => n17775, A2 => n12207, B1 => n17772, B2 => 
                           n14833, ZN => n12073);
   U6391 : AOI221_X1 port map( B1 => registers_48_3_port, B2 => n17637, C1 => 
                           registers_4_3_port, C2 => n17634, A => n11944, ZN =>
                           n11937);
   U6392 : OAI22_X1 port map( A1 => n17631, A2 => n15498, B1 => n17628, B2 => 
                           n14638, ZN => n11944);
   U6393 : AOI221_X1 port map( B1 => registers_23_3_port, B2 => n17781, C1 => 
                           registers_22_3_port, C2 => n17778, A => n11920, ZN 
                           => n11913);
   U6394 : OAI22_X1 port map( A1 => n17775, A2 => n12208, B1 => n17772, B2 => 
                           n14834, ZN => n11920);
   U6395 : AOI221_X1 port map( B1 => registers_48_4_port, B2 => n17637, C1 => 
                           registers_4_4_port, C2 => n17634, A => n10501, ZN =>
                           n10494);
   U6396 : OAI22_X1 port map( A1 => n17631, A2 => n15499, B1 => n17628, B2 => 
                           n14639, ZN => n10501);
   U6397 : AOI221_X1 port map( B1 => registers_23_4_port, B2 => n17781, C1 => 
                           registers_22_4_port, C2 => n17778, A => n10477, ZN 
                           => n10470);
   U6398 : OAI22_X1 port map( A1 => n17775, A2 => n12195, B1 => n17772, B2 => 
                           n14823, ZN => n10477);
   U6399 : AOI221_X1 port map( B1 => registers_48_5_port, B2 => n17637, C1 => 
                           registers_4_5_port, C2 => n17634, A => n10391, ZN =>
                           n10384);
   U6400 : OAI22_X1 port map( A1 => n17631, A2 => n15358, B1 => n17628, B2 => 
                           n14681, ZN => n10391);
   U6401 : AOI221_X1 port map( B1 => registers_23_5_port, B2 => n17781, C1 => 
                           registers_22_5_port, C2 => n17778, A => n10367, ZN 
                           => n10360);
   U6402 : OAI22_X1 port map( A1 => n17775, A2 => n12209, B1 => n17772, B2 => 
                           n14835, ZN => n10367);
   U6403 : AOI221_X1 port map( B1 => registers_48_6_port, B2 => n17637, C1 => 
                           registers_4_6_port, C2 => n17634, A => n10279, ZN =>
                           n10272);
   U6404 : OAI22_X1 port map( A1 => n17631, A2 => n15500, B1 => n17628, B2 => 
                           n14682, ZN => n10279);
   U6405 : AOI221_X1 port map( B1 => registers_23_6_port, B2 => n17781, C1 => 
                           registers_22_6_port, C2 => n17778, A => n10255, ZN 
                           => n10248);
   U6406 : OAI22_X1 port map( A1 => n17775, A2 => n12210, B1 => n17772, B2 => 
                           n14836, ZN => n10255);
   U6407 : AOI221_X1 port map( B1 => registers_48_7_port, B2 => n17637, C1 => 
                           registers_4_7_port, C2 => n17634, A => n7643, ZN => 
                           n7636);
   U6408 : OAI22_X1 port map( A1 => n17631, A2 => n15501, B1 => n17628, B2 => 
                           n14683, ZN => n7643);
   U6409 : AOI221_X1 port map( B1 => registers_23_7_port, B2 => n17781, C1 => 
                           registers_22_7_port, C2 => n17778, A => n7619, ZN =>
                           n7612);
   U6410 : OAI22_X1 port map( A1 => n17775, A2 => n12211, B1 => n17772, B2 => 
                           n14837, ZN => n7619);
   U6411 : AOI221_X1 port map( B1 => registers_48_8_port, B2 => n17637, C1 => 
                           registers_4_8_port, C2 => n17634, A => n7528, ZN => 
                           n7521);
   U6412 : OAI22_X1 port map( A1 => n17631, A2 => n15502, B1 => n17628, B2 => 
                           n14684, ZN => n7528);
   U6413 : AOI221_X1 port map( B1 => registers_23_8_port, B2 => n17781, C1 => 
                           registers_22_8_port, C2 => n17778, A => n7504, ZN =>
                           n7497);
   U6414 : OAI22_X1 port map( A1 => n17775, A2 => n12212, B1 => n17772, B2 => 
                           n14838, ZN => n7504);
   U6415 : AOI221_X1 port map( B1 => registers_48_9_port, B2 => n17637, C1 => 
                           registers_4_9_port, C2 => n17634, A => n7419, ZN => 
                           n7412);
   U6416 : OAI22_X1 port map( A1 => n17631, A2 => n15503, B1 => n17628, B2 => 
                           n14685, ZN => n7419);
   U6417 : AOI221_X1 port map( B1 => registers_23_9_port, B2 => n17781, C1 => 
                           registers_22_9_port, C2 => n17778, A => n7395, ZN =>
                           n7388);
   U6418 : OAI22_X1 port map( A1 => n17775, A2 => n12213, B1 => n17772, B2 => 
                           n14839, ZN => n7395);
   U6419 : AOI221_X1 port map( B1 => registers_48_10_port, B2 => n17637, C1 => 
                           registers_4_10_port, C2 => n17634, A => n7310, ZN =>
                           n7303);
   U6420 : OAI22_X1 port map( A1 => n17631, A2 => n15504, B1 => n17628, B2 => 
                           n14686, ZN => n7310);
   U6421 : AOI221_X1 port map( B1 => registers_23_10_port, B2 => n17781, C1 => 
                           registers_22_10_port, C2 => n17778, A => n7286, ZN 
                           => n7279);
   U6422 : OAI22_X1 port map( A1 => n17775, A2 => n12214, B1 => n17772, B2 => 
                           n14840, ZN => n7286);
   U6423 : AOI221_X1 port map( B1 => registers_48_11_port, B2 => n17638, C1 => 
                           registers_4_11_port, C2 => n17635, A => n7196, ZN =>
                           n7189);
   U6424 : OAI22_X1 port map( A1 => n17632, A2 => n15505, B1 => n17629, B2 => 
                           n14687, ZN => n7196);
   U6425 : AOI221_X1 port map( B1 => registers_23_11_port, B2 => n17782, C1 => 
                           registers_22_11_port, C2 => n17779, A => n7172, ZN 
                           => n7165);
   U6426 : OAI22_X1 port map( A1 => n17776, A2 => n12215, B1 => n17773, B2 => 
                           n14841, ZN => n7172);
   U6427 : AOI221_X1 port map( B1 => registers_48_12_port, B2 => n17638, C1 => 
                           registers_4_12_port, C2 => n17635, A => n7087, ZN =>
                           n7080);
   U6428 : OAI22_X1 port map( A1 => n17632, A2 => n15506, B1 => n17629, B2 => 
                           n14688, ZN => n7087);
   U6429 : AOI221_X1 port map( B1 => registers_23_12_port, B2 => n17782, C1 => 
                           registers_22_12_port, C2 => n17779, A => n7063, ZN 
                           => n7056);
   U6430 : OAI22_X1 port map( A1 => n17776, A2 => n12253, B1 => n17773, B2 => 
                           n14842, ZN => n7063);
   U6431 : AOI221_X1 port map( B1 => registers_48_13_port, B2 => n17638, C1 => 
                           registers_4_13_port, C2 => n17635, A => n6978, ZN =>
                           n6971);
   U6432 : OAI22_X1 port map( A1 => n17632, A2 => n15507, B1 => n17629, B2 => 
                           n14689, ZN => n6978);
   U6433 : AOI221_X1 port map( B1 => registers_23_13_port, B2 => n17782, C1 => 
                           registers_22_13_port, C2 => n17779, A => n6954, ZN 
                           => n6947);
   U6434 : OAI22_X1 port map( A1 => n17776, A2 => n12254, B1 => n17773, B2 => 
                           n14843, ZN => n6954);
   U6435 : AOI221_X1 port map( B1 => registers_48_14_port, B2 => n17638, C1 => 
                           registers_4_14_port, C2 => n17635, A => n6869, ZN =>
                           n6862);
   U6436 : OAI22_X1 port map( A1 => n17632, A2 => n15508, B1 => n17629, B2 => 
                           n14690, ZN => n6869);
   U6437 : AOI221_X1 port map( B1 => registers_23_14_port, B2 => n17782, C1 => 
                           registers_22_14_port, C2 => n17779, A => n6845, ZN 
                           => n6838);
   U6438 : OAI22_X1 port map( A1 => n17776, A2 => n12255, B1 => n17773, B2 => 
                           n14844, ZN => n6845);
   U6439 : AOI221_X1 port map( B1 => registers_48_15_port, B2 => n17638, C1 => 
                           registers_4_15_port, C2 => n17635, A => n6760, ZN =>
                           n6753);
   U6440 : OAI22_X1 port map( A1 => n17632, A2 => n15509, B1 => n17629, B2 => 
                           n14691, ZN => n6760);
   U6441 : AOI221_X1 port map( B1 => registers_23_15_port, B2 => n17782, C1 => 
                           registers_22_15_port, C2 => n17779, A => n6736, ZN 
                           => n6729);
   U6442 : OAI22_X1 port map( A1 => n17776, A2 => n12256, B1 => n17773, B2 => 
                           n14845, ZN => n6736);
   U6443 : AOI221_X1 port map( B1 => registers_48_16_port, B2 => n17638, C1 => 
                           registers_4_16_port, C2 => n17635, A => n6622, ZN =>
                           n6612);
   U6444 : OAI22_X1 port map( A1 => n17632, A2 => n15510, B1 => n17629, B2 => 
                           n14692, ZN => n6622);
   U6445 : AOI221_X1 port map( B1 => registers_23_16_port, B2 => n17782, C1 => 
                           registers_22_16_port, C2 => n17779, A => n6576, ZN 
                           => n6566);
   U6446 : OAI22_X1 port map( A1 => n17776, A2 => n12257, B1 => n17773, B2 => 
                           n14846, ZN => n6576);
   U6447 : AOI221_X1 port map( B1 => registers_48_17_port, B2 => n17638, C1 => 
                           registers_4_17_port, C2 => n17635, A => n6436, ZN =>
                           n6426);
   U6448 : OAI22_X1 port map( A1 => n17632, A2 => n15511, B1 => n17629, B2 => 
                           n14693, ZN => n6436);
   U6449 : AOI221_X1 port map( B1 => registers_23_17_port, B2 => n17782, C1 => 
                           registers_22_17_port, C2 => n17779, A => n6391, ZN 
                           => n6381);
   U6450 : OAI22_X1 port map( A1 => n17776, A2 => n12258, B1 => n17773, B2 => 
                           n14847, ZN => n6391);
   U6451 : AOI221_X1 port map( B1 => registers_48_18_port, B2 => n17638, C1 => 
                           registers_4_18_port, C2 => n17635, A => n6249, ZN =>
                           n6239);
   U6452 : OAI22_X1 port map( A1 => n17632, A2 => n15512, B1 => n17629, B2 => 
                           n14694, ZN => n6249);
   U6453 : AOI221_X1 port map( B1 => registers_23_18_port, B2 => n17782, C1 => 
                           registers_22_18_port, C2 => n17779, A => n6204, ZN 
                           => n6195);
   U6454 : OAI22_X1 port map( A1 => n17776, A2 => n12301, B1 => n17773, B2 => 
                           n14848, ZN => n6204);
   U6455 : AOI221_X1 port map( B1 => registers_48_19_port, B2 => n17638, C1 => 
                           registers_4_19_port, C2 => n17635, A => n6062, ZN =>
                           n6052);
   U6456 : OAI22_X1 port map( A1 => n17632, A2 => n15513, B1 => n17629, B2 => 
                           n14695, ZN => n6062);
   U6457 : AOI221_X1 port map( B1 => registers_23_19_port, B2 => n17782, C1 => 
                           registers_22_19_port, C2 => n17779, A => n6032, ZN 
                           => n6008);
   U6458 : OAI22_X1 port map( A1 => n17776, A2 => n12303, B1 => n17773, B2 => 
                           n14849, ZN => n6032);
   U6459 : AOI221_X1 port map( B1 => registers_48_20_port, B2 => n17638, C1 => 
                           registers_4_20_port, C2 => n17635, A => n5877, ZN =>
                           n5867);
   U6460 : OAI22_X1 port map( A1 => n17632, A2 => n15514, B1 => n17629, B2 => 
                           n14696, ZN => n5877);
   U6461 : AOI221_X1 port map( B1 => registers_23_20_port, B2 => n17782, C1 => 
                           registers_22_20_port, C2 => n17779, A => n5845, ZN 
                           => n5821);
   U6462 : OAI22_X1 port map( A1 => n17776, A2 => n12304, B1 => n17773, B2 => 
                           n14850, ZN => n5845);
   U6463 : AOI221_X1 port map( B1 => registers_48_21_port, B2 => n17638, C1 => 
                           registers_4_21_port, C2 => n17635, A => n5691, ZN =>
                           n5681);
   U6464 : OAI22_X1 port map( A1 => n17632, A2 => n15515, B1 => n17629, B2 => 
                           n14697, ZN => n5691);
   U6465 : AOI221_X1 port map( B1 => registers_23_21_port, B2 => n17782, C1 => 
                           registers_22_21_port, C2 => n17779, A => n5658, ZN 
                           => n5636);
   U6466 : OAI22_X1 port map( A1 => n17776, A2 => n12305, B1 => n17773, B2 => 
                           n14851, ZN => n5658);
   U6467 : AOI221_X1 port map( B1 => registers_48_22_port, B2 => n17638, C1 => 
                           registers_4_22_port, C2 => n17635, A => n5504, ZN =>
                           n5494);
   U6468 : OAI22_X1 port map( A1 => n17632, A2 => n15516, B1 => n17629, B2 => 
                           n14698, ZN => n5504);
   U6469 : AOI221_X1 port map( B1 => registers_23_22_port, B2 => n17782, C1 => 
                           registers_22_22_port, C2 => n17779, A => n5471, ZN 
                           => n5464);
   U6470 : OAI22_X1 port map( A1 => n17776, A2 => n12306, B1 => n17773, B2 => 
                           n14852, ZN => n5471);
   U6471 : AOI221_X1 port map( B1 => registers_48_31_port, B2 => n17637, C1 => 
                           registers_4_31_port, C2 => n17634, A => n14210, ZN 
                           => n14187);
   U6472 : OAI22_X1 port map( A1 => n17631, A2 => n15517, B1 => n17628, B2 => 
                           n14699, ZN => n14210);
   U6473 : AOI221_X1 port map( B1 => registers_23_31_port, B2 => n17781, C1 => 
                           registers_22_31_port, C2 => n17778, A => n14106, ZN 
                           => n14080);
   U6474 : OAI22_X1 port map( A1 => n17775, A2 => n12307, B1 => n17772, B2 => 
                           n14853, ZN => n14106);
   U6475 : NOR2_X1 port map( A1 => n14097, A2 => call, ZN => n14092);
   U6476 : NOR2_X1 port map( A1 => n14003, A2 => r590_carry_5_port, ZN => 
                           n14196);
   U6477 : NOR2_X1 port map( A1 => N9909, A2 => n10190, ZN => n14129);
   U6478 : AOI21_X1 port map( B1 => n14103, B2 => n14095, A => n14192, ZN => 
                           n4223);
   U6479 : AND3_X1 port map( A1 => n14193, A2 => call, A3 => n14194, ZN => 
                           n14192);
   U6480 : AOI22_X1 port map( A1 => net226843, A2 => n16466, B1 => 
                           registers_68_0_port, B2 => n16463, ZN => n12416);
   U6481 : AOI221_X1 port map( B1 => net226842, B2 => n16687, C1 => net226833, 
                           C2 => n16682, A => n12419, ZN => n12418);
   U6482 : AOI221_X1 port map( B1 => net226835, B2 => n16675, C1 => net226834, 
                           C2 => n16670, A => n12425, ZN => n12417);
   U6483 : AOI22_X1 port map( A1 => net227456, A2 => n16466, B1 => 
                           registers_68_31_port, B2 => n16463, ZN => n10513);
   U6484 : AOI221_X1 port map( B1 => net227454, B2 => n16687, C1 => net227453, 
                           C2 => n16682, A => n10518, ZN => n10515);
   U6485 : AOI221_X1 port map( B1 => net227457, B2 => n16675, C1 => net227455, 
                           C2 => n16670, A => n10524, ZN => n10514);
   U6486 : AOI22_X1 port map( A1 => n16216, A2 => net227330, B1 => n16211, B2 
                           => registers_68_24_port, ZN => n12889);
   U6487 : AOI221_X1 port map( B1 => n16435, B2 => net227328, C1 => n16432, C2 
                           => net227327, A => n12892, ZN => n12891);
   U6488 : AOI221_X1 port map( B1 => n16423, B2 => net227331, C1 => n16420, C2 
                           => net227329, A => n12893, ZN => n12890);
   U6489 : AOI22_X1 port map( A1 => n16216, A2 => net227348, B1 => n16211, B2 
                           => registers_68_25_port, ZN => n12847);
   U6490 : AOI221_X1 port map( B1 => n16435, B2 => net227346, C1 => n16432, C2 
                           => net227345, A => n12850, ZN => n12849);
   U6491 : AOI221_X1 port map( B1 => n16423, B2 => net227349, C1 => n16420, C2 
                           => net227347, A => n12851, ZN => n12848);
   U6492 : AOI22_X1 port map( A1 => n16216, A2 => net227366, B1 => n16211, B2 
                           => registers_68_26_port, ZN => n12805);
   U6493 : AOI221_X1 port map( B1 => n16435, B2 => net227364, C1 => n16432, C2 
                           => net227363, A => n12808, ZN => n12807);
   U6494 : AOI221_X1 port map( B1 => n16423, B2 => net227367, C1 => n16420, C2 
                           => net227365, A => n12809, ZN => n12806);
   U6495 : AOI22_X1 port map( A1 => n16216, A2 => net227384, B1 => n16211, B2 
                           => registers_68_27_port, ZN => n12763);
   U6496 : AOI221_X1 port map( B1 => n16435, B2 => net227382, C1 => n16432, C2 
                           => net227381, A => n12766, ZN => n12765);
   U6497 : AOI221_X1 port map( B1 => n16423, B2 => net227385, C1 => n16420, C2 
                           => net227383, A => n12767, ZN => n12764);
   U6498 : AOI22_X1 port map( A1 => n16216, A2 => net227402, B1 => n16211, B2 
                           => registers_68_28_port, ZN => n12721);
   U6499 : AOI221_X1 port map( B1 => n16435, B2 => net227400, C1 => n16432, C2 
                           => net227399, A => n12724, ZN => n12723);
   U6500 : AOI221_X1 port map( B1 => n16423, B2 => net227403, C1 => n16420, C2 
                           => net227401, A => n12725, ZN => n12722);
   U6501 : AOI22_X1 port map( A1 => n16216, A2 => net227420, B1 => n16211, B2 
                           => registers_68_29_port, ZN => n12679);
   U6502 : AOI221_X1 port map( B1 => n16435, B2 => net227418, C1 => n16432, C2 
                           => net227417, A => n12682, ZN => n12681);
   U6503 : AOI221_X1 port map( B1 => n16423, B2 => net227421, C1 => n16420, C2 
                           => net227419, A => n12683, ZN => n12680);
   U6504 : AOI22_X1 port map( A1 => n16216, A2 => net227438, B1 => n16211, B2 
                           => registers_68_30_port, ZN => n12635);
   U6505 : AOI221_X1 port map( B1 => n16435, B2 => net227436, C1 => n16432, C2 
                           => net227435, A => n12638, ZN => n12637);
   U6506 : AOI221_X1 port map( B1 => n16423, B2 => net227439, C1 => n16420, C2 
                           => net227437, A => n12639, ZN => n12636);
   U6507 : AOI22_X1 port map( A1 => n16216, A2 => net227456, B1 => n16211, B2 
                           => registers_68_31_port, ZN => n12516);
   U6508 : AOI221_X1 port map( B1 => n16435, B2 => net227454, C1 => n16432, C2 
                           => net227453, A => n12521, ZN => n12518);
   U6509 : AOI221_X1 port map( B1 => n16423, B2 => net227457, C1 => n16420, C2 
                           => net227455, A => n12526, ZN => n12517);
   U6510 : AOI22_X1 port map( A1 => n16468, A2 => net226988, B1 => n16465, B2 
                           => registers_68_5_port, ZN => n11757);
   U6511 : AOI221_X1 port map( B1 => n16687, B2 => net226986, C1 => n16684, C2 
                           => net226985, A => n11760, ZN => n11759);
   U6512 : AOI221_X1 port map( B1 => n16675, B2 => net226989, C1 => n16672, C2 
                           => net226987, A => n11761, ZN => n11758);
   U6513 : AOI22_X1 port map( A1 => n16468, A2 => net227006, B1 => n16465, B2 
                           => registers_68_6_port, ZN => n11714);
   U6514 : AOI221_X1 port map( B1 => n16687, B2 => net227004, C1 => n16684, C2 
                           => net227003, A => n11717, ZN => n11716);
   U6515 : AOI221_X1 port map( B1 => n16675, B2 => net227007, C1 => n16672, C2 
                           => net227005, A => n11718, ZN => n11715);
   U6516 : NOR2_X1 port map( A1 => n14201, A2 => call, ZN => n14152);
   U6517 : AOI21_X1 port map( B1 => n14151, B2 => n14092, A => n14169, ZN => 
                           n4202);
   U6518 : AND3_X1 port map( A1 => n14140, A2 => call, A3 => n14170, ZN => 
                           n14169);
   U6519 : NOR2_X1 port map( A1 => n10189, A2 => n10187, ZN => n14128);
   U6520 : NOR2_X1 port map( A1 => N9908, A2 => n10187, ZN => n14146);
   U6521 : OAI21_X1 port map( B1 => n14090, B2 => n14201, A => n14211, ZN => 
                           n4240);
   U6522 : NOR2_X1 port map( A1 => n14089, A2 => call, ZN => n14149);
   U6523 : NOR2_X1 port map( A1 => n14098, A2 => call, ZN => n14150);
   U6524 : AOI221_X1 port map( B1 => registers_56_23_port, B2 => n17675, C1 => 
                           registers_55_23_port, C2 => n17672, A => n5314, ZN 
                           => n5313);
   U6525 : OAI22_X1 port map( A1 => n17669, A2 => n15518, B1 => n17666, B2 => 
                           n14817, ZN => n5314);
   U6526 : AOI221_X1 port map( B1 => registers_56_24_port, B2 => n17675, C1 => 
                           registers_55_24_port, C2 => n17672, A => n5142, ZN 
                           => n5141);
   U6527 : OAI22_X1 port map( A1 => n17669, A2 => n15519, B1 => n17666, B2 => 
                           n14818, ZN => n5142);
   U6528 : AOI221_X1 port map( B1 => registers_56_25_port, B2 => n17675, C1 => 
                           registers_55_25_port, C2 => n17672, A => n5028, ZN 
                           => n5027);
   U6529 : OAI22_X1 port map( A1 => n17669, A2 => n15520, B1 => n17666, B2 => 
                           n14819, ZN => n5028);
   U6530 : AOI221_X1 port map( B1 => registers_56_30_port, B2 => n17675, C1 => 
                           registers_55_30_port, C2 => n17672, A => n4221, ZN 
                           => n4218);
   U6531 : OAI22_X1 port map( A1 => n17669, A2 => n15315, B1 => n17666, B2 => 
                           n14632, ZN => n4221);
   U6532 : AOI221_X1 port map( B1 => net227344, B2 => n16315, C1 => 
                           registers_44_24_port, C2 => n16312, A => n12919, ZN 
                           => n12918);
   U6533 : OAI22_X1 port map( A1 => n16309, A2 => n15144, B1 => n16306, B2 => 
                           n14527, ZN => n12919);
   U6534 : AOI221_X1 port map( B1 => registers_7_24_port, B2 => n16228, C1 => 
                           registers_42_24_port, C2 => n16225, A => n12930, ZN 
                           => n12923);
   U6535 : OAI22_X1 port map( A1 => n16222, A2 => n15233, B1 => n16219, B2 => 
                           n14352, ZN => n12930);
   U6536 : AOI221_X1 port map( B1 => net227362, B2 => n16315, C1 => 
                           registers_44_25_port, C2 => n16312, A => n12877, ZN 
                           => n12876);
   U6537 : OAI22_X1 port map( A1 => n16309, A2 => n15145, B1 => n16306, B2 => 
                           n14528, ZN => n12877);
   U6538 : AOI221_X1 port map( B1 => registers_7_25_port, B2 => n16228, C1 => 
                           registers_42_25_port, C2 => n16225, A => n12888, ZN 
                           => n12881);
   U6539 : OAI22_X1 port map( A1 => n16222, A2 => n15234, B1 => n16219, B2 => 
                           n14353, ZN => n12888);
   U6540 : AOI221_X1 port map( B1 => net227380, B2 => n16315, C1 => 
                           registers_44_26_port, C2 => n16312, A => n12835, ZN 
                           => n12834);
   U6541 : OAI22_X1 port map( A1 => n16309, A2 => n15146, B1 => n16306, B2 => 
                           n14529, ZN => n12835);
   U6542 : AOI221_X1 port map( B1 => registers_7_26_port, B2 => n16228, C1 => 
                           registers_42_26_port, C2 => n16225, A => n12846, ZN 
                           => n12839);
   U6543 : OAI22_X1 port map( A1 => n16222, A2 => n15235, B1 => n16219, B2 => 
                           n14354, ZN => n12846);
   U6544 : AOI221_X1 port map( B1 => net227398, B2 => n16315, C1 => 
                           registers_44_27_port, C2 => n16312, A => n12793, ZN 
                           => n12792);
   U6545 : OAI22_X1 port map( A1 => n16309, A2 => n15147, B1 => n16306, B2 => 
                           n14530, ZN => n12793);
   U6546 : AOI221_X1 port map( B1 => registers_7_27_port, B2 => n16228, C1 => 
                           registers_42_27_port, C2 => n16225, A => n12804, ZN 
                           => n12797);
   U6547 : OAI22_X1 port map( A1 => n16222, A2 => n15236, B1 => n16219, B2 => 
                           n14355, ZN => n12804);
   U6548 : AOI221_X1 port map( B1 => net227416, B2 => n16315, C1 => 
                           registers_44_28_port, C2 => n16312, A => n12751, ZN 
                           => n12750);
   U6549 : OAI22_X1 port map( A1 => n16309, A2 => n15148, B1 => n16306, B2 => 
                           n14531, ZN => n12751);
   U6550 : AOI221_X1 port map( B1 => registers_7_28_port, B2 => n16228, C1 => 
                           registers_42_28_port, C2 => n16225, A => n12762, ZN 
                           => n12755);
   U6551 : OAI22_X1 port map( A1 => n16222, A2 => n15237, B1 => n16219, B2 => 
                           n14356, ZN => n12762);
   U6552 : AOI221_X1 port map( B1 => net227434, B2 => n16315, C1 => 
                           registers_44_29_port, C2 => n16312, A => n12709, ZN 
                           => n12708);
   U6553 : OAI22_X1 port map( A1 => n16309, A2 => n15149, B1 => n16306, B2 => 
                           n14532, ZN => n12709);
   U6554 : AOI221_X1 port map( B1 => registers_7_29_port, B2 => n16228, C1 => 
                           registers_42_29_port, C2 => n16225, A => n12720, ZN 
                           => n12713);
   U6555 : OAI22_X1 port map( A1 => n16222, A2 => n15238, B1 => n16219, B2 => 
                           n14357, ZN => n12720);
   U6556 : AOI221_X1 port map( B1 => net227452, B2 => n16315, C1 => 
                           registers_44_30_port, C2 => n16312, A => n12666, ZN 
                           => n12665);
   U6557 : OAI22_X1 port map( A1 => n16309, A2 => n14871, B1 => n16306, B2 => 
                           n14069, ZN => n12666);
   U6558 : AOI221_X1 port map( B1 => registers_7_30_port, B2 => n16228, C1 => 
                           registers_42_30_port, C2 => n16225, A => n12678, ZN 
                           => n12671);
   U6559 : OAI22_X1 port map( A1 => n16222, A2 => n14874, B1 => n16219, B2 => 
                           n14055, ZN => n12678);
   U6560 : AOI221_X1 port map( B1 => net227470, B2 => n16315, C1 => 
                           registers_44_31_port, C2 => n16312, A => n12588, ZN 
                           => n12585);
   U6561 : OAI22_X1 port map( A1 => n16309, A2 => n15150, B1 => n16306, B2 => 
                           n14533, ZN => n12588);
   U6562 : AOI221_X1 port map( B1 => registers_7_31_port, B2 => n16228, C1 => 
                           registers_42_31_port, C2 => n16225, A => n12630, ZN 
                           => n12608);
   U6563 : OAI22_X1 port map( A1 => n16222, A2 => n15239, B1 => n16219, B2 => 
                           n14358, ZN => n12630);
   U6564 : AOI221_X1 port map( B1 => registers_50_0_port, B2 => n16277, C1 => 
                           net226846, C2 => n16274, A => n13959, ZN => n13948);
   U6565 : OAI22_X1 port map( A1 => n16271, A2 => n12356, B1 => n16268, B2 => 
                           n14938, ZN => n13959);
   U6566 : AOI221_X1 port map( B1 => registers_5_0_port, B2 => n16250, C1 => 
                           registers_59_0_port, C2 => n16247, A => n13971, ZN 
                           => n13966);
   U6567 : OAI22_X1 port map( A1 => n16244, A2 => n12357, B1 => n16241, B2 => 
                           n14910, ZN => n13971);
   U6568 : AOI221_X1 port map( B1 => registers_50_1_port, B2 => n16277, C1 => 
                           net226859, C2 => n16274, A => n13888, ZN => n13881);
   U6569 : OAI22_X1 port map( A1 => n16271, A2 => n12358, B1 => n16268, B2 => 
                           n14939, ZN => n13888);
   U6570 : AOI221_X1 port map( B1 => registers_5_1_port, B2 => n16250, C1 => 
                           registers_59_1_port, C2 => n16247, A => n13894, ZN 
                           => n13891);
   U6571 : OAI22_X1 port map( A1 => n16244, A2 => n12359, B1 => n16241, B2 => 
                           n14911, ZN => n13894);
   U6572 : AOI221_X1 port map( B1 => registers_50_2_port, B2 => n16277, C1 => 
                           net226885, C2 => n16274, A => n13846, ZN => n13839);
   U6573 : OAI22_X1 port map( A1 => n16271, A2 => n12360, B1 => n16268, B2 => 
                           n14940, ZN => n13846);
   U6574 : AOI221_X1 port map( B1 => registers_5_2_port, B2 => n16250, C1 => 
                           registers_59_2_port, C2 => n16247, A => n13852, ZN 
                           => n13849);
   U6575 : OAI22_X1 port map( A1 => n16244, A2 => n12361, B1 => n16241, B2 => 
                           n14912, ZN => n13852);
   U6576 : AOI221_X1 port map( B1 => registers_50_3_port, B2 => n16277, C1 => 
                           net226898, C2 => n16274, A => n13804, ZN => n13797);
   U6577 : OAI22_X1 port map( A1 => n16271, A2 => n12340, B1 => n16268, B2 => 
                           n14941, ZN => n13804);
   U6578 : AOI221_X1 port map( B1 => registers_5_3_port, B2 => n16250, C1 => 
                           registers_59_3_port, C2 => n16247, A => n13810, ZN 
                           => n13807);
   U6579 : OAI22_X1 port map( A1 => n16244, A2 => n12362, B1 => n16241, B2 => 
                           n14863, ZN => n13810);
   U6580 : AOI221_X1 port map( B1 => registers_50_4_port, B2 => n16277, C1 => 
                           net226980, C2 => n16274, A => n13762, ZN => n13755);
   U6581 : OAI22_X1 port map( A1 => n16271, A2 => n12341, B1 => n16268, B2 => 
                           n14866, ZN => n13762);
   U6582 : AOI221_X1 port map( B1 => registers_5_4_port, B2 => n16250, C1 => 
                           registers_59_4_port, C2 => n16247, A => n13768, ZN 
                           => n13765);
   U6583 : OAI22_X1 port map( A1 => n16244, A2 => n12363, B1 => n16241, B2 => 
                           n14864, ZN => n13768);
   U6584 : AOI221_X1 port map( B1 => registers_50_5_port, B2 => n16277, C1 => 
                           net227000, C2 => n16274, A => n13720, ZN => n13713);
   U6585 : OAI22_X1 port map( A1 => n16271, A2 => n12364, B1 => n16268, B2 => 
                           n14867, ZN => n13720);
   U6586 : AOI221_X1 port map( B1 => registers_5_5_port, B2 => n16250, C1 => 
                           registers_59_5_port, C2 => n16247, A => n13726, ZN 
                           => n13723);
   U6587 : OAI22_X1 port map( A1 => n16244, A2 => n12365, B1 => n16241, B2 => 
                           n14865, ZN => n13726);
   U6588 : AOI221_X1 port map( B1 => registers_50_6_port, B2 => n16277, C1 => 
                           net227011, C2 => n16274, A => n13678, ZN => n13671);
   U6589 : OAI22_X1 port map( A1 => n16271, A2 => n12366, B1 => n16268, B2 => 
                           n14942, ZN => n13678);
   U6590 : AOI221_X1 port map( B1 => registers_5_6_port, B2 => n16250, C1 => 
                           registers_59_6_port, C2 => n16247, A => n13684, ZN 
                           => n13681);
   U6591 : OAI22_X1 port map( A1 => n16244, A2 => n12367, B1 => n16241, B2 => 
                           n14913, ZN => n13684);
   U6592 : AOI221_X1 port map( B1 => registers_50_7_port, B2 => n16277, C1 => 
                           net227029, C2 => n16274, A => n13636, ZN => n13629);
   U6593 : OAI22_X1 port map( A1 => n16271, A2 => n12368, B1 => n16268, B2 => 
                           n14943, ZN => n13636);
   U6594 : AOI221_X1 port map( B1 => registers_5_7_port, B2 => n16250, C1 => 
                           registers_59_7_port, C2 => n16247, A => n13642, ZN 
                           => n13639);
   U6595 : OAI22_X1 port map( A1 => n16244, A2 => n12369, B1 => n16241, B2 => 
                           n14914, ZN => n13642);
   U6596 : AOI221_X1 port map( B1 => registers_50_8_port, B2 => n16277, C1 => 
                           net227047, C2 => n16274, A => n13594, ZN => n13587);
   U6597 : OAI22_X1 port map( A1 => n16271, A2 => n12407, B1 => n16268, B2 => 
                           n14944, ZN => n13594);
   U6598 : AOI221_X1 port map( B1 => registers_5_8_port, B2 => n16250, C1 => 
                           registers_59_8_port, C2 => n16247, A => n13600, ZN 
                           => n13597);
   U6599 : OAI22_X1 port map( A1 => n16244, A2 => n12408, B1 => n16241, B2 => 
                           n14915, ZN => n13600);
   U6600 : AOI221_X1 port map( B1 => registers_50_9_port, B2 => n16277, C1 => 
                           net227065, C2 => n16274, A => n13552, ZN => n13545);
   U6601 : OAI22_X1 port map( A1 => n16271, A2 => n12409, B1 => n16268, B2 => 
                           n14945, ZN => n13552);
   U6602 : AOI221_X1 port map( B1 => registers_5_9_port, B2 => n16250, C1 => 
                           registers_59_9_port, C2 => n16247, A => n13558, ZN 
                           => n13555);
   U6603 : OAI22_X1 port map( A1 => n16244, A2 => n12410, B1 => n16241, B2 => 
                           n14916, ZN => n13558);
   U6604 : AOI221_X1 port map( B1 => registers_50_10_port, B2 => n16277, C1 => 
                           net227083, C2 => n16274, A => n13510, ZN => n13503);
   U6605 : OAI22_X1 port map( A1 => n16271, A2 => n12411, B1 => n16268, B2 => 
                           n14946, ZN => n13510);
   U6606 : AOI221_X1 port map( B1 => registers_5_10_port, B2 => n16250, C1 => 
                           registers_59_10_port, C2 => n16247, A => n13516, ZN 
                           => n13513);
   U6607 : OAI22_X1 port map( A1 => n16244, A2 => n12551, B1 => n16241, B2 => 
                           n14917, ZN => n13516);
   U6608 : AOI221_X1 port map( B1 => registers_50_11_port, B2 => n16277, C1 => 
                           net227101, C2 => n16274, A => n13468, ZN => n13461);
   U6609 : OAI22_X1 port map( A1 => n16271, A2 => n12600, B1 => n16268, B2 => 
                           n14947, ZN => n13468);
   U6610 : AOI221_X1 port map( B1 => registers_5_11_port, B2 => n16250, C1 => 
                           registers_59_11_port, C2 => n16247, A => n13474, ZN 
                           => n13471);
   U6611 : OAI22_X1 port map( A1 => n16244, A2 => n12602, B1 => n16241, B2 => 
                           n14918, ZN => n13474);
   U6612 : AOI221_X1 port map( B1 => registers_50_12_port, B2 => n16278, C1 => 
                           net227119, C2 => n16275, A => n13426, ZN => n13419);
   U6613 : OAI22_X1 port map( A1 => n16272, A2 => n12652, B1 => n16269, B2 => 
                           n14948, ZN => n13426);
   U6614 : AOI221_X1 port map( B1 => registers_5_12_port, B2 => n16251, C1 => 
                           registers_59_12_port, C2 => n16248, A => n13432, ZN 
                           => n13429);
   U6615 : OAI22_X1 port map( A1 => n16245, A2 => n12669, B1 => n16242, B2 => 
                           n14919, ZN => n13432);
   U6616 : AOI221_X1 port map( B1 => registers_50_13_port, B2 => n16278, C1 => 
                           net227137, C2 => n16275, A => n13384, ZN => n13377);
   U6617 : OAI22_X1 port map( A1 => n16272, A2 => n13996, B1 => n16269, B2 => 
                           n14949, ZN => n13384);
   U6618 : AOI221_X1 port map( B1 => registers_5_13_port, B2 => n16251, C1 => 
                           registers_59_13_port, C2 => n16248, A => n13390, ZN 
                           => n13387);
   U6619 : OAI22_X1 port map( A1 => n16245, A2 => n13999, B1 => n16242, B2 => 
                           n14920, ZN => n13390);
   U6620 : AOI221_X1 port map( B1 => registers_50_14_port, B2 => n16278, C1 => 
                           net227155, C2 => n16275, A => n13342, ZN => n13335);
   U6621 : OAI22_X1 port map( A1 => n16272, A2 => n14008, B1 => n16269, B2 => 
                           n14950, ZN => n13342);
   U6622 : AOI221_X1 port map( B1 => registers_5_14_port, B2 => n16251, C1 => 
                           registers_59_14_port, C2 => n16248, A => n13348, ZN 
                           => n13345);
   U6623 : OAI22_X1 port map( A1 => n16245, A2 => n14014, B1 => n16242, B2 => 
                           n14921, ZN => n13348);
   U6624 : AOI221_X1 port map( B1 => registers_50_15_port, B2 => n16278, C1 => 
                           net227173, C2 => n16275, A => n13300, ZN => n13293);
   U6625 : OAI22_X1 port map( A1 => n16272, A2 => n14015, B1 => n16269, B2 => 
                           n14951, ZN => n13300);
   U6626 : AOI221_X1 port map( B1 => registers_5_15_port, B2 => n16251, C1 => 
                           registers_59_15_port, C2 => n16248, A => n13306, ZN 
                           => n13303);
   U6627 : OAI22_X1 port map( A1 => n16245, A2 => n14032, B1 => n16242, B2 => 
                           n14922, ZN => n13306);
   U6628 : AOI221_X1 port map( B1 => registers_50_16_port, B2 => n16278, C1 => 
                           net227191, C2 => n16275, A => n13258, ZN => n13251);
   U6629 : OAI22_X1 port map( A1 => n16272, A2 => n14035, B1 => n16269, B2 => 
                           n14952, ZN => n13258);
   U6630 : AOI221_X1 port map( B1 => registers_5_16_port, B2 => n16251, C1 => 
                           registers_59_16_port, C2 => n16248, A => n13264, ZN 
                           => n13261);
   U6631 : OAI22_X1 port map( A1 => n16245, A2 => n14036, B1 => n16242, B2 => 
                           n14923, ZN => n13264);
   U6632 : AOI221_X1 port map( B1 => registers_50_17_port, B2 => n16278, C1 => 
                           net227209, C2 => n16275, A => n13216, ZN => n13209);
   U6633 : OAI22_X1 port map( A1 => n16272, A2 => n14037, B1 => n16269, B2 => 
                           n14953, ZN => n13216);
   U6634 : AOI221_X1 port map( B1 => registers_5_17_port, B2 => n16251, C1 => 
                           registers_59_17_port, C2 => n16248, A => n13222, ZN 
                           => n13219);
   U6635 : OAI22_X1 port map( A1 => n16245, A2 => n14038, B1 => n16242, B2 => 
                           n14924, ZN => n13222);
   U6636 : AOI221_X1 port map( B1 => registers_50_18_port, B2 => n16278, C1 => 
                           net227227, C2 => n16275, A => n13174, ZN => n13167);
   U6637 : OAI22_X1 port map( A1 => n16272, A2 => n14039, B1 => n16269, B2 => 
                           n14954, ZN => n13174);
   U6638 : AOI221_X1 port map( B1 => registers_5_18_port, B2 => n16251, C1 => 
                           registers_59_18_port, C2 => n16248, A => n13180, ZN 
                           => n13177);
   U6639 : OAI22_X1 port map( A1 => n16245, A2 => n14040, B1 => n16242, B2 => 
                           n14925, ZN => n13180);
   U6640 : AOI221_X1 port map( B1 => registers_50_19_port, B2 => n16278, C1 => 
                           net227245, C2 => n16275, A => n13132, ZN => n13125);
   U6641 : OAI22_X1 port map( A1 => n16272, A2 => n14041, B1 => n16269, B2 => 
                           n14955, ZN => n13132);
   U6642 : AOI221_X1 port map( B1 => registers_5_19_port, B2 => n16251, C1 => 
                           registers_59_19_port, C2 => n16248, A => n13138, ZN 
                           => n13135);
   U6643 : OAI22_X1 port map( A1 => n16245, A2 => n14042, B1 => n16242, B2 => 
                           n14926, ZN => n13138);
   U6644 : AOI221_X1 port map( B1 => registers_50_20_port, B2 => n16278, C1 => 
                           net227263, C2 => n16275, A => n13090, ZN => n13083);
   U6645 : OAI22_X1 port map( A1 => n16272, A2 => n14043, B1 => n16269, B2 => 
                           n14956, ZN => n13090);
   U6646 : AOI221_X1 port map( B1 => registers_5_20_port, B2 => n16251, C1 => 
                           registers_59_20_port, C2 => n16248, A => n13096, ZN 
                           => n13093);
   U6647 : OAI22_X1 port map( A1 => n16245, A2 => n14044, B1 => n16242, B2 => 
                           n14927, ZN => n13096);
   U6648 : AOI221_X1 port map( B1 => registers_50_21_port, B2 => n16278, C1 => 
                           net227281, C2 => n16275, A => n13048, ZN => n13041);
   U6649 : OAI22_X1 port map( A1 => n16272, A2 => n14045, B1 => n16269, B2 => 
                           n14957, ZN => n13048);
   U6650 : AOI221_X1 port map( B1 => registers_5_21_port, B2 => n16251, C1 => 
                           registers_59_21_port, C2 => n16248, A => n13054, ZN 
                           => n13051);
   U6651 : OAI22_X1 port map( A1 => n16245, A2 => n14046, B1 => n16242, B2 => 
                           n14928, ZN => n13054);
   U6652 : AOI221_X1 port map( B1 => registers_50_22_port, B2 => n16278, C1 => 
                           net227299, C2 => n16275, A => n13006, ZN => n12999);
   U6653 : OAI22_X1 port map( A1 => n16272, A2 => n14047, B1 => n16269, B2 => 
                           n14958, ZN => n13006);
   U6654 : AOI221_X1 port map( B1 => registers_5_22_port, B2 => n16251, C1 => 
                           registers_59_22_port, C2 => n16248, A => n13012, ZN 
                           => n13009);
   U6655 : OAI22_X1 port map( A1 => n16245, A2 => n14048, B1 => n16242, B2 => 
                           n14929, ZN => n13012);
   U6656 : AOI221_X1 port map( B1 => registers_50_23_port, B2 => n16278, C1 => 
                           net227317, C2 => n16275, A => n12964, ZN => n12957);
   U6657 : OAI22_X1 port map( A1 => n16272, A2 => n14049, B1 => n16269, B2 => 
                           n14959, ZN => n12964);
   U6658 : AOI221_X1 port map( B1 => registers_5_23_port, B2 => n16251, C1 => 
                           registers_59_23_port, C2 => n16248, A => n12970, ZN 
                           => n12967);
   U6659 : OAI22_X1 port map( A1 => n16245, A2 => n14050, B1 => n16242, B2 => 
                           n14930, ZN => n12970);
   U6660 : AOI221_X1 port map( B1 => registers_49_0_port, B2 => n16541, C1 => 
                           registers_51_0_port, C2 => n16538, A => n12476, ZN 
                           => n12468);
   U6661 : OAI22_X1 port map( A1 => n16535, A2 => n15521, B1 => n16532, B2 => 
                           n14547, ZN => n12476);
   U6662 : AOI221_X1 port map( B1 => registers_49_1_port, B2 => n16541, C1 => 
                           registers_51_1_port, C2 => n16538, A => n12291, ZN 
                           => n12286);
   U6663 : OAI22_X1 port map( A1 => n16535, A2 => n15522, B1 => n16532, B2 => 
                           n14548, ZN => n12291);
   U6664 : AOI221_X1 port map( B1 => registers_49_2_port, B2 => n16541, C1 => 
                           registers_51_2_port, C2 => n16538, A => n12138, ZN 
                           => n12133);
   U6665 : OAI22_X1 port map( A1 => n16535, A2 => n15523, B1 => n16532, B2 => 
                           n14549, ZN => n12138);
   U6666 : AOI221_X1 port map( B1 => registers_49_3_port, B2 => n16541, C1 => 
                           registers_51_3_port, C2 => n16538, A => n11985, ZN 
                           => n11980);
   U6667 : OAI22_X1 port map( A1 => n16535, A2 => n15524, B1 => n16532, B2 => 
                           n14536, ZN => n11985);
   U6668 : AOI221_X1 port map( B1 => registers_49_4_port, B2 => n16541, C1 => 
                           registers_51_4_port, C2 => n16538, A => n11832, ZN 
                           => n11827);
   U6669 : OAI22_X1 port map( A1 => n16535, A2 => n15525, B1 => n16532, B2 => 
                           n14550, ZN => n11832);
   U6670 : AOI221_X1 port map( B1 => registers_49_5_port, B2 => n16541, C1 => 
                           registers_51_5_port, C2 => n16538, A => n11789, ZN 
                           => n11784);
   U6671 : OAI22_X1 port map( A1 => n16535, A2 => n15526, B1 => n16532, B2 => 
                           n14537, ZN => n11789);
   U6672 : AOI221_X1 port map( B1 => registers_49_6_port, B2 => n16541, C1 => 
                           registers_51_6_port, C2 => n16538, A => n11746, ZN 
                           => n11741);
   U6673 : OAI22_X1 port map( A1 => n16535, A2 => n15527, B1 => n16532, B2 => 
                           n14551, ZN => n11746);
   U6674 : AOI221_X1 port map( B1 => registers_49_7_port, B2 => n16541, C1 => 
                           registers_51_7_port, C2 => n16538, A => n11703, ZN 
                           => n11698);
   U6675 : OAI22_X1 port map( A1 => n16535, A2 => n15528, B1 => n16532, B2 => 
                           n14552, ZN => n11703);
   U6676 : AOI221_X1 port map( B1 => registers_49_8_port, B2 => n16541, C1 => 
                           registers_51_8_port, C2 => n16538, A => n11660, ZN 
                           => n11655);
   U6677 : OAI22_X1 port map( A1 => n16535, A2 => n15529, B1 => n16532, B2 => 
                           n14553, ZN => n11660);
   U6678 : AOI221_X1 port map( B1 => registers_49_9_port, B2 => n16541, C1 => 
                           registers_51_9_port, C2 => n16538, A => n11617, ZN 
                           => n11612);
   U6679 : OAI22_X1 port map( A1 => n16535, A2 => n15530, B1 => n16532, B2 => 
                           n14554, ZN => n11617);
   U6680 : AOI221_X1 port map( B1 => registers_49_10_port, B2 => n16541, C1 => 
                           registers_51_10_port, C2 => n16538, A => n11574, ZN 
                           => n11569);
   U6681 : OAI22_X1 port map( A1 => n16535, A2 => n15531, B1 => n16532, B2 => 
                           n14555, ZN => n11574);
   U6682 : AOI221_X1 port map( B1 => registers_49_11_port, B2 => n16541, C1 => 
                           registers_51_11_port, C2 => n16538, A => n11531, ZN 
                           => n11526);
   U6683 : OAI22_X1 port map( A1 => n16535, A2 => n15532, B1 => n16532, B2 => 
                           n14556, ZN => n11531);
   U6684 : AOI221_X1 port map( B1 => registers_49_12_port, B2 => n16542, C1 => 
                           registers_51_12_port, C2 => n16539, A => n11488, ZN 
                           => n11483);
   U6685 : OAI22_X1 port map( A1 => n16536, A2 => n15533, B1 => n16533, B2 => 
                           n14557, ZN => n11488);
   U6686 : AOI221_X1 port map( B1 => registers_49_13_port, B2 => n16542, C1 => 
                           registers_51_13_port, C2 => n16539, A => n11444, ZN 
                           => n11439);
   U6687 : OAI22_X1 port map( A1 => n16536, A2 => n15534, B1 => n16533, B2 => 
                           n14558, ZN => n11444);
   U6688 : AOI221_X1 port map( B1 => registers_49_14_port, B2 => n16542, C1 => 
                           registers_51_14_port, C2 => n16539, A => n11401, ZN 
                           => n11396);
   U6689 : OAI22_X1 port map( A1 => n16536, A2 => n15535, B1 => n16533, B2 => 
                           n14559, ZN => n11401);
   U6690 : AOI221_X1 port map( B1 => registers_49_15_port, B2 => n16542, C1 => 
                           registers_51_15_port, C2 => n16539, A => n11358, ZN 
                           => n11353);
   U6691 : OAI22_X1 port map( A1 => n16536, A2 => n15536, B1 => n16533, B2 => 
                           n14560, ZN => n11358);
   U6692 : AOI221_X1 port map( B1 => registers_49_16_port, B2 => n16542, C1 => 
                           registers_51_16_port, C2 => n16539, A => n11315, ZN 
                           => n11310);
   U6693 : OAI22_X1 port map( A1 => n16536, A2 => n15537, B1 => n16533, B2 => 
                           n14561, ZN => n11315);
   U6694 : AOI221_X1 port map( B1 => registers_49_17_port, B2 => n16542, C1 => 
                           registers_51_17_port, C2 => n16539, A => n11272, ZN 
                           => n11267);
   U6695 : OAI22_X1 port map( A1 => n16536, A2 => n15538, B1 => n16533, B2 => 
                           n14562, ZN => n11272);
   U6696 : AOI221_X1 port map( B1 => registers_49_18_port, B2 => n16542, C1 => 
                           registers_51_18_port, C2 => n16539, A => n11229, ZN 
                           => n11224);
   U6697 : OAI22_X1 port map( A1 => n16536, A2 => n15539, B1 => n16533, B2 => 
                           n14563, ZN => n11229);
   U6698 : AOI221_X1 port map( B1 => registers_49_19_port, B2 => n16542, C1 => 
                           registers_51_19_port, C2 => n16539, A => n11186, ZN 
                           => n11181);
   U6699 : OAI22_X1 port map( A1 => n16536, A2 => n15540, B1 => n16533, B2 => 
                           n14564, ZN => n11186);
   U6700 : AOI221_X1 port map( B1 => registers_49_20_port, B2 => n16542, C1 => 
                           registers_51_20_port, C2 => n16539, A => n11143, ZN 
                           => n11138);
   U6701 : OAI22_X1 port map( A1 => n16536, A2 => n15541, B1 => n16533, B2 => 
                           n14565, ZN => n11143);
   U6702 : AOI221_X1 port map( B1 => registers_49_21_port, B2 => n16542, C1 => 
                           registers_51_21_port, C2 => n16539, A => n11100, ZN 
                           => n11095);
   U6703 : OAI22_X1 port map( A1 => n16536, A2 => n15542, B1 => n16533, B2 => 
                           n14566, ZN => n11100);
   U6704 : AOI221_X1 port map( B1 => registers_49_22_port, B2 => n16542, C1 => 
                           registers_51_22_port, C2 => n16539, A => n11057, ZN 
                           => n11052);
   U6705 : OAI22_X1 port map( A1 => n16536, A2 => n15543, B1 => n16533, B2 => 
                           n14567, ZN => n11057);
   U6706 : AOI221_X1 port map( B1 => registers_49_23_port, B2 => n16542, C1 => 
                           registers_51_23_port, C2 => n16539, A => n11014, ZN 
                           => n11009);
   U6707 : OAI22_X1 port map( A1 => n16536, A2 => n15544, B1 => n16533, B2 => 
                           n14568, ZN => n11014);
   U6708 : AOI221_X1 port map( B1 => net226841, B2 => n17697, C1 => 
                           registers_9_0_port, C2 => n17694, A => n12397, ZN =>
                           n12392);
   U6709 : OAI22_X1 port map( A1 => n17691, A2 => n15758, B1 => n17688, B2 => 
                           n12171, ZN => n12397);
   U6710 : AOI221_X1 port map( B1 => net226864, B2 => n17697, C1 => 
                           registers_9_1_port, C2 => n17694, A => n12243, ZN =>
                           n12238);
   U6711 : OAI22_X1 port map( A1 => n17691, A2 => n15759, B1 => n17688, B2 => 
                           n12172, ZN => n12243);
   U6712 : AOI221_X1 port map( B1 => net226882, B2 => n17697, C1 => 
                           registers_9_2_port, C2 => n17694, A => n12088, ZN =>
                           n12083);
   U6713 : OAI22_X1 port map( A1 => n17691, A2 => n15760, B1 => n17688, B2 => 
                           n12173, ZN => n12088);
   U6714 : AOI221_X1 port map( B1 => net226902, B2 => n17697, C1 => 
                           registers_9_3_port, C2 => n17694, A => n11935, ZN =>
                           n11930);
   U6715 : OAI22_X1 port map( A1 => n17691, A2 => n15761, B1 => n17688, B2 => 
                           n12174, ZN => n11935);
   U6716 : AOI221_X1 port map( B1 => net226975, B2 => n17697, C1 => 
                           registers_9_4_port, C2 => n17694, A => n10492, ZN =>
                           n10487);
   U6717 : OAI22_X1 port map( A1 => n17691, A2 => n15762, B1 => n17688, B2 => 
                           n12175, ZN => n10492);
   U6718 : AOI221_X1 port map( B1 => net226995, B2 => n17697, C1 => 
                           registers_9_5_port, C2 => n17694, A => n10382, ZN =>
                           n10377);
   U6719 : OAI22_X1 port map( A1 => n17691, A2 => n15763, B1 => n17688, B2 => 
                           n12162, ZN => n10382);
   U6720 : AOI221_X1 port map( B1 => net227019, B2 => n17697, C1 => 
                           registers_9_6_port, C2 => n17694, A => n10270, ZN =>
                           n10265);
   U6721 : OAI22_X1 port map( A1 => n17691, A2 => n15764, B1 => n17688, B2 => 
                           n12176, ZN => n10270);
   U6722 : AOI221_X1 port map( B1 => net227037, B2 => n17697, C1 => 
                           registers_9_7_port, C2 => n17694, A => n7634, ZN => 
                           n7629);
   U6723 : OAI22_X1 port map( A1 => n17691, A2 => n15765, B1 => n17688, B2 => 
                           n12177, ZN => n7634);
   U6724 : AOI221_X1 port map( B1 => net227055, B2 => n17697, C1 => 
                           registers_9_8_port, C2 => n17694, A => n7519, ZN => 
                           n7514);
   U6725 : OAI22_X1 port map( A1 => n17691, A2 => n15766, B1 => n17688, B2 => 
                           n12178, ZN => n7519);
   U6726 : AOI221_X1 port map( B1 => net227073, B2 => n17697, C1 => 
                           registers_9_9_port, C2 => n17694, A => n7410, ZN => 
                           n7405);
   U6727 : OAI22_X1 port map( A1 => n17691, A2 => n15767, B1 => n17688, B2 => 
                           n12179, ZN => n7410);
   U6728 : AOI221_X1 port map( B1 => net227091, B2 => n17697, C1 => 
                           registers_9_10_port, C2 => n17694, A => n7301, ZN =>
                           n7296);
   U6729 : OAI22_X1 port map( A1 => n17691, A2 => n15768, B1 => n17688, B2 => 
                           n12180, ZN => n7301);
   U6730 : AOI221_X1 port map( B1 => net227109, B2 => n17698, C1 => 
                           registers_9_11_port, C2 => n17695, A => n7187, ZN =>
                           n7182);
   U6731 : OAI22_X1 port map( A1 => n17692, A2 => n15769, B1 => n17689, B2 => 
                           n12181, ZN => n7187);
   U6732 : AOI221_X1 port map( B1 => net227127, B2 => n17698, C1 => 
                           registers_9_12_port, C2 => n17695, A => n7078, ZN =>
                           n7073);
   U6733 : OAI22_X1 port map( A1 => n17692, A2 => n15770, B1 => n17689, B2 => 
                           n12182, ZN => n7078);
   U6734 : AOI221_X1 port map( B1 => net227145, B2 => n17698, C1 => 
                           registers_9_13_port, C2 => n17695, A => n6969, ZN =>
                           n6964);
   U6735 : OAI22_X1 port map( A1 => n17692, A2 => n15771, B1 => n17689, B2 => 
                           n12183, ZN => n6969);
   U6736 : AOI221_X1 port map( B1 => net227163, B2 => n17698, C1 => 
                           registers_9_14_port, C2 => n17695, A => n6860, ZN =>
                           n6855);
   U6737 : OAI22_X1 port map( A1 => n17692, A2 => n15772, B1 => n17689, B2 => 
                           n12185, ZN => n6860);
   U6738 : AOI221_X1 port map( B1 => net227181, B2 => n17698, C1 => 
                           registers_9_15_port, C2 => n17695, A => n6751, ZN =>
                           n6746);
   U6739 : OAI22_X1 port map( A1 => n17692, A2 => n15773, B1 => n17689, B2 => 
                           n12186, ZN => n6751);
   U6740 : AOI221_X1 port map( B1 => net227199, B2 => n17698, C1 => 
                           registers_9_16_port, C2 => n17695, A => n6609, ZN =>
                           n6603);
   U6741 : OAI22_X1 port map( A1 => n17692, A2 => n15774, B1 => n17689, B2 => 
                           n12187, ZN => n6609);
   U6742 : AOI221_X1 port map( B1 => net227217, B2 => n17698, C1 => 
                           registers_9_17_port, C2 => n17695, A => n6423, ZN =>
                           n6416);
   U6743 : OAI22_X1 port map( A1 => n17692, A2 => n15775, B1 => n17689, B2 => 
                           n12188, ZN => n6423);
   U6744 : AOI221_X1 port map( B1 => net227235, B2 => n17698, C1 => 
                           registers_9_18_port, C2 => n17695, A => n6237, ZN =>
                           n6229);
   U6745 : OAI22_X1 port map( A1 => n17692, A2 => n15776, B1 => n17689, B2 => 
                           n12189, ZN => n6237);
   U6746 : AOI221_X1 port map( B1 => net227253, B2 => n17698, C1 => 
                           registers_9_19_port, C2 => n17695, A => n6050, ZN =>
                           n6043);
   U6747 : OAI22_X1 port map( A1 => n17692, A2 => n15777, B1 => n17689, B2 => 
                           n12190, ZN => n6050);
   U6748 : AOI221_X1 port map( B1 => net227271, B2 => n17698, C1 => 
                           registers_9_20_port, C2 => n17695, A => n5863, ZN =>
                           n5858);
   U6749 : OAI22_X1 port map( A1 => n17692, A2 => n15778, B1 => n17689, B2 => 
                           n12191, ZN => n5863);
   U6750 : AOI221_X1 port map( B1 => net227289, B2 => n17698, C1 => 
                           registers_9_21_port, C2 => n17695, A => n5678, ZN =>
                           n5671);
   U6751 : OAI22_X1 port map( A1 => n17692, A2 => n15779, B1 => n17689, B2 => 
                           n12192, ZN => n5678);
   U6752 : AOI221_X1 port map( B1 => net227307, B2 => n17698, C1 => 
                           registers_9_22_port, C2 => n17695, A => n5492, ZN =>
                           n5484);
   U6753 : OAI22_X1 port map( A1 => n17692, A2 => n15780, B1 => n17689, B2 => 
                           n12193, ZN => n5492);
   U6754 : AOI221_X1 port map( B1 => net227469, B2 => n17697, C1 => 
                           registers_9_31_port, C2 => n17694, A => n14168, ZN 
                           => n14154);
   U6755 : OAI22_X1 port map( A1 => n17691, A2 => n15781, B1 => n17688, B2 => 
                           n12194, ZN => n14168);
   U6756 : NOR3_X1 port map( A1 => n13994, A2 => n12514, A3 => n13995, ZN => 
                           n13993);
   U6757 : XNOR2_X1 port map( A => n13984, B => add_wr(2), ZN => n13994);
   U6758 : NOR3_X1 port map( A1 => n12513, A2 => n12514, A3 => n12515, ZN => 
                           n12512);
   U6759 : XNOR2_X1 port map( A => n12503, B => add_wr(2), ZN => n12513);
   U6760 : NOR3_X1 port map( A1 => n14030, A2 => n14031, A3 => n17824, ZN => 
                           n14029);
   U6761 : XNOR2_X1 port map( A => swp_1_port, B => n10189, ZN => n14031);
   U6762 : XNOR2_X1 port map( A => swp_4_port, B => n14820, ZN => n14030);
   U6763 : NOR2_X1 port map( A1 => n10190, A2 => n10188, ZN => n14016);
   U6764 : NOR2_X1 port map( A1 => n13986, A2 => add_rd2(0), ZN => n13904);
   U6765 : INV_X1 port map( A => n13987, ZN => n13986);
   U6766 : NOR2_X1 port map( A1 => n12505, A2 => add_rd1(0), ZN => n12423);
   U6767 : INV_X1 port map( A => n12506, ZN => n12505);
   U6768 : NOR2_X1 port map( A1 => add_rd2(2), A2 => add_rd2(1), ZN => n13985);
   U6769 : NOR2_X1 port map( A1 => add_rd1(2), A2 => add_rd1(1), ZN => n12504);
   U6770 : OAI22_X1 port map( A1 => n17557, A2 => n16199, B1 => n16439, B2 => 
                           n17548, ZN => n7797);
   U6771 : OAI22_X1 port map( A1 => n17612, A2 => n16111, B1 => n16439, B2 => 
                           n17603, ZN => n7799);
   U6772 : OAI22_X1 port map( A1 => n16875, A2 => n15911, B1 => n16439, B2 => 
                           n16866, ZN => n7805);
   U6773 : OAI22_X1 port map( A1 => n17159, A2 => n15791, B1 => n16440, B2 => 
                           n17150, ZN => n7817);
   U6774 : OAI22_X1 port map( A1 => n17225, A2 => n15881, B1 => n16441, B2 => 
                           n17216, ZN => n7820);
   U6775 : OAI22_X1 port map( A1 => n17277, A2 => n15792, B1 => n16441, B2 => 
                           n17268, ZN => n7822);
   U6776 : OAI22_X1 port map( A1 => n17543, A2 => n16115, B1 => n16445, B2 => 
                           n17534, ZN => n7834);
   U6777 : OAI22_X1 port map( A1 => n17598, A2 => n16116, B1 => n16445, B2 => 
                           n17589, ZN => n7873);
   U6778 : OAI22_X1 port map( A1 => n16909, A2 => n15969, B1 => n16445, B2 => 
                           n16900, ZN => n7881);
   U6779 : OAI22_X1 port map( A1 => n16998, A2 => n15912, B1 => n16446, B2 => 
                           n16989, ZN => n7885);
   U6780 : OAI22_X1 port map( A1 => n17225, A2 => n15882, B1 => n16447, B2 => 
                           n17216, ZN => n7894);
   U6781 : OAI22_X1 port map( A1 => n17277, A2 => n15793, B1 => n16447, B2 => 
                           n17268, ZN => n7896);
   U6782 : OAI22_X1 port map( A1 => n17543, A2 => n16117, B1 => n16451, B2 => 
                           n17534, ZN => n7908);
   U6783 : OAI22_X1 port map( A1 => n17557, A2 => n16200, B1 => n16451, B2 => 
                           n17548, ZN => n7909);
   U6784 : OAI22_X1 port map( A1 => n17571, A2 => n16207, B1 => n16451, B2 => 
                           n17562, ZN => n7910);
   U6785 : OAI22_X1 port map( A1 => n16875, A2 => n15913, B1 => n16451, B2 => 
                           n16866, ZN => n7954);
   U6786 : OAI22_X1 port map( A1 => n17159, A2 => n15794, B1 => n16452, B2 => 
                           n17150, ZN => n7966);
   U6787 : OAI22_X1 port map( A1 => n17225, A2 => n15883, B1 => n16453, B2 => 
                           n17216, ZN => n7968);
   U6788 : OAI22_X1 port map( A1 => n17530, A2 => n15795, B1 => n17522, B2 => 
                           n16438, ZN => n7796);
   U6789 : OAI22_X1 port map( A1 => n17530, A2 => n15796, B1 => n17522, B2 => 
                           n16444, ZN => n7871);
   U6790 : OAI22_X1 port map( A1 => n17530, A2 => n15797, B1 => n17521, B2 => 
                           n16450, ZN => n7947);
   U6791 : OAI22_X1 port map( A1 => n17529, A2 => n15798, B1 => n17521, B2 => 
                           n16459, ZN => n8029);
   U6792 : OAI22_X1 port map( A1 => n17529, A2 => n15799, B1 => n17522, B2 => 
                           n16712, ZN => n8157);
   U6793 : OAI22_X1 port map( A1 => n17529, A2 => n15800, B1 => n17522, B2 => 
                           n16721, ZN => n8229);
   U6794 : OAI22_X1 port map( A1 => n17530, A2 => n15801, B1 => n17521, B2 => 
                           n16702, ZN => n10125);
   U6795 : OAI22_X1 port map( A1 => n17626, A2 => n16201, B1 => n17618, B2 => 
                           n16436, ZN => n7763);
   U6796 : OAI22_X1 port map( A1 => n17998, A2 => n15998, B1 => n17990, B2 => 
                           n16436, ZN => n7768);
   U6797 : OAI22_X1 port map( A1 => n17626, A2 => n16202, B1 => n17618, B2 => 
                           n16442, ZN => n7838);
   U6798 : OAI22_X1 port map( A1 => n17998, A2 => n15999, B1 => n17990, B2 => 
                           n16442, ZN => n7843);
   U6799 : OAI22_X1 port map( A1 => n17626, A2 => n16203, B1 => n17618, B2 => 
                           n16448, ZN => n7914);
   U6800 : OAI22_X1 port map( A1 => n17998, A2 => n16000, B1 => n17990, B2 => 
                           n16448, ZN => n7919);
   U6801 : OAI22_X1 port map( A1 => n17626, A2 => n16204, B1 => n17618, B2 => 
                           n16456, ZN => n7988);
   U6802 : OAI22_X1 port map( A1 => n17625, A2 => n16124, B1 => n17618, B2 => 
                           n16709, ZN => n8116);
   U6803 : OAI22_X1 port map( A1 => n17625, A2 => n16125, B1 => n17618, B2 => 
                           n16718, ZN => n8188);
   U6804 : OAI22_X1 port map( A1 => n17998, A2 => n16001, B1 => n17990, B2 => 
                           n16725, ZN => n8269);
   U6805 : OAI22_X1 port map( A1 => n17997, A2 => n16002, B1 => n17990, B2 => 
                           n16732, ZN => n8341);
   U6806 : OAI22_X1 port map( A1 => n17997, A2 => n16003, B1 => n17990, B2 => 
                           n16744, ZN => n8485);
   U6807 : OAI22_X1 port map( A1 => n17529, A2 => n15802, B1 => n17522, B2 => 
                           n16730, ZN => n8325);
   U6808 : OAI22_X1 port map( A1 => n16875, A2 => n15914, B1 => n16867, B2 => 
                           n16442, ZN => n7844);
   U6809 : OAI22_X1 port map( A1 => n16874, A2 => n15915, B1 => n16867, B2 => 
                           n16456, ZN => n7992);
   U6810 : OAI22_X1 port map( A1 => n16874, A2 => n15916, B1 => n16867, B2 => 
                           n16725, ZN => n8272);
   U6811 : OAI22_X1 port map( A1 => n16874, A2 => n15917, B1 => n16867, B2 => 
                           n16732, ZN => n8344);
   U6812 : OAI22_X1 port map( A1 => n16874, A2 => n15918, B1 => n16867, B2 => 
                           n16738, ZN => n8416);
   U6813 : OAI22_X1 port map( A1 => n16873, A2 => n15919, B1 => n16867, B2 => 
                           n16744, ZN => n8488);
   U6814 : OAI22_X1 port map( A1 => n16875, A2 => n15920, B1 => n16867, B2 => 
                           n16706, ZN => n10072);
   U6815 : OAI22_X1 port map( A1 => n16909, A2 => n15970, B1 => n16901, B2 => 
                           n16436, ZN => n7771);
   U6816 : OAI22_X1 port map( A1 => n16998, A2 => n15921, B1 => n16990, B2 => 
                           n16437, ZN => n7775);
   U6817 : OAI22_X1 port map( A1 => n17159, A2 => n15803, B1 => n17151, B2 => 
                           n16443, ZN => n7856);
   U6818 : OAI22_X1 port map( A1 => n16909, A2 => n15971, B1 => n16901, B2 => 
                           n16448, ZN => n7921);
   U6819 : OAI22_X1 port map( A1 => n16998, A2 => n15922, B1 => n16990, B2 => 
                           n16449, ZN => n7925);
   U6820 : OAI22_X1 port map( A1 => n17277, A2 => n15804, B1 => n17269, B2 => 
                           n16450, ZN => n7936);
   U6821 : OAI22_X1 port map( A1 => n16908, A2 => n15972, B1 => n16901, B2 => 
                           n16457, ZN => n7995);
   U6822 : OAI22_X1 port map( A1 => n17224, A2 => n15884, B1 => n17217, B2 => 
                           n16458, ZN => n8006);
   U6823 : OAI22_X1 port map( A1 => n17276, A2 => n15805, B1 => n17269, B2 => 
                           n16458, ZN => n8010);
   U6824 : OAI22_X1 port map( A1 => n16997, A2 => n15923, B1 => n16990, B2 => 
                           n16710, ZN => n8123);
   U6825 : OAI22_X1 port map( A1 => n17158, A2 => n15806, B1 => n17151, B2 => 
                           n16718, ZN => n8200);
   U6826 : OAI22_X1 port map( A1 => n17224, A2 => n15885, B1 => n17217, B2 => 
                           n16719, ZN => n8206);
   U6827 : OAI22_X1 port map( A1 => n17276, A2 => n15807, B1 => n17269, B2 => 
                           n16719, ZN => n8210);
   U6828 : OAI22_X1 port map( A1 => n16908, A2 => n15973, B1 => n16901, B2 => 
                           n16726, ZN => n8275);
   U6829 : OAI22_X1 port map( A1 => n16997, A2 => n15924, B1 => n16990, B2 => 
                           n16726, ZN => n8283);
   U6830 : OAI22_X1 port map( A1 => n17158, A2 => n15808, B1 => n17151, B2 => 
                           n16727, ZN => n8296);
   U6831 : OAI22_X1 port map( A1 => n17224, A2 => n15886, B1 => n17217, B2 => 
                           n16728, ZN => n8302);
   U6832 : OAI22_X1 port map( A1 => n17276, A2 => n15809, B1 => n17269, B2 => 
                           n16728, ZN => n8306);
   U6833 : OAI22_X1 port map( A1 => n16908, A2 => n15974, B1 => n16901, B2 => 
                           n16732, ZN => n8347);
   U6834 : OAI22_X1 port map( A1 => n16997, A2 => n15925, B1 => n16990, B2 => 
                           n16733, ZN => n8355);
   U6835 : OAI22_X1 port map( A1 => n17158, A2 => n15810, B1 => n17151, B2 => 
                           n16734, ZN => n8368);
   U6836 : OAI22_X1 port map( A1 => n17224, A2 => n15887, B1 => n17217, B2 => 
                           n16735, ZN => n8374);
   U6837 : OAI22_X1 port map( A1 => n17276, A2 => n15811, B1 => n17269, B2 => 
                           n16735, ZN => n8378);
   U6838 : OAI22_X1 port map( A1 => n17158, A2 => n15812, B1 => n17151, B2 => 
                           n16740, ZN => n8440);
   U6839 : OAI22_X1 port map( A1 => n17223, A2 => n15888, B1 => n17217, B2 => 
                           n16741, ZN => n8446);
   U6840 : OAI22_X1 port map( A1 => n16909, A2 => n15975, B1 => n16901, B2 => 
                           n16706, ZN => n10075);
   U6841 : OAI22_X1 port map( A1 => n16998, A2 => n15926, B1 => n16990, B2 => 
                           n16706, ZN => n10083);
   U6842 : OAI22_X1 port map( A1 => n17159, A2 => n15813, B1 => n17151, B2 => 
                           n16704, ZN => n10096);
   U6843 : OAI22_X1 port map( A1 => n17225, A2 => n15889, B1 => n17217, B2 => 
                           n16704, ZN => n10102);
   U6844 : OAI22_X1 port map( A1 => n17277, A2 => n15814, B1 => n17269, B2 => 
                           n16704, ZN => n10106);
   U6845 : OAI22_X1 port map( A1 => n17543, A2 => n16118, B1 => n17535, B2 => 
                           n16436, ZN => n7760);
   U6846 : OAI22_X1 port map( A1 => n17542, A2 => n16119, B1 => n17535, B2 => 
                           n16456, ZN => n7982);
   U6847 : OAI22_X1 port map( A1 => n17542, A2 => n16036, B1 => n17535, B2 => 
                           n16709, ZN => n8110);
   U6848 : OAI22_X1 port map( A1 => n17542, A2 => n16037, B1 => n17535, B2 => 
                           n16718, ZN => n8182);
   U6849 : OAI22_X1 port map( A1 => n17542, A2 => n16038, B1 => n17535, B2 => 
                           n16731, ZN => n8326);
   U6850 : OAI22_X1 port map( A1 => n17541, A2 => n16039, B1 => n17535, B2 => 
                           n16737, ZN => n8398);
   U6851 : OAI22_X1 port map( A1 => n17571, A2 => n16208, B1 => n17563, B2 => 
                           n16436, ZN => n7761);
   U6852 : OAI22_X1 port map( A1 => n17598, A2 => n16120, B1 => n17590, B2 => 
                           n16436, ZN => n7762);
   U6853 : OAI22_X1 port map( A1 => n17557, A2 => n16205, B1 => n17549, B2 => 
                           n16442, ZN => n7835);
   U6854 : OAI22_X1 port map( A1 => n17571, A2 => n16209, B1 => n17563, B2 => 
                           n16442, ZN => n7836);
   U6855 : OAI22_X1 port map( A1 => n17612, A2 => n16112, B1 => n17604, B2 => 
                           n16442, ZN => n7837);
   U6856 : OAI22_X1 port map( A1 => n17598, A2 => n16121, B1 => n17590, B2 => 
                           n16448, ZN => n7912);
   U6857 : OAI22_X1 port map( A1 => n17612, A2 => n16113, B1 => n17604, B2 => 
                           n16448, ZN => n7913);
   U6858 : OAI22_X1 port map( A1 => n17557, A2 => n16206, B1 => n17549, B2 => 
                           n16456, ZN => n7983);
   U6859 : OAI22_X1 port map( A1 => n17571, A2 => n16210, B1 => n17563, B2 => 
                           n16456, ZN => n7984);
   U6860 : OAI22_X1 port map( A1 => n17598, A2 => n16122, B1 => n17590, B2 => 
                           n16456, ZN => n7986);
   U6861 : OAI22_X1 port map( A1 => n17612, A2 => n16114, B1 => n17604, B2 => 
                           n16456, ZN => n7987);
   U6862 : OAI22_X1 port map( A1 => n17556, A2 => n16126, B1 => n17549, B2 => 
                           n16709, ZN => n8111);
   U6863 : OAI22_X1 port map( A1 => n17570, A2 => n16174, B1 => n17563, B2 => 
                           n16709, ZN => n8112);
   U6864 : OAI22_X1 port map( A1 => n17597, A2 => n16040, B1 => n17590, B2 => 
                           n16709, ZN => n8114);
   U6865 : OAI22_X1 port map( A1 => n17611, A2 => n16086, B1 => n17604, B2 => 
                           n16709, ZN => n8115);
   U6866 : OAI22_X1 port map( A1 => n17556, A2 => n16127, B1 => n17549, B2 => 
                           n16718, ZN => n8183);
   U6867 : OAI22_X1 port map( A1 => n17570, A2 => n16175, B1 => n17563, B2 => 
                           n16718, ZN => n8184);
   U6868 : OAI22_X1 port map( A1 => n17597, A2 => n16041, B1 => n17590, B2 => 
                           n16718, ZN => n8186);
   U6869 : OAI22_X1 port map( A1 => n17611, A2 => n16087, B1 => n17604, B2 => 
                           n16718, ZN => n8187);
   U6870 : OAI22_X1 port map( A1 => n17556, A2 => n16128, B1 => n17549, B2 => 
                           n16731, ZN => n8327);
   U6871 : OAI22_X1 port map( A1 => n16908, A2 => n15976, B1 => n16901, B2 => 
                           n16738, ZN => n8419);
   U6872 : OAI22_X1 port map( A1 => n16997, A2 => n15927, B1 => n16990, B2 => 
                           n16739, ZN => n8427);
   U6873 : OAI22_X1 port map( A1 => n17275, A2 => n15815, B1 => n17269, B2 => 
                           n16741, ZN => n8450);
   U6874 : OAI22_X1 port map( A1 => n16907, A2 => n15977, B1 => n16901, B2 => 
                           n16744, ZN => n8491);
   U6875 : OAI22_X1 port map( A1 => n16996, A2 => n15928, B1 => n16990, B2 => 
                           n16745, ZN => n8499);
   U6876 : OAI22_X1 port map( A1 => n17157, A2 => n15816, B1 => n17151, B2 => 
                           n16746, ZN => n8512);
   U6877 : OAI22_X1 port map( A1 => n17223, A2 => n15890, B1 => n17217, B2 => 
                           n16747, ZN => n8518);
   U6878 : OAI22_X1 port map( A1 => n17275, A2 => n15817, B1 => n17269, B2 => 
                           n16747, ZN => n8522);
   U6879 : OAI22_X1 port map( A1 => n16907, A2 => n15978, B1 => n16901, B2 => 
                           n16750, ZN => n8563);
   U6880 : OAI22_X1 port map( A1 => n16996, A2 => n15929, B1 => n16990, B2 => 
                           n16751, ZN => n8571);
   U6881 : OAI22_X1 port map( A1 => n17157, A2 => n15818, B1 => n17151, B2 => 
                           n16752, ZN => n8584);
   U6882 : OAI22_X1 port map( A1 => n17223, A2 => n15891, B1 => n17217, B2 => 
                           n16753, ZN => n8590);
   U6883 : OAI22_X1 port map( A1 => n17275, A2 => n15819, B1 => n17269, B2 => 
                           n16753, ZN => n8594);
   U6884 : OAI22_X1 port map( A1 => n16907, A2 => n15979, B1 => n16901, B2 => 
                           n16756, ZN => n8635);
   U6885 : OAI22_X1 port map( A1 => n16996, A2 => n15930, B1 => n16990, B2 => 
                           n16757, ZN => n8643);
   U6886 : OAI22_X1 port map( A1 => n17157, A2 => n15820, B1 => n17151, B2 => 
                           n16758, ZN => n8656);
   U6887 : OAI22_X1 port map( A1 => n17223, A2 => n15892, B1 => n17217, B2 => 
                           n16759, ZN => n8662);
   U6888 : OAI22_X1 port map( A1 => n17275, A2 => n15821, B1 => n17269, B2 => 
                           n16759, ZN => n8666);
   U6889 : OAI22_X1 port map( A1 => n16907, A2 => n15980, B1 => n16901, B2 => 
                           n16762, ZN => n8707);
   U6890 : OAI22_X1 port map( A1 => n16996, A2 => n15931, B1 => n16990, B2 => 
                           n16763, ZN => n8715);
   U6891 : OAI22_X1 port map( A1 => n17157, A2 => n15822, B1 => n17151, B2 => 
                           n16764, ZN => n8728);
   U6892 : OAI22_X1 port map( A1 => n17222, A2 => n15893, B1 => n17217, B2 => 
                           n16765, ZN => n8734);
   U6893 : OAI22_X1 port map( A1 => n17274, A2 => n15823, B1 => n17269, B2 => 
                           n16765, ZN => n8738);
   U6894 : OAI22_X1 port map( A1 => n16906, A2 => n15981, B1 => n16901, B2 => 
                           n16768, ZN => n8779);
   U6895 : OAI22_X1 port map( A1 => n16995, A2 => n15932, B1 => n16990, B2 => 
                           n16769, ZN => n8787);
   U6896 : OAI22_X1 port map( A1 => n17156, A2 => n15824, B1 => n17151, B2 => 
                           n16770, ZN => n8800);
   U6897 : OAI22_X1 port map( A1 => n17222, A2 => n15894, B1 => n17217, B2 => 
                           n16771, ZN => n8806);
   U6898 : OAI22_X1 port map( A1 => n17274, A2 => n15825, B1 => n17269, B2 => 
                           n16771, ZN => n8810);
   U6899 : OAI22_X1 port map( A1 => n16906, A2 => n15982, B1 => n16901, B2 => 
                           n16774, ZN => n8851);
   U6900 : OAI22_X1 port map( A1 => n16995, A2 => n15933, B1 => n16990, B2 => 
                           n16775, ZN => n8859);
   U6901 : OAI22_X1 port map( A1 => n17156, A2 => n15826, B1 => n17151, B2 => 
                           n16776, ZN => n8872);
   U6902 : OAI22_X1 port map( A1 => n17222, A2 => n15895, B1 => n17217, B2 => 
                           n16777, ZN => n8878);
   U6903 : OAI22_X1 port map( A1 => n17274, A2 => n15827, B1 => n17269, B2 => 
                           n16777, ZN => n8882);
   U6904 : OAI22_X1 port map( A1 => n16906, A2 => n15983, B1 => n16901, B2 => 
                           n16780, ZN => n8923);
   U6905 : OAI22_X1 port map( A1 => n16995, A2 => n15934, B1 => n16990, B2 => 
                           n16781, ZN => n8931);
   U6906 : OAI22_X1 port map( A1 => n17156, A2 => n15828, B1 => n17151, B2 => 
                           n16782, ZN => n8944);
   U6907 : OAI22_X1 port map( A1 => n17221, A2 => n15896, B1 => n17217, B2 => 
                           n16783, ZN => n8950);
   U6908 : OAI22_X1 port map( A1 => n17273, A2 => n15829, B1 => n17269, B2 => 
                           n16783, ZN => n8954);
   U6909 : OAI22_X1 port map( A1 => n16905, A2 => n15984, B1 => n16901, B2 => 
                           n16786, ZN => n8995);
   U6910 : OAI22_X1 port map( A1 => n16994, A2 => n15935, B1 => n16990, B2 => 
                           n16787, ZN => n9003);
   U6911 : OAI22_X1 port map( A1 => n17155, A2 => n15830, B1 => n17151, B2 => 
                           n16788, ZN => n9016);
   U6912 : OAI22_X1 port map( A1 => n17221, A2 => n15897, B1 => n17217, B2 => 
                           n16789, ZN => n9022);
   U6913 : OAI22_X1 port map( A1 => n17273, A2 => n15831, B1 => n17269, B2 => 
                           n16789, ZN => n9026);
   U6914 : OAI22_X1 port map( A1 => n16905, A2 => n15985, B1 => n16901, B2 => 
                           n16792, ZN => n9067);
   U6915 : OAI22_X1 port map( A1 => n16994, A2 => n15936, B1 => n16990, B2 => 
                           n16793, ZN => n9075);
   U6916 : OAI22_X1 port map( A1 => n17155, A2 => n15832, B1 => n17151, B2 => 
                           n16794, ZN => n9088);
   U6917 : OAI22_X1 port map( A1 => n17221, A2 => n15898, B1 => n17217, B2 => 
                           n16795, ZN => n9094);
   U6918 : OAI22_X1 port map( A1 => n17273, A2 => n15833, B1 => n17269, B2 => 
                           n16795, ZN => n9098);
   U6919 : OAI22_X1 port map( A1 => n16905, A2 => n15986, B1 => n16901, B2 => 
                           n16798, ZN => n9139);
   U6920 : OAI22_X1 port map( A1 => n16994, A2 => n15937, B1 => n16990, B2 => 
                           n16799, ZN => n9147);
   U6921 : OAI22_X1 port map( A1 => n17155, A2 => n15834, B1 => n17151, B2 => 
                           n16800, ZN => n9160);
   U6922 : OAI22_X1 port map( A1 => n17221, A2 => n15899, B1 => n17217, B2 => 
                           n16801, ZN => n9166);
   U6923 : OAI22_X1 port map( A1 => n17273, A2 => n15835, B1 => n17269, B2 => 
                           n16801, ZN => n9170);
   U6924 : OAI22_X1 port map( A1 => n16905, A2 => n15987, B1 => n16901, B2 => 
                           n16804, ZN => n9211);
   U6925 : OAI22_X1 port map( A1 => n16994, A2 => n15938, B1 => n16990, B2 => 
                           n16805, ZN => n9219);
   U6926 : OAI22_X1 port map( A1 => n17155, A2 => n15836, B1 => n17151, B2 => 
                           n16806, ZN => n9232);
   U6927 : OAI22_X1 port map( A1 => n17220, A2 => n15900, B1 => n17217, B2 => 
                           n16807, ZN => n9238);
   U6928 : OAI22_X1 port map( A1 => n17272, A2 => n15837, B1 => n17269, B2 => 
                           n16807, ZN => n9242);
   U6929 : OAI22_X1 port map( A1 => n17154, A2 => n15838, B1 => n17151, B2 => 
                           n16812, ZN => n9304);
   U6930 : OAI22_X1 port map( A1 => n17220, A2 => n15901, B1 => n17217, B2 => 
                           n16813, ZN => n9310);
   U6931 : OAI22_X1 port map( A1 => n16906, A2 => n15988, B1 => n16901, B2 => 
                           n17513, ZN => n9931);
   U6932 : OAI22_X1 port map( A1 => n16995, A2 => n15939, B1 => n16990, B2 => 
                           n17514, ZN => n9939);
   U6933 : OAI22_X1 port map( A1 => n17156, A2 => n15839, B1 => n17151, B2 => 
                           n17515, ZN => n9952);
   U6934 : OAI22_X1 port map( A1 => n17222, A2 => n15902, B1 => n17217, B2 => 
                           n17516, ZN => n9958);
   U6935 : OAI22_X1 port map( A1 => n17274, A2 => n15840, B1 => n17269, B2 => 
                           n17516, ZN => n9962);
   U6936 : NAND2_X1 port map( A1 => add_wr(2), A2 => n14223, ZN => n12413);
   U6937 : OAI22_X1 port map( A1 => net227474, A2 => n14007, B1 => n14009, B2 
                           => n14012, ZN => n10136);
   U6938 : XNOR2_X1 port map( A => N9641, B => n10189, ZN => n14012);
   U6939 : OAI22_X1 port map( A1 => net227475, A2 => n14007, B1 => n14009, B2 
                           => n14010, ZN => n10137);
   U6940 : OAI22_X1 port map( A1 => n17220, A2 => n15903, B1 => n17216, B2 => 
                           n16819, ZN => n9382);
   U6941 : OAI22_X1 port map( A1 => n17220, A2 => n15904, B1 => n17216, B2 => 
                           n16825, ZN => n9454);
   U6942 : OAI22_X1 port map( A1 => n17219, A2 => n15905, B1 => n17216, B2 => 
                           n16831, ZN => n9526);
   U6943 : OAI22_X1 port map( A1 => n17219, A2 => n15906, B1 => n17216, B2 => 
                           n16837, ZN => n9598);
   U6944 : OAI22_X1 port map( A1 => n17219, A2 => n15907, B1 => n17216, B2 => 
                           n16843, ZN => n9670);
   U6945 : OAI22_X1 port map( A1 => n17219, A2 => n15908, B1 => n17216, B2 => 
                           n16849, ZN => n9742);
   U6946 : OAI22_X1 port map( A1 => n17218, A2 => n15909, B1 => n17216, B2 => 
                           n16855, ZN => n9814);
   U6947 : OAI22_X1 port map( A1 => n17218, A2 => n15910, B1 => n17216, B2 => 
                           n16861, ZN => n9886);
   U6948 : OAI22_X1 port map( A1 => n17154, A2 => n15841, B1 => n17150, B2 => 
                           n16818, ZN => n9376);
   U6949 : OAI22_X1 port map( A1 => n17154, A2 => n15842, B1 => n17150, B2 => 
                           n16824, ZN => n9448);
   U6950 : OAI22_X1 port map( A1 => n17153, A2 => n15843, B1 => n17150, B2 => 
                           n16830, ZN => n9520);
   U6951 : OAI22_X1 port map( A1 => n17154, A2 => n15844, B1 => n17150, B2 => 
                           n16836, ZN => n9592);
   U6952 : OAI22_X1 port map( A1 => n17153, A2 => n15845, B1 => n17150, B2 => 
                           n16842, ZN => n9664);
   U6953 : OAI22_X1 port map( A1 => n17153, A2 => n15846, B1 => n17150, B2 => 
                           n16848, ZN => n9736);
   U6954 : OAI22_X1 port map( A1 => n17153, A2 => n15847, B1 => n17150, B2 => 
                           n16854, ZN => n9808);
   U6955 : OAI22_X1 port map( A1 => n17152, A2 => n15848, B1 => n17150, B2 => 
                           n16860, ZN => n9880);
   U6956 : OAI22_X1 port map( A1 => n17272, A2 => n15849, B1 => n17268, B2 => 
                           n16813, ZN => n9314);
   U6957 : OAI22_X1 port map( A1 => n17272, A2 => n15850, B1 => n17268, B2 => 
                           n16819, ZN => n9386);
   U6958 : OAI22_X1 port map( A1 => n16870, A2 => n15940, B1 => n16866, B2 => 
                           n16822, ZN => n9424);
   U6959 : OAI22_X1 port map( A1 => n17272, A2 => n15851, B1 => n17268, B2 => 
                           n16825, ZN => n9458);
   U6960 : OAI22_X1 port map( A1 => n16870, A2 => n15941, B1 => n16866, B2 => 
                           n16828, ZN => n9496);
   U6961 : OAI22_X1 port map( A1 => n17271, A2 => n15852, B1 => n17268, B2 => 
                           n16831, ZN => n9530);
   U6962 : OAI22_X1 port map( A1 => n16869, A2 => n15942, B1 => n16866, B2 => 
                           n16834, ZN => n9568);
   U6963 : OAI22_X1 port map( A1 => n17271, A2 => n15853, B1 => n17268, B2 => 
                           n16837, ZN => n9602);
   U6964 : OAI22_X1 port map( A1 => n16869, A2 => n15943, B1 => n16866, B2 => 
                           n16840, ZN => n9640);
   U6965 : OAI22_X1 port map( A1 => n17271, A2 => n15854, B1 => n17268, B2 => 
                           n16843, ZN => n9674);
   U6966 : OAI22_X1 port map( A1 => n16869, A2 => n15944, B1 => n16866, B2 => 
                           n16846, ZN => n9712);
   U6967 : OAI22_X1 port map( A1 => n17271, A2 => n15855, B1 => n17268, B2 => 
                           n16849, ZN => n9746);
   U6968 : OAI22_X1 port map( A1 => n16869, A2 => n15945, B1 => n16866, B2 => 
                           n16852, ZN => n9784);
   U6969 : OAI22_X1 port map( A1 => n17270, A2 => n15856, B1 => n17268, B2 => 
                           n16855, ZN => n9818);
   U6970 : OAI22_X1 port map( A1 => n16868, A2 => n15946, B1 => n16866, B2 => 
                           n16858, ZN => n9856);
   U6971 : OAI22_X1 port map( A1 => n17270, A2 => n15857, B1 => n17268, B2 => 
                           n16861, ZN => n9890);
   U6972 : OAI22_X1 port map( A1 => n15782, A2 => n16868, B1 => n16866, B2 => 
                           n18031, ZN => n10000);
   U6973 : OAI22_X1 port map( A1 => n17552, A2 => n16129, B1 => n17548, B2 => 
                           n16809, ZN => n9263);
   U6974 : OAI22_X1 port map( A1 => n17538, A2 => n16042, B1 => n17534, B2 => 
                           n16815, ZN => n9334);
   U6975 : OAI22_X1 port map( A1 => n17552, A2 => n16130, B1 => n17548, B2 => 
                           n16815, ZN => n9335);
   U6976 : OAI22_X1 port map( A1 => n17537, A2 => n16043, B1 => n17534, B2 => 
                           n16827, ZN => n9478);
   U6977 : OAI22_X1 port map( A1 => n17552, A2 => n16131, B1 => n17548, B2 => 
                           n16827, ZN => n9479);
   U6978 : OAI22_X1 port map( A1 => n17537, A2 => n16044, B1 => n17534, B2 => 
                           n16833, ZN => n9550);
   U6979 : OAI22_X1 port map( A1 => n17551, A2 => n16132, B1 => n17548, B2 => 
                           n16833, ZN => n9551);
   U6980 : OAI22_X1 port map( A1 => n17538, A2 => n16045, B1 => n17534, B2 => 
                           n16839, ZN => n9622);
   U6981 : OAI22_X1 port map( A1 => n17552, A2 => n16133, B1 => n17548, B2 => 
                           n16839, ZN => n9623);
   U6982 : OAI22_X1 port map( A1 => n17537, A2 => n16046, B1 => n17534, B2 => 
                           n16845, ZN => n9694);
   U6983 : OAI22_X1 port map( A1 => n17551, A2 => n16134, B1 => n17548, B2 => 
                           n16845, ZN => n9695);
   U6984 : OAI22_X1 port map( A1 => n17536, A2 => n16047, B1 => n17534, B2 => 
                           n16851, ZN => n9766);
   U6985 : OAI22_X1 port map( A1 => n17551, A2 => n16135, B1 => n17548, B2 => 
                           n16851, ZN => n9767);
   U6986 : OAI22_X1 port map( A1 => n17537, A2 => n16048, B1 => n17534, B2 => 
                           n16857, ZN => n9838);
   U6987 : OAI22_X1 port map( A1 => n17551, A2 => n16136, B1 => n17548, B2 => 
                           n16857, ZN => n9839);
   U6988 : OAI22_X1 port map( A1 => n17536, A2 => n16049, B1 => n17534, B2 => 
                           n17512, ZN => n9910_port);
   U6989 : OAI22_X1 port map( A1 => n17550, A2 => n16137, B1 => n17548, B2 => 
                           n17512, ZN => n9911);
   U6990 : OAI22_X1 port map( A1 => n17543, A2 => n16123, B1 => n17534, B2 => 
                           n16702, ZN => n10054);
   U6991 : OAI22_X1 port map( A1 => n16904, A2 => n15989, B1 => n16900, B2 => 
                           n16810, ZN => n9283);
   U6992 : OAI22_X1 port map( A1 => n16993, A2 => n15947, B1 => n16989, B2 => 
                           n16811, ZN => n9291);
   U6993 : OAI22_X1 port map( A1 => n16904, A2 => n15990, B1 => n16900, B2 => 
                           n16816, ZN => n9355);
   U6994 : OAI22_X1 port map( A1 => n16993, A2 => n15948, B1 => n16989, B2 => 
                           n16817, ZN => n9363);
   U6995 : OAI22_X1 port map( A1 => n16904, A2 => n15991, B1 => n16900, B2 => 
                           n16822, ZN => n9427);
   U6996 : OAI22_X1 port map( A1 => n16993, A2 => n15949, B1 => n16989, B2 => 
                           n16823, ZN => n9435);
   U6997 : OAI22_X1 port map( A1 => n16904, A2 => n15992, B1 => n16900, B2 => 
                           n16828, ZN => n9499);
   U6998 : OAI22_X1 port map( A1 => n16992, A2 => n15950, B1 => n16989, B2 => 
                           n16829, ZN => n9507);
   U6999 : OAI22_X1 port map( A1 => n16903, A2 => n15993, B1 => n16900, B2 => 
                           n16834, ZN => n9571);
   U7000 : OAI22_X1 port map( A1 => n16993, A2 => n15951, B1 => n16989, B2 => 
                           n16835, ZN => n9579);
   U7001 : OAI22_X1 port map( A1 => n16903, A2 => n15994, B1 => n16900, B2 => 
                           n16840, ZN => n9643);
   U7002 : OAI22_X1 port map( A1 => n16992, A2 => n15952, B1 => n16989, B2 => 
                           n16841, ZN => n9651);
   U7003 : OAI22_X1 port map( A1 => n16903, A2 => n15995, B1 => n16900, B2 => 
                           n16846, ZN => n9715);
   U7004 : OAI22_X1 port map( A1 => n16992, A2 => n15953, B1 => n16989, B2 => 
                           n16847, ZN => n9723);
   U7005 : OAI22_X1 port map( A1 => n16903, A2 => n15996, B1 => n16900, B2 => 
                           n16852, ZN => n9787);
   U7006 : OAI22_X1 port map( A1 => n16992, A2 => n15954, B1 => n16989, B2 => 
                           n16853, ZN => n9795);
   U7007 : OAI22_X1 port map( A1 => n16902, A2 => n15997, B1 => n16900, B2 => 
                           n16858, ZN => n9859);
   U7008 : OAI22_X1 port map( A1 => n16991, A2 => n15955, B1 => n16989, B2 => 
                           n16859, ZN => n9867);
   U7009 : OAI22_X1 port map( A1 => n17567, A2 => n16176, B1 => n17562, B2 => 
                           n16803, ZN => n9192);
   U7010 : OAI22_X1 port map( A1 => n17594, A2 => n16050, B1 => n17589, B2 => 
                           n16803, ZN => n9194);
   U7011 : OAI22_X1 port map( A1 => n17608, A2 => n16088, B1 => n17603, B2 => 
                           n16803, ZN => n9195);
   U7012 : OAI22_X1 port map( A1 => n17566, A2 => n16177, B1 => n17562, B2 => 
                           n16809, ZN => n9264);
   U7013 : OAI22_X1 port map( A1 => n17593, A2 => n16051, B1 => n17589, B2 => 
                           n16809, ZN => n9266);
   U7014 : OAI22_X1 port map( A1 => n17607, A2 => n16089, B1 => n17603, B2 => 
                           n16809, ZN => n9267);
   U7015 : OAI22_X1 port map( A1 => n17566, A2 => n16178, B1 => n17562, B2 => 
                           n16815, ZN => n9336);
   U7016 : OAI22_X1 port map( A1 => n17593, A2 => n16052, B1 => n17589, B2 => 
                           n16815, ZN => n9338);
   U7017 : OAI22_X1 port map( A1 => n17607, A2 => n16090, B1 => n17603, B2 => 
                           n16815, ZN => n9339);
   U7018 : OAI22_X1 port map( A1 => n17566, A2 => n16179, B1 => n17562, B2 => 
                           n16827, ZN => n9480);
   U7019 : OAI22_X1 port map( A1 => n17593, A2 => n16053, B1 => n17589, B2 => 
                           n16827, ZN => n9482);
   U7020 : OAI22_X1 port map( A1 => n17607, A2 => n16091, B1 => n17603, B2 => 
                           n16827, ZN => n9483);
   U7021 : OAI22_X1 port map( A1 => n17565, A2 => n16180, B1 => n17562, B2 => 
                           n16833, ZN => n9552);
   U7022 : OAI22_X1 port map( A1 => n17592, A2 => n16054, B1 => n17589, B2 => 
                           n16833, ZN => n9554);
   U7023 : OAI22_X1 port map( A1 => n17606, A2 => n16092, B1 => n17603, B2 => 
                           n16833, ZN => n9555);
   U7024 : OAI22_X1 port map( A1 => n17566, A2 => n16181, B1 => n17562, B2 => 
                           n16839, ZN => n9624);
   U7025 : OAI22_X1 port map( A1 => n17593, A2 => n16055, B1 => n17589, B2 => 
                           n16839, ZN => n9626);
   U7026 : OAI22_X1 port map( A1 => n17607, A2 => n16093, B1 => n17603, B2 => 
                           n16839, ZN => n9627);
   U7027 : OAI22_X1 port map( A1 => n17565, A2 => n16182, B1 => n17562, B2 => 
                           n16845, ZN => n9696);
   U7028 : OAI22_X1 port map( A1 => n17592, A2 => n16056, B1 => n17589, B2 => 
                           n16845, ZN => n9698);
   U7029 : OAI22_X1 port map( A1 => n17606, A2 => n16094, B1 => n17603, B2 => 
                           n16845, ZN => n9699);
   U7030 : OAI22_X1 port map( A1 => n17565, A2 => n16183, B1 => n17562, B2 => 
                           n16851, ZN => n9768);
   U7031 : OAI22_X1 port map( A1 => n17592, A2 => n16057, B1 => n17589, B2 => 
                           n16851, ZN => n9770);
   U7032 : OAI22_X1 port map( A1 => n17606, A2 => n16095, B1 => n17603, B2 => 
                           n16851, ZN => n9771);
   U7033 : OAI22_X1 port map( A1 => n17565, A2 => n16184, B1 => n17562, B2 => 
                           n16857, ZN => n9840);
   U7034 : OAI22_X1 port map( A1 => n17592, A2 => n16058, B1 => n17589, B2 => 
                           n16857, ZN => n9842);
   U7035 : OAI22_X1 port map( A1 => n17606, A2 => n16096, B1 => n17603, B2 => 
                           n16857, ZN => n9843);
   U7036 : OAI22_X1 port map( A1 => n17564, A2 => n16185, B1 => n17562, B2 => 
                           n17512, ZN => n9912);
   U7037 : OAI22_X1 port map( A1 => n17591, A2 => n16059, B1 => n17589, B2 => 
                           n17512, ZN => n9914);
   U7038 : OAI22_X1 port map( A1 => n17605, A2 => n16097, B1 => n17603, B2 => 
                           n17512, ZN => n9915);
   U7039 : OAI22_X1 port map( A1 => n17994, A2 => n16004, B1 => n17989, B2 => 
                           n16810, ZN => n9277);
   U7040 : OAI22_X1 port map( A1 => n17994, A2 => n16005, B1 => n17989, B2 => 
                           n16816, ZN => n9349);
   U7041 : OAI22_X1 port map( A1 => n17993, A2 => n16006, B1 => n17989, B2 => 
                           n16828, ZN => n9493);
   U7042 : OAI22_X1 port map( A1 => n17993, A2 => n16007, B1 => n17989, B2 => 
                           n16834, ZN => n9565);
   U7043 : OAI22_X1 port map( A1 => n17993, A2 => n16008, B1 => n17989, B2 => 
                           n16840, ZN => n9637);
   U7044 : OAI22_X1 port map( A1 => n17992, A2 => n16009, B1 => n17989, B2 => 
                           n16846, ZN => n9709);
   U7045 : OAI22_X1 port map( A1 => n17992, A2 => n16010, B1 => n17989, B2 => 
                           n16852, ZN => n9781);
   U7046 : OAI22_X1 port map( A1 => n17992, A2 => n16011, B1 => n17989, B2 => 
                           n16858, ZN => n9853);
   U7047 : OAI22_X1 port map( A1 => n17993, A2 => n16012, B1 => n17989, B2 => 
                           n17513, ZN => n9925_port);
   U7048 : OAI22_X1 port map( A1 => n17528, A2 => n15858, B1 => n17522, B2 => 
                           n16736, ZN => n8397);
   U7049 : OAI22_X1 port map( A1 => n17528, A2 => n15859, B1 => n17522, B2 => 
                           n16742, ZN => n8469);
   U7050 : OAI22_X1 port map( A1 => n17528, A2 => n15860, B1 => n17522, B2 => 
                           n16748, ZN => n8541);
   U7051 : OAI22_X1 port map( A1 => n17528, A2 => n15861, B1 => n17522, B2 => 
                           n16754, ZN => n8613);
   U7052 : OAI22_X1 port map( A1 => n17527, A2 => n15862, B1 => n17522, B2 => 
                           n16760, ZN => n8685);
   U7053 : OAI22_X1 port map( A1 => n17527, A2 => n15863, B1 => n17522, B2 => 
                           n16766, ZN => n8757);
   U7054 : OAI22_X1 port map( A1 => n17527, A2 => n15864, B1 => n17522, B2 => 
                           n16772, ZN => n8829);
   U7055 : OAI22_X1 port map( A1 => n17526, A2 => n15865, B1 => n17522, B2 => 
                           n16778, ZN => n8901);
   U7056 : OAI22_X1 port map( A1 => n17526, A2 => n15866, B1 => n17522, B2 => 
                           n16784, ZN => n8973);
   U7057 : OAI22_X1 port map( A1 => n17526, A2 => n15867, B1 => n17522, B2 => 
                           n16790, ZN => n9045);
   U7058 : OAI22_X1 port map( A1 => n17526, A2 => n15868, B1 => n17522, B2 => 
                           n16796, ZN => n9117);
   U7059 : OAI22_X1 port map( A1 => n17525, A2 => n15869, B1 => n17521, B2 => 
                           n16802, ZN => n9189);
   U7060 : OAI22_X1 port map( A1 => n17525, A2 => n15870, B1 => n17521, B2 => 
                           n16808, ZN => n9261);
   U7061 : OAI22_X1 port map( A1 => n17525, A2 => n15871, B1 => n17521, B2 => 
                           n16814, ZN => n9333);
   U7062 : OAI22_X1 port map( A1 => n17525, A2 => n15872, B1 => n17521, B2 => 
                           n16820, ZN => n9405);
   U7063 : OAI22_X1 port map( A1 => n17524, A2 => n15873, B1 => n17521, B2 => 
                           n16826, ZN => n9477);
   U7064 : OAI22_X1 port map( A1 => n17524, A2 => n15874, B1 => n17521, B2 => 
                           n16832, ZN => n9549);
   U7065 : OAI22_X1 port map( A1 => n17524, A2 => n15875, B1 => n17521, B2 => 
                           n16838, ZN => n9621);
   U7066 : OAI22_X1 port map( A1 => n17524, A2 => n15876, B1 => n17521, B2 => 
                           n16844, ZN => n9693);
   U7067 : OAI22_X1 port map( A1 => n17523, A2 => n15877, B1 => n17521, B2 => 
                           n16850, ZN => n9765);
   U7068 : OAI22_X1 port map( A1 => n17523, A2 => n15878, B1 => n17521, B2 => 
                           n16856, ZN => n9837);
   U7069 : OAI22_X1 port map( A1 => n17523, A2 => n15879, B1 => n17521, B2 => 
                           n16862, ZN => n9909_port);
   U7070 : OAI22_X1 port map( A1 => n17527, A2 => n15880, B1 => n17521, B2 => 
                           n17517, ZN => n9981);
   U7071 : OAI22_X1 port map( A1 => n17622, A2 => n16138, B1 => n17617, B2 => 
                           n16797, ZN => n9124);
   U7072 : OAI22_X1 port map( A1 => n17622, A2 => n16139, B1 => n17617, B2 => 
                           n16803, ZN => n9196);
   U7073 : OAI22_X1 port map( A1 => n17621, A2 => n16140, B1 => n17617, B2 => 
                           n16809, ZN => n9268);
   U7074 : OAI22_X1 port map( A1 => n17621, A2 => n16141, B1 => n17617, B2 => 
                           n16815, ZN => n9340);
   U7075 : OAI22_X1 port map( A1 => n17621, A2 => n16142, B1 => n17617, B2 => 
                           n16827, ZN => n9484);
   U7076 : OAI22_X1 port map( A1 => n17620, A2 => n16143, B1 => n17617, B2 => 
                           n16833, ZN => n9556);
   U7077 : OAI22_X1 port map( A1 => n17621, A2 => n16144, B1 => n17617, B2 => 
                           n16839, ZN => n9628);
   U7078 : OAI22_X1 port map( A1 => n17620, A2 => n16145, B1 => n17617, B2 => 
                           n16845, ZN => n9700);
   U7079 : OAI22_X1 port map( A1 => n17620, A2 => n16146, B1 => n17617, B2 => 
                           n16851, ZN => n9772);
   U7080 : OAI22_X1 port map( A1 => n17620, A2 => n16147, B1 => n17617, B2 => 
                           n16857, ZN => n9844);
   U7081 : OAI22_X1 port map( A1 => n17619, A2 => n16148, B1 => n17617, B2 => 
                           n17512, ZN => n9916);
   U7082 : OAI22_X1 port map( A1 => n17625, A2 => n16149, B1 => n17618, B2 => 
                           n16731, ZN => n8332);
   U7083 : OAI22_X1 port map( A1 => n17625, A2 => n16150, B1 => n17618, B2 => 
                           n16737, ZN => n8404);
   U7084 : OAI22_X1 port map( A1 => n17997, A2 => n16013, B1 => n17990, B2 => 
                           n16738, ZN => n8413);
   U7085 : OAI22_X1 port map( A1 => n17624, A2 => n16151, B1 => n17618, B2 => 
                           n16743, ZN => n8476);
   U7086 : OAI22_X1 port map( A1 => n17624, A2 => n16152, B1 => n17618, B2 => 
                           n16749, ZN => n8548);
   U7087 : OAI22_X1 port map( A1 => n17997, A2 => n16014, B1 => n17990, B2 => 
                           n16750, ZN => n8557);
   U7088 : OAI22_X1 port map( A1 => n17624, A2 => n16153, B1 => n17618, B2 => 
                           n16755, ZN => n8620);
   U7089 : OAI22_X1 port map( A1 => n17996, A2 => n16015, B1 => n17990, B2 => 
                           n16756, ZN => n8629);
   U7090 : OAI22_X1 port map( A1 => n17624, A2 => n16154, B1 => n17618, B2 => 
                           n16761, ZN => n8692);
   U7091 : OAI22_X1 port map( A1 => n17996, A2 => n16016, B1 => n17990, B2 => 
                           n16762, ZN => n8701);
   U7092 : OAI22_X1 port map( A1 => n17623, A2 => n16155, B1 => n17618, B2 => 
                           n16767, ZN => n8764);
   U7093 : OAI22_X1 port map( A1 => n17996, A2 => n16017, B1 => n17990, B2 => 
                           n16768, ZN => n8773);
   U7094 : OAI22_X1 port map( A1 => n17623, A2 => n16156, B1 => n17618, B2 => 
                           n16773, ZN => n8836);
   U7095 : OAI22_X1 port map( A1 => n17996, A2 => n16018, B1 => n17990, B2 => 
                           n16774, ZN => n8845);
   U7096 : OAI22_X1 port map( A1 => n17623, A2 => n16157, B1 => n17618, B2 => 
                           n16779, ZN => n8908);
   U7097 : OAI22_X1 port map( A1 => n17995, A2 => n16019, B1 => n17990, B2 => 
                           n16780, ZN => n8917);
   U7098 : OAI22_X1 port map( A1 => n17622, A2 => n16158, B1 => n17618, B2 => 
                           n16785, ZN => n8980);
   U7099 : OAI22_X1 port map( A1 => n17995, A2 => n16020, B1 => n17990, B2 => 
                           n16786, ZN => n8989);
   U7100 : OAI22_X1 port map( A1 => n17622, A2 => n16159, B1 => n17618, B2 => 
                           n16791, ZN => n9052);
   U7101 : OAI22_X1 port map( A1 => n17995, A2 => n16021, B1 => n17990, B2 => 
                           n16792, ZN => n9061);
   U7102 : OAI22_X1 port map( A1 => n17994, A2 => n16022, B1 => n17990, B2 => 
                           n16798, ZN => n9133);
   U7103 : OAI22_X1 port map( A1 => n17994, A2 => n16023, B1 => n17990, B2 => 
                           n16804, ZN => n9205);
   U7104 : OAI22_X1 port map( A1 => n17623, A2 => n16160, B1 => n17618, B2 => 
                           n16821, ZN => n9412);
   U7105 : OAI22_X1 port map( A1 => n17995, A2 => n16024, B1 => n17990, B2 => 
                           n16822, ZN => n9421);
   U7106 : OAI22_X1 port map( A1 => n10189, A2 => n14033, B1 => n7588, B2 => 
                           n14034, ZN => n10128);
   U7107 : OAI22_X1 port map( A1 => n7725, A2 => n17833, B1 => n12370, B2 => 
                           n17824, ZN => n7764);
   U7108 : NOR4_X1 port map( A1 => n12371, A2 => n12372, A3 => n12373, A4 => 
                           n12374, ZN => n12370);
   U7109 : NAND4_X1 port map( A1 => n12375, A2 => n12376, A3 => n12377, A4 => 
                           n12378, ZN => n12374);
   U7110 : NAND4_X1 port map( A1 => n12399, A2 => n12400, A3 => n12401, A4 => 
                           n12402, ZN => n12371);
   U7111 : OAI22_X1 port map( A1 => n7724, A2 => n17833, B1 => n12216, B2 => 
                           n17824, ZN => n7839);
   U7112 : NOR4_X1 port map( A1 => n12217, A2 => n12218, A3 => n12219, A4 => 
                           n12220, ZN => n12216);
   U7113 : NAND4_X1 port map( A1 => n12221, A2 => n12222, A3 => n12223, A4 => 
                           n12224, ZN => n12220);
   U7114 : NAND4_X1 port map( A1 => n12245, A2 => n12246, A3 => n12247, A4 => 
                           n12248, ZN => n12217);
   U7115 : OAI22_X1 port map( A1 => n7695, A2 => n17826, B1 => n4091, B2 => 
                           n17824, ZN => n9989);
   U7116 : NOR4_X1 port map( A1 => n4095, A2 => n4098, A3 => n4099, A4 => n4100
                           , ZN => n4091);
   U7117 : NAND4_X1 port map( A1 => n4101, A2 => n4102, A3 => n4103, A4 => 
                           n4106, ZN => n4100);
   U7118 : NAND4_X1 port map( A1 => n4213, A2 => n4214, A3 => n4217, A4 => 
                           n4218, ZN => n4095);
   U7119 : OAI22_X1 port map( A1 => net227471, A2 => n14007, B1 => n14019, B2 
                           => n14009, ZN => n10133);
   U7120 : AOI21_X1 port map( B1 => n14021, B2 => r590_carry_5_port, A => 
                           n14011, ZN => n14019);
   U7121 : OAI22_X1 port map( A1 => net227472, A2 => n14007, B1 => n14018, B2 
                           => n14009, ZN => n10134);
   U7122 : XNOR2_X1 port map( A => n10187, B => n14017, ZN => n14018);
   U7123 : OAI22_X1 port map( A1 => net227473, A2 => n14007, B1 => n14013, B2 
                           => n14009, ZN => n10135);
   U7124 : AOI211_X1 port map( C1 => N9909, C2 => N9908, A => n14016, B => 
                           n14017, ZN => n14013);
   U7125 : OAI22_X1 port map( A1 => net227476, A2 => n14007, B1 => N9641, B2 =>
                           n14009, ZN => n10138);
   U7126 : OAI22_X1 port map( A1 => n7723, A2 => n17833, B1 => n12061, B2 => 
                           n17823, ZN => n7915);
   U7127 : NOR4_X1 port map( A1 => n12062, A2 => n12063, A3 => n12064, A4 => 
                           n12065, ZN => n12061);
   U7128 : NAND4_X1 port map( A1 => n12066, A2 => n12067, A3 => n12068, A4 => 
                           n12069, ZN => n12065);
   U7129 : NAND4_X1 port map( A1 => n12090, A2 => n12091, A3 => n12092, A4 => 
                           n12093, ZN => n12062);
   U7130 : OAI22_X1 port map( A1 => n7722, A2 => n17832, B1 => n11908, B2 => 
                           n17825, ZN => n7989);
   U7131 : NOR4_X1 port map( A1 => n11909, A2 => n11910, A3 => n11911, A4 => 
                           n11912, ZN => n11908);
   U7132 : NAND4_X1 port map( A1 => n11913, A2 => n11914, A3 => n11915, A4 => 
                           n11916, ZN => n11912);
   U7133 : NAND4_X1 port map( A1 => n11937, A2 => n11938, A3 => n11939, A4 => 
                           n11940, ZN => n11909);
   U7134 : OAI22_X1 port map( A1 => n7721, A2 => n17832, B1 => n10465, B2 => 
                           n17823, ZN => n8117);
   U7135 : NOR4_X1 port map( A1 => n10466, A2 => n10467, A3 => n10468, A4 => 
                           n10469, ZN => n10465);
   U7136 : NAND4_X1 port map( A1 => n10470, A2 => n10471, A3 => n10472, A4 => 
                           n10473, ZN => n10469);
   U7137 : NAND4_X1 port map( A1 => n10494, A2 => n10495, A3 => n10496, A4 => 
                           n10497, ZN => n10466);
   U7138 : OAI22_X1 port map( A1 => n7720, A2 => n17832, B1 => n10355, B2 => 
                           n17825, ZN => n8189);
   U7139 : NOR4_X1 port map( A1 => n10356, A2 => n10357, A3 => n10358, A4 => 
                           n10359, ZN => n10355);
   U7140 : NAND4_X1 port map( A1 => n10360, A2 => n10361, A3 => n10362, A4 => 
                           n10363, ZN => n10359);
   U7141 : NAND4_X1 port map( A1 => n10384, A2 => n10385, A3 => n10386, A4 => 
                           n10387, ZN => n10356);
   U7142 : OAI22_X1 port map( A1 => n7719, A2 => n17832, B1 => n10243, B2 => 
                           n17823, ZN => n8261);
   U7143 : NOR4_X1 port map( A1 => n10244, A2 => n10245, A3 => n10246, A4 => 
                           n10247, ZN => n10243);
   U7144 : NAND4_X1 port map( A1 => n10248, A2 => n10249, A3 => n10250, A4 => 
                           n10251, ZN => n10247);
   U7145 : NAND4_X1 port map( A1 => n10272, A2 => n10273, A3 => n10274, A4 => 
                           n10275, ZN => n10244);
   U7146 : OAI22_X1 port map( A1 => n7718, A2 => n17831, B1 => n7607, B2 => 
                           n17825, ZN => n8333);
   U7147 : NOR4_X1 port map( A1 => n7608, A2 => n7609, A3 => n7610, A4 => n7611
                           , ZN => n7607);
   U7148 : NAND4_X1 port map( A1 => n7612, A2 => n7613, A3 => n7614, A4 => 
                           n7615, ZN => n7611);
   U7149 : NAND4_X1 port map( A1 => n7636, A2 => n7637, A3 => n7638, A4 => 
                           n7639, ZN => n7608);
   U7150 : OAI22_X1 port map( A1 => n7717, A2 => n17831, B1 => n7492, B2 => 
                           n17823, ZN => n8405);
   U7151 : NOR4_X1 port map( A1 => n7493, A2 => n7494, A3 => n7495, A4 => n7496
                           , ZN => n7492);
   U7152 : NAND4_X1 port map( A1 => n7497, A2 => n7498, A3 => n7499, A4 => 
                           n7500, ZN => n7496);
   U7153 : NAND4_X1 port map( A1 => n7521, A2 => n7522, A3 => n7523, A4 => 
                           n7524, ZN => n7493);
   U7154 : OAI22_X1 port map( A1 => n7716, A2 => n17831, B1 => n7383, B2 => 
                           n17825, ZN => n8477);
   U7155 : NOR4_X1 port map( A1 => n7384, A2 => n7385, A3 => n7386, A4 => n7387
                           , ZN => n7383);
   U7156 : NAND4_X1 port map( A1 => n7388, A2 => n7389, A3 => n7390, A4 => 
                           n7391, ZN => n7387);
   U7157 : NAND4_X1 port map( A1 => n7412, A2 => n7413, A3 => n7414, A4 => 
                           n7415, ZN => n7384);
   U7158 : OAI22_X1 port map( A1 => n7715, A2 => n17831, B1 => n7274, B2 => 
                           n17823, ZN => n8549);
   U7159 : NOR4_X1 port map( A1 => n7275, A2 => n7276, A3 => n7277, A4 => n7278
                           , ZN => n7274);
   U7160 : NAND4_X1 port map( A1 => n7279, A2 => n7280, A3 => n7281, A4 => 
                           n7282, ZN => n7278);
   U7161 : NAND4_X1 port map( A1 => n7303, A2 => n7304, A3 => n7305, A4 => 
                           n7306, ZN => n7275);
   U7162 : OAI22_X1 port map( A1 => n7714, A2 => n17830, B1 => n7160, B2 => 
                           n17823, ZN => n8621);
   U7163 : NOR4_X1 port map( A1 => n7161, A2 => n7162, A3 => n7163, A4 => n7164
                           , ZN => n7160);
   U7164 : NAND4_X1 port map( A1 => n7165, A2 => n7166, A3 => n7167, A4 => 
                           n7168, ZN => n7164);
   U7165 : NAND4_X1 port map( A1 => n7189, A2 => n7190, A3 => n7191, A4 => 
                           n7192, ZN => n7161);
   U7166 : OAI22_X1 port map( A1 => n7713, A2 => n17830, B1 => n7051, B2 => 
                           n17823, ZN => n8693);
   U7167 : NOR4_X1 port map( A1 => n7052, A2 => n7053, A3 => n7054, A4 => n7055
                           , ZN => n7051);
   U7168 : NAND4_X1 port map( A1 => n7056, A2 => n7057, A3 => n7058, A4 => 
                           n7059, ZN => n7055);
   U7169 : NAND4_X1 port map( A1 => n7080, A2 => n7081, A3 => n7082, A4 => 
                           n7083, ZN => n7052);
   U7170 : OAI22_X1 port map( A1 => n7712, A2 => n17830, B1 => n6942, B2 => 
                           n17825, ZN => n8765);
   U7171 : NOR4_X1 port map( A1 => n6943, A2 => n6944, A3 => n6945, A4 => n6946
                           , ZN => n6942);
   U7172 : NAND4_X1 port map( A1 => n6947, A2 => n6948, A3 => n6949, A4 => 
                           n6950, ZN => n6946);
   U7173 : NAND4_X1 port map( A1 => n6971, A2 => n6972, A3 => n6973, A4 => 
                           n6974, ZN => n6943);
   U7174 : OAI22_X1 port map( A1 => n7711, A2 => n17830, B1 => n6833, B2 => 
                           n17823, ZN => n8837);
   U7175 : NOR4_X1 port map( A1 => n6834, A2 => n6835, A3 => n6836, A4 => n6837
                           , ZN => n6833);
   U7176 : NAND4_X1 port map( A1 => n6838, A2 => n6839, A3 => n6840, A4 => 
                           n6841, ZN => n6837);
   U7177 : NAND4_X1 port map( A1 => n6862, A2 => n6863, A3 => n6864, A4 => 
                           n6865, ZN => n6834);
   U7178 : OAI22_X1 port map( A1 => n7710, A2 => n17829, B1 => n6724, B2 => 
                           n17823, ZN => n8909);
   U7179 : NOR4_X1 port map( A1 => n6725, A2 => n6726, A3 => n6727, A4 => n6728
                           , ZN => n6724);
   U7180 : NAND4_X1 port map( A1 => n6729, A2 => n6730, A3 => n6731, A4 => 
                           n6732, ZN => n6728);
   U7181 : NAND4_X1 port map( A1 => n6753, A2 => n6754, A3 => n6755, A4 => 
                           n6756, ZN => n6725);
   U7182 : OAI22_X1 port map( A1 => n7709, A2 => n17829, B1 => n6560, B2 => 
                           n17825, ZN => n8981);
   U7183 : NOR4_X1 port map( A1 => n6562, A2 => n6563, A3 => n6564, A4 => n6565
                           , ZN => n6560);
   U7184 : NAND4_X1 port map( A1 => n6566, A2 => n6568, A3 => n6570, A4 => 
                           n6572, ZN => n6565);
   U7185 : NAND4_X1 port map( A1 => n6612, A2 => n6614, A3 => n6615, A4 => 
                           n6616, ZN => n6562);
   U7186 : OAI22_X1 port map( A1 => n7708, A2 => n17829, B1 => n6374, B2 => 
                           n17823, ZN => n9053);
   U7187 : NOR4_X1 port map( A1 => n6375, A2 => n6376, A3 => n6377, A4 => n6379
                           , ZN => n6374);
   U7188 : NAND4_X1 port map( A1 => n6381, A2 => n6383, A3 => n6384, A4 => 
                           n6385, ZN => n6379);
   U7189 : NAND4_X1 port map( A1 => n6426, A2 => n6427, A3 => n6428, A4 => 
                           n6429, ZN => n6375);
   U7190 : OAI22_X1 port map( A1 => n7707, A2 => n17829, B1 => n6187, B2 => 
                           n17825, ZN => n9125);
   U7191 : NOR4_X1 port map( A1 => n6188, A2 => n6190, A3 => n6192, A4 => n6194
                           , ZN => n6187);
   U7192 : NAND4_X1 port map( A1 => n6195, A2 => n6196, A3 => n6197, A4 => 
                           n6198, ZN => n6194);
   U7193 : NAND4_X1 port map( A1 => n6239, A2 => n6240, A3 => n6241, A4 => 
                           n6244, ZN => n6188);
   U7194 : OAI22_X1 port map( A1 => n7706, A2 => n17828, B1 => n6001, B2 => 
                           n17825, ZN => n9197);
   U7195 : NOR4_X1 port map( A1 => n6003, A2 => n6005, A3 => n6006, A4 => n6007
                           , ZN => n6001);
   U7196 : NAND4_X1 port map( A1 => n6008, A2 => n6009, A3 => n6010, A4 => 
                           n6013, ZN => n6007);
   U7197 : NAND4_X1 port map( A1 => n6052, A2 => n6055, A3 => n6056, A4 => 
                           n6058, ZN => n6003);
   U7198 : OAI22_X1 port map( A1 => n7705, A2 => n17828, B1 => n5816, B2 => 
                           n17823, ZN => n9269);
   U7199 : NOR4_X1 port map( A1 => n5817, A2 => n5818, A3 => n5819, A4 => n5820
                           , ZN => n5816);
   U7200 : NAND4_X1 port map( A1 => n5821, A2 => n5824, A3 => n5825, A4 => 
                           n5826, ZN => n5820);
   U7201 : NAND4_X1 port map( A1 => n5867, A2 => n5869, A3 => n5870, A4 => 
                           n5871, ZN => n5817);
   U7202 : OAI22_X1 port map( A1 => n7704, A2 => n17828, B1 => n5629, B2 => 
                           n17823, ZN => n9341);
   U7203 : NOR4_X1 port map( A1 => n5630, A2 => n5631, A3 => n5632, A4 => n5635
                           , ZN => n5629);
   U7204 : NAND4_X1 port map( A1 => n5636, A2 => n5637, A3 => n5653, A4 => 
                           n5654, ZN => n5635);
   U7205 : NAND4_X1 port map( A1 => n5681, A2 => n5682, A3 => n5683, A4 => 
                           n5684, ZN => n5630);
   U7206 : OAI22_X1 port map( A1 => n7703, A2 => n17828, B1 => n5442, B2 => 
                           n17823, ZN => n9413);
   U7207 : NOR4_X1 port map( A1 => n5443, A2 => n5446, A3 => n5447, A4 => n5448
                           , ZN => n5442);
   U7208 : NAND4_X1 port map( A1 => n5464, A2 => n5465, A3 => n5466, A4 => 
                           n5467, ZN => n5448);
   U7209 : NAND4_X1 port map( A1 => n5494, A2 => n5495, A3 => n5497, A4 => 
                           n5499, ZN => n5443);
   U7210 : OAI22_X1 port map( A1 => n7702, A2 => n17827, B1 => n5257, B2 => 
                           n17823, ZN => n9485);
   U7211 : NOR4_X1 port map( A1 => n5259, A2 => n5274, A3 => n5275, A4 => n5276
                           , ZN => n5257);
   U7212 : NAND4_X1 port map( A1 => n5277, A2 => n5278, A3 => n5279, A4 => 
                           n5280, ZN => n5276);
   U7213 : NAND4_X1 port map( A1 => n5309, A2 => n5311, A3 => n5312, A4 => 
                           n5313, ZN => n5259);
   U7214 : OAI22_X1 port map( A1 => n7701, A2 => n17827, B1 => n5106, B2 => 
                           n17825, ZN => n9557);
   U7215 : NOR4_X1 port map( A1 => n5107, A2 => n5108, A3 => n5109, A4 => n5110
                           , ZN => n5106);
   U7216 : NAND4_X1 port map( A1 => n5111, A2 => n5112, A3 => n5113, A4 => 
                           n5115, ZN => n5110);
   U7217 : NAND4_X1 port map( A1 => n5138, A2 => n5139, A3 => n5140, A4 => 
                           n5141, ZN => n5107);
   U7218 : OAI22_X1 port map( A1 => n7700, A2 => n17827, B1 => n4993, B2 => 
                           n17825, ZN => n9629);
   U7219 : NOR4_X1 port map( A1 => n4994, A2 => n4995, A3 => n4996, A4 => n4997
                           , ZN => n4993);
   U7220 : NAND4_X1 port map( A1 => n4998, A2 => n4999, A3 => n5000, A4 => 
                           n5001, ZN => n4997);
   U7221 : NAND4_X1 port map( A1 => n5024, A2 => n5025, A3 => n5026, A4 => 
                           n5027, ZN => n4994);
   U7222 : OAI22_X1 port map( A1 => n3043, A2 => n14033, B1 => n7592, B2 => 
                           n14034, ZN => n10132);
   U7223 : OAI22_X1 port map( A1 => n10190, A2 => n14033, B1 => n7587, B2 => 
                           n14034, ZN => n10127);
   U7224 : OAI22_X1 port map( A1 => n10188, A2 => n14033, B1 => n7589, B2 => 
                           n14034, ZN => n10129);
   U7225 : OAI22_X1 port map( A1 => n10187, A2 => n14033, B1 => n7590, B2 => 
                           n14034, ZN => n10130);
   U7226 : OAI22_X1 port map( A1 => n14820, A2 => n14033, B1 => n7591, B2 => 
                           n14034, ZN => n10131);
   U7227 : OAI22_X1 port map( A1 => n17535, A2 => n18027, B1 => n17536, B2 => 
                           n16025, ZN => n9982);
   U7228 : OAI22_X1 port map( A1 => n17549, A2 => n18027, B1 => n17550, B2 => 
                           n16030, ZN => n9983);
   U7229 : OAI22_X1 port map( A1 => n17563, A2 => n18027, B1 => n17564, B2 => 
                           n16032, ZN => n9984);
   U7230 : OAI22_X1 port map( A1 => n17590, A2 => n18027, B1 => n17591, B2 => 
                           n16026, ZN => n9986);
   U7231 : OAI22_X1 port map( A1 => n17604, A2 => n18026, B1 => n17605, B2 => 
                           n16027, ZN => n9987);
   U7232 : OAI22_X1 port map( A1 => n17618, A2 => n18026, B1 => n17619, B2 => 
                           n16031, ZN => n9988);
   U7233 : OAI22_X1 port map( A1 => n17990, A2 => n18026, B1 => n17991, B2 => 
                           n15789, ZN => n9997);
   U7234 : OAI22_X1 port map( A1 => n16901, A2 => n18031, B1 => n15788, B2 => 
                           n16902, ZN => n10003);
   U7235 : OAI22_X1 port map( A1 => n16990, A2 => n18031, B1 => n15787, B2 => 
                           n16991, ZN => n10011);
   U7236 : OAI22_X1 port map( A1 => n17151, A2 => n18029, B1 => n15783, B2 => 
                           n17152, ZN => n10024);
   U7237 : OAI22_X1 port map( A1 => n17217, A2 => n18029, B1 => n15786, B2 => 
                           n17218, ZN => n10030);
   U7238 : OAI22_X1 port map( A1 => n17269, A2 => n18029, B1 => n15784, B2 => 
                           n17270, ZN => n10034);
   U7239 : OAI22_X1 port map( A1 => n17549, A2 => n16701, B1 => n17550, B2 => 
                           n16033, ZN => n10055);
   U7240 : OAI22_X1 port map( A1 => n17563, A2 => n16701, B1 => n17564, B2 => 
                           n16035, ZN => n10056);
   U7241 : OAI22_X1 port map( A1 => n17590, A2 => n16701, B1 => n17591, B2 => 
                           n16029, ZN => n10058);
   U7242 : OAI22_X1 port map( A1 => n17604, A2 => n16701, B1 => n17605, B2 => 
                           n16028, ZN => n10059);
   U7243 : OAI22_X1 port map( A1 => n17618, A2 => n16701, B1 => n17619, B2 => 
                           n16034, ZN => n10060);
   U7244 : OAI22_X1 port map( A1 => n17990, A2 => n16702, B1 => n17991, B2 => 
                           n15790, ZN => n10069);
   U7245 : OAI22_X1 port map( A1 => n17570, A2 => n16186, B1 => n17563, B2 => 
                           n16731, ZN => n8328);
   U7246 : OAI22_X1 port map( A1 => n17597, A2 => n16060, B1 => n17590, B2 => 
                           n16731, ZN => n8330);
   U7247 : OAI22_X1 port map( A1 => n17611, A2 => n16098, B1 => n17604, B2 => 
                           n16731, ZN => n8331);
   U7248 : OAI22_X1 port map( A1 => n17556, A2 => n16161, B1 => n17549, B2 => 
                           n16737, ZN => n8399);
   U7249 : OAI22_X1 port map( A1 => n17570, A2 => n16187, B1 => n17563, B2 => 
                           n16737, ZN => n8400);
   U7250 : OAI22_X1 port map( A1 => n17597, A2 => n16061, B1 => n17590, B2 => 
                           n16737, ZN => n8402);
   U7251 : OAI22_X1 port map( A1 => n17611, A2 => n16099, B1 => n17604, B2 => 
                           n16737, ZN => n8403);
   U7252 : OAI22_X1 port map( A1 => n17541, A2 => n16062, B1 => n17535, B2 => 
                           n16743, ZN => n8470);
   U7253 : OAI22_X1 port map( A1 => n17555, A2 => n16162, B1 => n17549, B2 => 
                           n16743, ZN => n8471);
   U7254 : OAI22_X1 port map( A1 => n17569, A2 => n16188, B1 => n17563, B2 => 
                           n16743, ZN => n8472);
   U7255 : OAI22_X1 port map( A1 => n17596, A2 => n16063, B1 => n17590, B2 => 
                           n16743, ZN => n8474);
   U7256 : OAI22_X1 port map( A1 => n17610, A2 => n16100, B1 => n17604, B2 => 
                           n16743, ZN => n8475);
   U7257 : OAI22_X1 port map( A1 => n17541, A2 => n16064, B1 => n17535, B2 => 
                           n16749, ZN => n8542);
   U7258 : OAI22_X1 port map( A1 => n17555, A2 => n16163, B1 => n17549, B2 => 
                           n16749, ZN => n8543);
   U7259 : OAI22_X1 port map( A1 => n17569, A2 => n16189, B1 => n17563, B2 => 
                           n16749, ZN => n8544);
   U7260 : OAI22_X1 port map( A1 => n17596, A2 => n16065, B1 => n17590, B2 => 
                           n16749, ZN => n8546);
   U7261 : OAI22_X1 port map( A1 => n17610, A2 => n16101, B1 => n17604, B2 => 
                           n16749, ZN => n8547);
   U7262 : OAI22_X1 port map( A1 => n16873, A2 => n15956, B1 => n16867, B2 => 
                           n16750, ZN => n8560);
   U7263 : OAI22_X1 port map( A1 => n17541, A2 => n16066, B1 => n17535, B2 => 
                           n16755, ZN => n8614);
   U7264 : OAI22_X1 port map( A1 => n17555, A2 => n16164, B1 => n17549, B2 => 
                           n16755, ZN => n8615);
   U7265 : OAI22_X1 port map( A1 => n17569, A2 => n16190, B1 => n17563, B2 => 
                           n16755, ZN => n8616);
   U7266 : OAI22_X1 port map( A1 => n17596, A2 => n16067, B1 => n17590, B2 => 
                           n16755, ZN => n8618);
   U7267 : OAI22_X1 port map( A1 => n17610, A2 => n16102, B1 => n17604, B2 => 
                           n16755, ZN => n8619);
   U7268 : OAI22_X1 port map( A1 => n16873, A2 => n15957, B1 => n16867, B2 => 
                           n16756, ZN => n8632);
   U7269 : OAI22_X1 port map( A1 => n17540, A2 => n16068, B1 => n17535, B2 => 
                           n16761, ZN => n8686);
   U7270 : OAI22_X1 port map( A1 => n17555, A2 => n16165, B1 => n17549, B2 => 
                           n16761, ZN => n8687);
   U7271 : OAI22_X1 port map( A1 => n17569, A2 => n16191, B1 => n17563, B2 => 
                           n16761, ZN => n8688);
   U7272 : OAI22_X1 port map( A1 => n17596, A2 => n16069, B1 => n17590, B2 => 
                           n16761, ZN => n8690);
   U7273 : OAI22_X1 port map( A1 => n17610, A2 => n16103, B1 => n17604, B2 => 
                           n16761, ZN => n8691);
   U7274 : OAI22_X1 port map( A1 => n16873, A2 => n15958, B1 => n16867, B2 => 
                           n16762, ZN => n8704);
   U7275 : OAI22_X1 port map( A1 => n17540, A2 => n16070, B1 => n17535, B2 => 
                           n16767, ZN => n8758);
   U7276 : OAI22_X1 port map( A1 => n17554, A2 => n16166, B1 => n17549, B2 => 
                           n16767, ZN => n8759);
   U7277 : OAI22_X1 port map( A1 => n17568, A2 => n16192, B1 => n17563, B2 => 
                           n16767, ZN => n8760);
   U7278 : OAI22_X1 port map( A1 => n17595, A2 => n16071, B1 => n17590, B2 => 
                           n16767, ZN => n8762);
   U7279 : OAI22_X1 port map( A1 => n17609, A2 => n16104, B1 => n17604, B2 => 
                           n16767, ZN => n8763);
   U7280 : OAI22_X1 port map( A1 => n16872, A2 => n15959, B1 => n16867, B2 => 
                           n16768, ZN => n8776);
   U7281 : OAI22_X1 port map( A1 => n17540, A2 => n16072, B1 => n17535, B2 => 
                           n16773, ZN => n8830);
   U7282 : OAI22_X1 port map( A1 => n17554, A2 => n16167, B1 => n17549, B2 => 
                           n16773, ZN => n8831);
   U7283 : OAI22_X1 port map( A1 => n17568, A2 => n16193, B1 => n17563, B2 => 
                           n16773, ZN => n8832);
   U7284 : OAI22_X1 port map( A1 => n17595, A2 => n16073, B1 => n17590, B2 => 
                           n16773, ZN => n8834);
   U7285 : OAI22_X1 port map( A1 => n17609, A2 => n16105, B1 => n17604, B2 => 
                           n16773, ZN => n8835);
   U7286 : OAI22_X1 port map( A1 => n16872, A2 => n15960, B1 => n16867, B2 => 
                           n16774, ZN => n8848);
   U7287 : OAI22_X1 port map( A1 => n17539, A2 => n16074, B1 => n17535, B2 => 
                           n16779, ZN => n8902);
   U7288 : OAI22_X1 port map( A1 => n17554, A2 => n16168, B1 => n17549, B2 => 
                           n16779, ZN => n8903);
   U7289 : OAI22_X1 port map( A1 => n17568, A2 => n16194, B1 => n17563, B2 => 
                           n16779, ZN => n8904);
   U7290 : OAI22_X1 port map( A1 => n17595, A2 => n16075, B1 => n17590, B2 => 
                           n16779, ZN => n8906);
   U7291 : OAI22_X1 port map( A1 => n17609, A2 => n16106, B1 => n17604, B2 => 
                           n16779, ZN => n8907);
   U7292 : OAI22_X1 port map( A1 => n16872, A2 => n15961, B1 => n16867, B2 => 
                           n16780, ZN => n8920);
   U7293 : OAI22_X1 port map( A1 => n17539, A2 => n16076, B1 => n17535, B2 => 
                           n16785, ZN => n8974);
   U7294 : OAI22_X1 port map( A1 => n17553, A2 => n16169, B1 => n17549, B2 => 
                           n16785, ZN => n8975);
   U7295 : OAI22_X1 port map( A1 => n17567, A2 => n16195, B1 => n17563, B2 => 
                           n16785, ZN => n8976);
   U7296 : OAI22_X1 port map( A1 => n17594, A2 => n16077, B1 => n17590, B2 => 
                           n16785, ZN => n8978);
   U7297 : OAI22_X1 port map( A1 => n17608, A2 => n16107, B1 => n17604, B2 => 
                           n16785, ZN => n8979);
   U7298 : OAI22_X1 port map( A1 => n16871, A2 => n15962, B1 => n16867, B2 => 
                           n16786, ZN => n8992);
   U7299 : OAI22_X1 port map( A1 => n17539, A2 => n16078, B1 => n17535, B2 => 
                           n16791, ZN => n9046);
   U7300 : OAI22_X1 port map( A1 => n17553, A2 => n16170, B1 => n17549, B2 => 
                           n16791, ZN => n9047);
   U7301 : OAI22_X1 port map( A1 => n17567, A2 => n16196, B1 => n17563, B2 => 
                           n16791, ZN => n9048);
   U7302 : OAI22_X1 port map( A1 => n17594, A2 => n16079, B1 => n17590, B2 => 
                           n16791, ZN => n9050);
   U7303 : OAI22_X1 port map( A1 => n17608, A2 => n16108, B1 => n17604, B2 => 
                           n16791, ZN => n9051);
   U7304 : OAI22_X1 port map( A1 => n16871, A2 => n15963, B1 => n16867, B2 => 
                           n16792, ZN => n9064);
   U7305 : OAI22_X1 port map( A1 => n17539, A2 => n16080, B1 => n17535, B2 => 
                           n16797, ZN => n9118);
   U7306 : OAI22_X1 port map( A1 => n17553, A2 => n16171, B1 => n17549, B2 => 
                           n16797, ZN => n9119);
   U7307 : OAI22_X1 port map( A1 => n17567, A2 => n16197, B1 => n17563, B2 => 
                           n16797, ZN => n9120);
   U7308 : OAI22_X1 port map( A1 => n17594, A2 => n16081, B1 => n17590, B2 => 
                           n16797, ZN => n9122);
   U7309 : OAI22_X1 port map( A1 => n17608, A2 => n16109, B1 => n17604, B2 => 
                           n16797, ZN => n9123);
   U7310 : OAI22_X1 port map( A1 => n16871, A2 => n15964, B1 => n16867, B2 => 
                           n16798, ZN => n9136);
   U7311 : OAI22_X1 port map( A1 => n17553, A2 => n16172, B1 => n17549, B2 => 
                           n16803, ZN => n9191);
   U7312 : OAI22_X1 port map( A1 => n16871, A2 => n15965, B1 => n16867, B2 => 
                           n16804, ZN => n9208);
   U7313 : OAI22_X1 port map( A1 => n17538, A2 => n16082, B1 => n17535, B2 => 
                           n16809, ZN => n9262);
   U7314 : OAI22_X1 port map( A1 => n16870, A2 => n15966, B1 => n16867, B2 => 
                           n16810, ZN => n9280);
   U7315 : OAI22_X1 port map( A1 => n16870, A2 => n15967, B1 => n16867, B2 => 
                           n16816, ZN => n9352);
   U7316 : OAI22_X1 port map( A1 => n17540, A2 => n16083, B1 => n17535, B2 => 
                           n16821, ZN => n9406);
   U7317 : OAI22_X1 port map( A1 => n17554, A2 => n16173, B1 => n17549, B2 => 
                           n16821, ZN => n9407);
   U7318 : OAI22_X1 port map( A1 => n17568, A2 => n16198, B1 => n17563, B2 => 
                           n16821, ZN => n9408);
   U7319 : OAI22_X1 port map( A1 => n17595, A2 => n16084, B1 => n17590, B2 => 
                           n16821, ZN => n9410);
   U7320 : OAI22_X1 port map( A1 => n17609, A2 => n16110, B1 => n17604, B2 => 
                           n16821, ZN => n9411);
   U7321 : OAI22_X1 port map( A1 => n16872, A2 => n15968, B1 => n16867, B2 => 
                           n17513, ZN => n9928);
   U7322 : OAI22_X1 port map( A1 => n17521, A2 => n18027, B1 => n15785, B2 => 
                           n17523, ZN => n10053);
   U7323 : OAI22_X1 port map( A1 => n17538, A2 => n16085, B1 => n17535, B2 => 
                           n16803, ZN => n9190);
   U7324 : NAND2_X1 port map( A1 => add_rd1(3), A2 => add_rd1(4), ZN => n12502)
                           ;
   U7325 : NOR2_X1 port map( A1 => n14265, A2 => n7592, ZN => n14231);
   U7326 : NAND4_X1 port map( A1 => n12509, A2 => n12510, A3 => n12511, A4 => 
                           n12512, ZN => n12492);
   U7327 : XNOR2_X1 port map( A => add_rd1(0), B => add_wr(0), ZN => n12510);
   U7328 : XNOR2_X1 port map( A => add_rd1(1), B => add_wr(1), ZN => n12511);
   U7329 : XNOR2_X1 port map( A => add_rd1(4), B => add_wr(4), ZN => n12509);
   U7330 : INV_X1 port map( A => n14023, ZN => n14025);
   U7331 : NAND2_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), ZN => n13983)
                           ;
   U7332 : NAND4_X1 port map( A1 => n13990, A2 => n13991, A3 => n13992, A4 => 
                           n13993, ZN => n13973);
   U7333 : XNOR2_X1 port map( A => add_rd2(4), B => add_wr(4), ZN => n13990);
   U7334 : XNOR2_X1 port map( A => add_rd2(0), B => add_wr(0), ZN => n13991);
   U7335 : XNOR2_X1 port map( A => add_rd2(1), B => add_wr(1), ZN => n13992);
   U7336 : NAND2_X1 port map( A1 => n14223, A2 => n14224, ZN => n14214);
   U7337 : INV_X1 port map( A => add_wr(2), ZN => n14224);
   U7338 : NAND2_X1 port map( A1 => n5522, A2 => n14821, ZN => n14006);
   U7339 : AOI21_X1 port map( B1 => n16414, B2 => net226799, A => n13907, ZN =>
                           n13906);
   U7340 : NOR4_X1 port map( A1 => n13908, A2 => n13909, A3 => n13910, A4 => 
                           n13911, ZN => n13907);
   U7341 : NAND4_X1 port map( A1 => n13964, A2 => n13965, A3 => n13966, A4 => 
                           n13967, ZN => n13908);
   U7342 : NAND4_X1 port map( A1 => n13948, A2 => n13949, A3 => n13950, A4 => 
                           n13951, ZN => n13909);
   U7343 : AOI21_X1 port map( B1 => n16417, B2 => net226800, A => n13860, ZN =>
                           n13859);
   U7344 : NOR4_X1 port map( A1 => n13861, A2 => n13862, A3 => n13863, A4 => 
                           n13864, ZN => n13860);
   U7345 : NAND4_X1 port map( A1 => n13889, A2 => n13890, A3 => n13891, A4 => 
                           n13892, ZN => n13861);
   U7346 : NAND4_X1 port map( A1 => n13881, A2 => n13882, A3 => n13883, A4 => 
                           n13884, ZN => n13862);
   U7347 : AOI21_X1 port map( B1 => n16417, B2 => net226801, A => n13818, ZN =>
                           n13817);
   U7348 : NOR4_X1 port map( A1 => n13819, A2 => n13820, A3 => n13821, A4 => 
                           n13822, ZN => n13818);
   U7349 : NAND4_X1 port map( A1 => n13847, A2 => n13848, A3 => n13849, A4 => 
                           n13850, ZN => n13819);
   U7350 : NAND4_X1 port map( A1 => n13839, A2 => n13840, A3 => n13841, A4 => 
                           n13842, ZN => n13820);
   U7351 : AOI21_X1 port map( B1 => n16417, B2 => net226802, A => n13776, ZN =>
                           n13775);
   U7352 : NOR4_X1 port map( A1 => n13777, A2 => n13778, A3 => n13779, A4 => 
                           n13780, ZN => n13776);
   U7353 : NAND4_X1 port map( A1 => n13805, A2 => n13806, A3 => n13807, A4 => 
                           n13808, ZN => n13777);
   U7354 : NAND4_X1 port map( A1 => n13797, A2 => n13798, A3 => n13799, A4 => 
                           n13800, ZN => n13778);
   U7355 : AOI21_X1 port map( B1 => n16416, B2 => net226803, A => n13734, ZN =>
                           n13733);
   U7356 : NOR4_X1 port map( A1 => n13735, A2 => n13736, A3 => n13737, A4 => 
                           n13738, ZN => n13734);
   U7357 : NAND4_X1 port map( A1 => n13763, A2 => n13764, A3 => n13765, A4 => 
                           n13766, ZN => n13735);
   U7358 : NAND4_X1 port map( A1 => n13755, A2 => n13756, A3 => n13757, A4 => 
                           n13758, ZN => n13736);
   U7359 : AOI21_X1 port map( B1 => n16416, B2 => net226804, A => n13692, ZN =>
                           n13691);
   U7360 : NOR4_X1 port map( A1 => n13693, A2 => n13694, A3 => n13695, A4 => 
                           n13696, ZN => n13692);
   U7361 : NAND4_X1 port map( A1 => n13721, A2 => n13722, A3 => n13723, A4 => 
                           n13724, ZN => n13693);
   U7362 : NAND4_X1 port map( A1 => n13713, A2 => n13714, A3 => n13715, A4 => 
                           n13716, ZN => n13694);
   U7363 : AOI21_X1 port map( B1 => n16416, B2 => net226805, A => n13650, ZN =>
                           n13649);
   U7364 : NOR4_X1 port map( A1 => n13651, A2 => n13652, A3 => n13653, A4 => 
                           n13654, ZN => n13650);
   U7365 : NAND4_X1 port map( A1 => n13679, A2 => n13680, A3 => n13681, A4 => 
                           n13682, ZN => n13651);
   U7366 : NAND4_X1 port map( A1 => n13671, A2 => n13672, A3 => n13673, A4 => 
                           n13674, ZN => n13652);
   U7367 : AOI21_X1 port map( B1 => n16416, B2 => net226806, A => n13608, ZN =>
                           n13607);
   U7368 : NOR4_X1 port map( A1 => n13609, A2 => n13610, A3 => n13611, A4 => 
                           n13612, ZN => n13608);
   U7369 : NAND4_X1 port map( A1 => n13637, A2 => n13638, A3 => n13639, A4 => 
                           n13640, ZN => n13609);
   U7370 : NAND4_X1 port map( A1 => n13629, A2 => n13630, A3 => n13631, A4 => 
                           n13632, ZN => n13610);
   U7371 : AOI21_X1 port map( B1 => n16416, B2 => net226807, A => n13566, ZN =>
                           n13565);
   U7372 : NOR4_X1 port map( A1 => n13567, A2 => n13568, A3 => n13569, A4 => 
                           n13570, ZN => n13566);
   U7373 : NAND4_X1 port map( A1 => n13595, A2 => n13596, A3 => n13597, A4 => 
                           n13598, ZN => n13567);
   U7374 : NAND4_X1 port map( A1 => n13587, A2 => n13588, A3 => n13589, A4 => 
                           n13590, ZN => n13568);
   U7375 : AOI21_X1 port map( B1 => n16416, B2 => net226808, A => n13524, ZN =>
                           n13523);
   U7376 : NOR4_X1 port map( A1 => n13525, A2 => n13526, A3 => n13527, A4 => 
                           n13528, ZN => n13524);
   U7377 : NAND4_X1 port map( A1 => n13553, A2 => n13554, A3 => n13555, A4 => 
                           n13556, ZN => n13525);
   U7378 : NAND4_X1 port map( A1 => n13545, A2 => n13546, A3 => n13547, A4 => 
                           n13548, ZN => n13526);
   U7379 : AOI21_X1 port map( B1 => n16416, B2 => net226809, A => n13482, ZN =>
                           n13481);
   U7380 : NOR4_X1 port map( A1 => n13483, A2 => n13484, A3 => n13485, A4 => 
                           n13486, ZN => n13482);
   U7381 : NAND4_X1 port map( A1 => n13511, A2 => n13512, A3 => n13513, A4 => 
                           n13514, ZN => n13483);
   U7382 : NAND4_X1 port map( A1 => n13503, A2 => n13504, A3 => n13505, A4 => 
                           n13506, ZN => n13484);
   U7383 : AOI21_X1 port map( B1 => n16416, B2 => net226810, A => n13440, ZN =>
                           n13439);
   U7384 : NOR4_X1 port map( A1 => n13441, A2 => n13442, A3 => n13443, A4 => 
                           n13444, ZN => n13440);
   U7385 : NAND4_X1 port map( A1 => n13469, A2 => n13470, A3 => n13471, A4 => 
                           n13472, ZN => n13441);
   U7386 : NAND4_X1 port map( A1 => n13461, A2 => n13462, A3 => n13463, A4 => 
                           n13464, ZN => n13442);
   U7387 : AOI21_X1 port map( B1 => n16416, B2 => net226811, A => n13398, ZN =>
                           n13397);
   U7388 : NOR4_X1 port map( A1 => n13399, A2 => n13400, A3 => n13401, A4 => 
                           n13402, ZN => n13398);
   U7389 : NAND4_X1 port map( A1 => n13427, A2 => n13428, A3 => n13429, A4 => 
                           n13430, ZN => n13399);
   U7390 : NAND4_X1 port map( A1 => n13419, A2 => n13420, A3 => n13421, A4 => 
                           n13422, ZN => n13400);
   U7391 : AOI21_X1 port map( B1 => n16416, B2 => net226812, A => n13356, ZN =>
                           n13355);
   U7392 : NOR4_X1 port map( A1 => n13357, A2 => n13358, A3 => n13359, A4 => 
                           n13360, ZN => n13356);
   U7393 : NAND4_X1 port map( A1 => n13385, A2 => n13386, A3 => n13387, A4 => 
                           n13388, ZN => n13357);
   U7394 : NAND4_X1 port map( A1 => n13377, A2 => n13378, A3 => n13379, A4 => 
                           n13380, ZN => n13358);
   U7395 : AOI21_X1 port map( B1 => n16416, B2 => net226813, A => n13314, ZN =>
                           n13313);
   U7396 : NOR4_X1 port map( A1 => n13315, A2 => n13316, A3 => n13317, A4 => 
                           n13318, ZN => n13314);
   U7397 : NAND4_X1 port map( A1 => n13343, A2 => n13344, A3 => n13345, A4 => 
                           n13346, ZN => n13315);
   U7398 : NAND4_X1 port map( A1 => n13335, A2 => n13336, A3 => n13337, A4 => 
                           n13338, ZN => n13316);
   U7399 : AOI21_X1 port map( B1 => n16416, B2 => net226814, A => n13272, ZN =>
                           n13271);
   U7400 : NOR4_X1 port map( A1 => n13273, A2 => n13274, A3 => n13275, A4 => 
                           n13276, ZN => n13272);
   U7401 : NAND4_X1 port map( A1 => n13301, A2 => n13302, A3 => n13303, A4 => 
                           n13304, ZN => n13273);
   U7402 : NAND4_X1 port map( A1 => n13293, A2 => n13294, A3 => n13295, A4 => 
                           n13296, ZN => n13274);
   U7403 : AOI21_X1 port map( B1 => n16416, B2 => net226815, A => n13230, ZN =>
                           n13229);
   U7404 : NOR4_X1 port map( A1 => n13231, A2 => n13232, A3 => n13233, A4 => 
                           n13234, ZN => n13230);
   U7405 : NAND4_X1 port map( A1 => n13259, A2 => n13260, A3 => n13261, A4 => 
                           n13262, ZN => n13231);
   U7406 : NAND4_X1 port map( A1 => n13251, A2 => n13252, A3 => n13253, A4 => 
                           n13254, ZN => n13232);
   U7407 : AOI21_X1 port map( B1 => n16415, B2 => net226816, A => n13188, ZN =>
                           n13187);
   U7408 : NOR4_X1 port map( A1 => n13189, A2 => n13190, A3 => n13191, A4 => 
                           n13192, ZN => n13188);
   U7409 : NAND4_X1 port map( A1 => n13217, A2 => n13218, A3 => n13219, A4 => 
                           n13220, ZN => n13189);
   U7410 : NAND4_X1 port map( A1 => n13209, A2 => n13210, A3 => n13211, A4 => 
                           n13212, ZN => n13190);
   U7411 : AOI21_X1 port map( B1 => n16415, B2 => net226817, A => n13146, ZN =>
                           n13145);
   U7412 : NOR4_X1 port map( A1 => n13147, A2 => n13148, A3 => n13149, A4 => 
                           n13150, ZN => n13146);
   U7413 : NAND4_X1 port map( A1 => n13175, A2 => n13176, A3 => n13177, A4 => 
                           n13178, ZN => n13147);
   U7414 : NAND4_X1 port map( A1 => n13167, A2 => n13168, A3 => n13169, A4 => 
                           n13170, ZN => n13148);
   U7415 : AOI21_X1 port map( B1 => n16415, B2 => net226818, A => n13104, ZN =>
                           n13103);
   U7416 : NOR4_X1 port map( A1 => n13105, A2 => n13106, A3 => n13107, A4 => 
                           n13108, ZN => n13104);
   U7417 : NAND4_X1 port map( A1 => n13133, A2 => n13134, A3 => n13135, A4 => 
                           n13136, ZN => n13105);
   U7418 : NAND4_X1 port map( A1 => n13125, A2 => n13126, A3 => n13127, A4 => 
                           n13128, ZN => n13106);
   U7419 : AOI21_X1 port map( B1 => n16415, B2 => net226819, A => n13062, ZN =>
                           n13061);
   U7420 : NOR4_X1 port map( A1 => n13063, A2 => n13064, A3 => n13065, A4 => 
                           n13066, ZN => n13062);
   U7421 : NAND4_X1 port map( A1 => n13091, A2 => n13092, A3 => n13093, A4 => 
                           n13094, ZN => n13063);
   U7422 : NAND4_X1 port map( A1 => n13083, A2 => n13084, A3 => n13085, A4 => 
                           n13086, ZN => n13064);
   U7423 : AOI21_X1 port map( B1 => n16415, B2 => net226820, A => n13020, ZN =>
                           n13019);
   U7424 : NOR4_X1 port map( A1 => n13021, A2 => n13022, A3 => n13023, A4 => 
                           n13024, ZN => n13020);
   U7425 : NAND4_X1 port map( A1 => n13049, A2 => n13050, A3 => n13051, A4 => 
                           n13052, ZN => n13021);
   U7426 : NAND4_X1 port map( A1 => n13041, A2 => n13042, A3 => n13043, A4 => 
                           n13044, ZN => n13022);
   U7427 : AOI21_X1 port map( B1 => n16415, B2 => net226821, A => n12978, ZN =>
                           n12977);
   U7428 : NOR4_X1 port map( A1 => n12979, A2 => n12980, A3 => n12981, A4 => 
                           n12982, ZN => n12978);
   U7429 : NAND4_X1 port map( A1 => n13007, A2 => n13008, A3 => n13009, A4 => 
                           n13010, ZN => n12979);
   U7430 : NAND4_X1 port map( A1 => n12999, A2 => n13000, A3 => n13001, A4 => 
                           n13002, ZN => n12980);
   U7431 : AOI21_X1 port map( B1 => n16415, B2 => net226822, A => n12936, ZN =>
                           n12935);
   U7432 : NOR4_X1 port map( A1 => n12937, A2 => n12938, A3 => n12939, A4 => 
                           n12940, ZN => n12936);
   U7433 : NAND4_X1 port map( A1 => n12965, A2 => n12966, A3 => n12967, A4 => 
                           n12968, ZN => n12937);
   U7434 : NAND4_X1 port map( A1 => n12957, A2 => n12958, A3 => n12959, A4 => 
                           n12960, ZN => n12938);
   U7435 : AOI21_X1 port map( B1 => n16415, B2 => net226823, A => n12894, ZN =>
                           n12893);
   U7436 : NOR4_X1 port map( A1 => n12895, A2 => n12896, A3 => n12897, A4 => 
                           n12898, ZN => n12894);
   U7437 : NAND4_X1 port map( A1 => n12923, A2 => n12924, A3 => n12925, A4 => 
                           n12926, ZN => n12895);
   U7438 : NAND4_X1 port map( A1 => n12915, A2 => n12916, A3 => n12917, A4 => 
                           n12918, ZN => n12896);
   U7439 : AOI21_X1 port map( B1 => n16415, B2 => net226824, A => n12852, ZN =>
                           n12851);
   U7440 : NOR4_X1 port map( A1 => n12853, A2 => n12854, A3 => n12855, A4 => 
                           n12856, ZN => n12852);
   U7441 : NAND4_X1 port map( A1 => n12881, A2 => n12882, A3 => n12883, A4 => 
                           n12884, ZN => n12853);
   U7442 : NAND4_X1 port map( A1 => n12873, A2 => n12874, A3 => n12875, A4 => 
                           n12876, ZN => n12854);
   U7443 : AOI21_X1 port map( B1 => n16415, B2 => net226825, A => n12810, ZN =>
                           n12809);
   U7444 : NOR4_X1 port map( A1 => n12811, A2 => n12812, A3 => n12813, A4 => 
                           n12814, ZN => n12810);
   U7445 : NAND4_X1 port map( A1 => n12839, A2 => n12840, A3 => n12841, A4 => 
                           n12842, ZN => n12811);
   U7446 : NAND4_X1 port map( A1 => n12831, A2 => n12832, A3 => n12833, A4 => 
                           n12834, ZN => n12812);
   U7447 : AOI21_X1 port map( B1 => n16415, B2 => net226826, A => n12768, ZN =>
                           n12767);
   U7448 : NOR4_X1 port map( A1 => n12769, A2 => n12770, A3 => n12771, A4 => 
                           n12772, ZN => n12768);
   U7449 : NAND4_X1 port map( A1 => n12797, A2 => n12798, A3 => n12799, A4 => 
                           n12800, ZN => n12769);
   U7450 : NAND4_X1 port map( A1 => n12789, A2 => n12790, A3 => n12791, A4 => 
                           n12792, ZN => n12770);
   U7451 : AOI21_X1 port map( B1 => n16414, B2 => net226827, A => n12726, ZN =>
                           n12725);
   U7452 : NOR4_X1 port map( A1 => n12727, A2 => n12728, A3 => n12729, A4 => 
                           n12730, ZN => n12726);
   U7453 : NAND4_X1 port map( A1 => n12755, A2 => n12756, A3 => n12757, A4 => 
                           n12758, ZN => n12727);
   U7454 : NAND4_X1 port map( A1 => n12747, A2 => n12748, A3 => n12749, A4 => 
                           n12750, ZN => n12728);
   U7455 : AOI21_X1 port map( B1 => n16415, B2 => net226828, A => n12684, ZN =>
                           n12683);
   U7456 : NOR4_X1 port map( A1 => n12685, A2 => n12686, A3 => n12687, A4 => 
                           n12688, ZN => n12684);
   U7457 : NAND4_X1 port map( A1 => n12713, A2 => n12714, A3 => n12715, A4 => 
                           n12716, ZN => n12685);
   U7458 : NAND4_X1 port map( A1 => n12705, A2 => n12706, A3 => n12707, A4 => 
                           n12708, ZN => n12686);
   U7459 : AOI21_X1 port map( B1 => n16414, B2 => net226829, A => n12640, ZN =>
                           n12639);
   U7460 : NOR4_X1 port map( A1 => n12641, A2 => n12642, A3 => n12643, A4 => 
                           n12644, ZN => n12640);
   U7461 : NAND4_X1 port map( A1 => n12671, A2 => n12672, A3 => n12673, A4 => 
                           n12674, ZN => n12641);
   U7462 : NAND4_X1 port map( A1 => n12662, A2 => n12663, A3 => n12664, A4 => 
                           n12665, ZN => n12642);
   U7463 : AOI21_X1 port map( B1 => n16415, B2 => net226830, A => n12528, ZN =>
                           n12526);
   U7464 : NOR4_X1 port map( A1 => n12529, A2 => n12530, A3 => n12531, A4 => 
                           n12532, ZN => n12528);
   U7465 : NAND4_X1 port map( A1 => n12608, A2 => n12609, A3 => n12610, A4 => 
                           n12611, ZN => n12529);
   U7466 : NAND4_X1 port map( A1 => n12582, A2 => n12583, A3 => n12584, A4 => 
                           n12585, ZN => n12530);
   U7467 : AOI21_X1 port map( B1 => n16666, B2 => net226831, A => n12426, ZN =>
                           n12425);
   U7468 : NOR4_X1 port map( A1 => n12427, A2 => n12428, A3 => n12429, A4 => 
                           n12430, ZN => n12426);
   U7469 : NAND4_X1 port map( A1 => n12483, A2 => n12484, A3 => n12485, A4 => 
                           n12486, ZN => n12427);
   U7470 : NAND4_X1 port map( A1 => n12467, A2 => n12468, A3 => n12469, A4 => 
                           n12470, ZN => n12428);
   U7471 : AOI21_X1 port map( B1 => n16669, B2 => net226851, A => n12264, ZN =>
                           n12263);
   U7472 : NOR4_X1 port map( A1 => n12265, A2 => n12266, A3 => n12267, A4 => 
                           n12268, ZN => n12264);
   U7473 : NAND4_X1 port map( A1 => n12293, A2 => n12294, A3 => n12295, A4 => 
                           n12296, ZN => n12265);
   U7474 : NAND4_X1 port map( A1 => n12285, A2 => n12286, A3 => n12287, A4 => 
                           n12288, ZN => n12266);
   U7475 : AOI21_X1 port map( B1 => n16669, B2 => net226871, A => n12111, ZN =>
                           n12110);
   U7476 : NOR4_X1 port map( A1 => n12112, A2 => n12113, A3 => n12114, A4 => 
                           n12115, ZN => n12111);
   U7477 : NAND4_X1 port map( A1 => n12140, A2 => n12141, A3 => n12142, A4 => 
                           n12143, ZN => n12112);
   U7478 : NAND4_X1 port map( A1 => n12132, A2 => n12133, A3 => n12134, A4 => 
                           n12135, ZN => n12113);
   U7479 : AOI21_X1 port map( B1 => n16669, B2 => net226891, A => n11958, ZN =>
                           n11957);
   U7480 : NOR4_X1 port map( A1 => n11959, A2 => n11960, A3 => n11961, A4 => 
                           n11962, ZN => n11958);
   U7481 : NAND4_X1 port map( A1 => n11987, A2 => n11988, A3 => n11989, A4 => 
                           n11990, ZN => n11959);
   U7482 : NAND4_X1 port map( A1 => n11979, A2 => n11980, A3 => n11981, A4 => 
                           n11982, ZN => n11960);
   U7483 : AOI21_X1 port map( B1 => n16668, B2 => net226911, A => n11805, ZN =>
                           n11804);
   U7484 : NOR4_X1 port map( A1 => n11806, A2 => n11807, A3 => n11808, A4 => 
                           n11809, ZN => n11805);
   U7485 : NAND4_X1 port map( A1 => n11834, A2 => n11835, A3 => n11836, A4 => 
                           n11837, ZN => n11806);
   U7486 : NAND4_X1 port map( A1 => n11826, A2 => n11827, A3 => n11828, A4 => 
                           n11829, ZN => n11807);
   U7487 : AOI21_X1 port map( B1 => n16668, B2 => net226913, A => n11762, ZN =>
                           n11761);
   U7488 : NOR4_X1 port map( A1 => n11763, A2 => n11764, A3 => n11765, A4 => 
                           n11766, ZN => n11762);
   U7489 : NAND4_X1 port map( A1 => n11791, A2 => n11792, A3 => n11793, A4 => 
                           n11794, ZN => n11763);
   U7490 : NAND4_X1 port map( A1 => n11783, A2 => n11784, A3 => n11785, A4 => 
                           n11786, ZN => n11764);
   U7491 : AOI21_X1 port map( B1 => n16668, B2 => net226915, A => n11719, ZN =>
                           n11718);
   U7492 : NOR4_X1 port map( A1 => n11720, A2 => n11721, A3 => n11722, A4 => 
                           n11723, ZN => n11719);
   U7493 : NAND4_X1 port map( A1 => n11748, A2 => n11749, A3 => n11750, A4 => 
                           n11751, ZN => n11720);
   U7494 : NAND4_X1 port map( A1 => n11740, A2 => n11741, A3 => n11742, A4 => 
                           n11743, ZN => n11721);
   U7495 : AOI21_X1 port map( B1 => n16668, B2 => net226917, A => n11676, ZN =>
                           n11675);
   U7496 : NOR4_X1 port map( A1 => n11677, A2 => n11678, A3 => n11679, A4 => 
                           n11680, ZN => n11676);
   U7497 : NAND4_X1 port map( A1 => n11705, A2 => n11706, A3 => n11707, A4 => 
                           n11708, ZN => n11677);
   U7498 : NAND4_X1 port map( A1 => n11697, A2 => n11698, A3 => n11699, A4 => 
                           n11700, ZN => n11678);
   U7499 : AOI21_X1 port map( B1 => n16668, B2 => net226919, A => n11633, ZN =>
                           n11632);
   U7500 : NOR4_X1 port map( A1 => n11634, A2 => n11635, A3 => n11636, A4 => 
                           n11637, ZN => n11633);
   U7501 : NAND4_X1 port map( A1 => n11662, A2 => n11663, A3 => n11664, A4 => 
                           n11665, ZN => n11634);
   U7502 : NAND4_X1 port map( A1 => n11654, A2 => n11655, A3 => n11656, A4 => 
                           n11657, ZN => n11635);
   U7503 : AOI21_X1 port map( B1 => n16668, B2 => net226921, A => n11590, ZN =>
                           n11589);
   U7504 : NOR4_X1 port map( A1 => n11591, A2 => n11592, A3 => n11593, A4 => 
                           n11594, ZN => n11590);
   U7505 : NAND4_X1 port map( A1 => n11619, A2 => n11620, A3 => n11621, A4 => 
                           n11622, ZN => n11591);
   U7506 : NAND4_X1 port map( A1 => n11611, A2 => n11612, A3 => n11613, A4 => 
                           n11614, ZN => n11592);
   U7507 : AOI21_X1 port map( B1 => n16668, B2 => net226923, A => n11547, ZN =>
                           n11546);
   U7508 : NOR4_X1 port map( A1 => n11548, A2 => n11549, A3 => n11550, A4 => 
                           n11551, ZN => n11547);
   U7509 : NAND4_X1 port map( A1 => n11576, A2 => n11577, A3 => n11578, A4 => 
                           n11579, ZN => n11548);
   U7510 : NAND4_X1 port map( A1 => n11568, A2 => n11569, A3 => n11570, A4 => 
                           n11571, ZN => n11549);
   U7511 : AOI21_X1 port map( B1 => n16668, B2 => net226925, A => n11504, ZN =>
                           n11503);
   U7512 : NOR4_X1 port map( A1 => n11505, A2 => n11506, A3 => n11507, A4 => 
                           n11508, ZN => n11504);
   U7513 : NAND4_X1 port map( A1 => n11533, A2 => n11534, A3 => n11535, A4 => 
                           n11536, ZN => n11505);
   U7514 : NAND4_X1 port map( A1 => n11525, A2 => n11526, A3 => n11527, A4 => 
                           n11528, ZN => n11506);
   U7515 : AOI21_X1 port map( B1 => n16668, B2 => net226927, A => n11460, ZN =>
                           n11459);
   U7516 : NOR4_X1 port map( A1 => n11462, A2 => n11463, A3 => n11464, A4 => 
                           n11465, ZN => n11460);
   U7517 : NAND4_X1 port map( A1 => n11490, A2 => n11491, A3 => n11492, A4 => 
                           n11493, ZN => n11462);
   U7518 : NAND4_X1 port map( A1 => n11482, A2 => n11483, A3 => n11484, A4 => 
                           n11485, ZN => n11463);
   U7519 : AOI21_X1 port map( B1 => n16668, B2 => net226929, A => n11417, ZN =>
                           n11416);
   U7520 : NOR4_X1 port map( A1 => n11418, A2 => n11419, A3 => n11420, A4 => 
                           n11421, ZN => n11417);
   U7521 : NAND4_X1 port map( A1 => n11446, A2 => n11447, A3 => n11448, A4 => 
                           n11449, ZN => n11418);
   U7522 : NAND4_X1 port map( A1 => n11438, A2 => n11439, A3 => n11440, A4 => 
                           n11441, ZN => n11419);
   U7523 : AOI21_X1 port map( B1 => n16668, B2 => net226931, A => n11374, ZN =>
                           n11373);
   U7524 : NOR4_X1 port map( A1 => n11375, A2 => n11376, A3 => n11377, A4 => 
                           n11378, ZN => n11374);
   U7525 : NAND4_X1 port map( A1 => n11403, A2 => n11404, A3 => n11405, A4 => 
                           n11406, ZN => n11375);
   U7526 : NAND4_X1 port map( A1 => n11395, A2 => n11396, A3 => n11397, A4 => 
                           n11398, ZN => n11376);
   U7527 : AOI21_X1 port map( B1 => n16668, B2 => net226933, A => n11331, ZN =>
                           n11330);
   U7528 : NOR4_X1 port map( A1 => n11332, A2 => n11333, A3 => n11334, A4 => 
                           n11335, ZN => n11331);
   U7529 : NAND4_X1 port map( A1 => n11360, A2 => n11361, A3 => n11362, A4 => 
                           n11363, ZN => n11332);
   U7530 : NAND4_X1 port map( A1 => n11352, A2 => n11353, A3 => n11354, A4 => 
                           n11355, ZN => n11333);
   U7531 : AOI21_X1 port map( B1 => n16668, B2 => net226935, A => n11288, ZN =>
                           n11287);
   U7532 : NOR4_X1 port map( A1 => n11289, A2 => n11290, A3 => n11291, A4 => 
                           n11292, ZN => n11288);
   U7533 : NAND4_X1 port map( A1 => n11317, A2 => n11318, A3 => n11319, A4 => 
                           n11320, ZN => n11289);
   U7534 : NAND4_X1 port map( A1 => n11309, A2 => n11310, A3 => n11311, A4 => 
                           n11312, ZN => n11290);
   U7535 : AOI21_X1 port map( B1 => n16667, B2 => net226937, A => n11245, ZN =>
                           n11244);
   U7536 : NOR4_X1 port map( A1 => n11246, A2 => n11247, A3 => n11248, A4 => 
                           n11249, ZN => n11245);
   U7537 : NAND4_X1 port map( A1 => n11274, A2 => n11275, A3 => n11276, A4 => 
                           n11277, ZN => n11246);
   U7538 : NAND4_X1 port map( A1 => n11266, A2 => n11267, A3 => n11268, A4 => 
                           n11269, ZN => n11247);
   U7539 : AOI21_X1 port map( B1 => n16667, B2 => net226939, A => n11202, ZN =>
                           n11201);
   U7540 : NOR4_X1 port map( A1 => n11203, A2 => n11204, A3 => n11205, A4 => 
                           n11206, ZN => n11202);
   U7541 : NAND4_X1 port map( A1 => n11231, A2 => n11232, A3 => n11233, A4 => 
                           n11234, ZN => n11203);
   U7542 : NAND4_X1 port map( A1 => n11223, A2 => n11224, A3 => n11225, A4 => 
                           n11226, ZN => n11204);
   U7543 : AOI21_X1 port map( B1 => n16667, B2 => net226941, A => n11159, ZN =>
                           n11158);
   U7544 : NOR4_X1 port map( A1 => n11160, A2 => n11161, A3 => n11162, A4 => 
                           n11163, ZN => n11159);
   U7545 : NAND4_X1 port map( A1 => n11188, A2 => n11189, A3 => n11190, A4 => 
                           n11191, ZN => n11160);
   U7546 : NAND4_X1 port map( A1 => n11180, A2 => n11181, A3 => n11182, A4 => 
                           n11183, ZN => n11161);
   U7547 : AOI21_X1 port map( B1 => n16667, B2 => net226943, A => n11116, ZN =>
                           n11115);
   U7548 : NOR4_X1 port map( A1 => n11117, A2 => n11118, A3 => n11119, A4 => 
                           n11120, ZN => n11116);
   U7549 : NAND4_X1 port map( A1 => n11145, A2 => n11146, A3 => n11147, A4 => 
                           n11148, ZN => n11117);
   U7550 : NAND4_X1 port map( A1 => n11137, A2 => n11138, A3 => n11139, A4 => 
                           n11140, ZN => n11118);
   U7551 : AOI21_X1 port map( B1 => n16667, B2 => net226945, A => n11073, ZN =>
                           n11072);
   U7552 : NOR4_X1 port map( A1 => n11074, A2 => n11075, A3 => n11076, A4 => 
                           n11077, ZN => n11073);
   U7553 : NAND4_X1 port map( A1 => n11102, A2 => n11103, A3 => n11104, A4 => 
                           n11105, ZN => n11074);
   U7554 : NAND4_X1 port map( A1 => n11094, A2 => n11095, A3 => n11096, A4 => 
                           n11097, ZN => n11075);
   U7555 : AOI21_X1 port map( B1 => n16667, B2 => net226947, A => n11030, ZN =>
                           n11029);
   U7556 : NOR4_X1 port map( A1 => n11031, A2 => n11032, A3 => n11033, A4 => 
                           n11034, ZN => n11030);
   U7557 : NAND4_X1 port map( A1 => n11059, A2 => n11060, A3 => n11061, A4 => 
                           n11062, ZN => n11031);
   U7558 : NAND4_X1 port map( A1 => n11051, A2 => n11052, A3 => n11053, A4 => 
                           n11054, ZN => n11032);
   U7559 : AOI21_X1 port map( B1 => n16667, B2 => net226949, A => n10987, ZN =>
                           n10986);
   U7560 : NOR4_X1 port map( A1 => n10988, A2 => n10989, A3 => n10990, A4 => 
                           n10991, ZN => n10987);
   U7561 : NAND4_X1 port map( A1 => n11016, A2 => n11017, A3 => n11018, A4 => 
                           n11019, ZN => n10988);
   U7562 : NAND4_X1 port map( A1 => n11008, A2 => n11009, A3 => n11010, A4 => 
                           n11011, ZN => n10989);
   U7563 : AOI21_X1 port map( B1 => n16667, B2 => net226951, A => n10944, ZN =>
                           n10943);
   U7564 : NOR4_X1 port map( A1 => n10945, A2 => n10946, A3 => n10947, A4 => 
                           n10948, ZN => n10944);
   U7565 : NAND4_X1 port map( A1 => n10973, A2 => n10974, A3 => n10975, A4 => 
                           n10976, ZN => n10945);
   U7566 : NAND4_X1 port map( A1 => n10965, A2 => n10966, A3 => n10967, A4 => 
                           n10968, ZN => n10946);
   U7567 : AOI21_X1 port map( B1 => n16667, B2 => net226953, A => n10901, ZN =>
                           n10900);
   U7568 : NOR4_X1 port map( A1 => n10902, A2 => n10903, A3 => n10904, A4 => 
                           n10905, ZN => n10901);
   U7569 : NAND4_X1 port map( A1 => n10930, A2 => n10931, A3 => n10932, A4 => 
                           n10933, ZN => n10902);
   U7570 : NAND4_X1 port map( A1 => n10922, A2 => n10923, A3 => n10924, A4 => 
                           n10925, ZN => n10903);
   U7571 : AOI21_X1 port map( B1 => n16667, B2 => net226955, A => n10858, ZN =>
                           n10857);
   U7572 : NOR4_X1 port map( A1 => n10859, A2 => n10860, A3 => n10861, A4 => 
                           n10862, ZN => n10858);
   U7573 : NAND4_X1 port map( A1 => n10887, A2 => n10888, A3 => n10889, A4 => 
                           n10890, ZN => n10859);
   U7574 : NAND4_X1 port map( A1 => n10879, A2 => n10880, A3 => n10881, A4 => 
                           n10882, ZN => n10860);
   U7575 : AOI21_X1 port map( B1 => n16667, B2 => net226957, A => n10815, ZN =>
                           n10814);
   U7576 : NOR4_X1 port map( A1 => n10816, A2 => n10817, A3 => n10818, A4 => 
                           n10819, ZN => n10815);
   U7577 : NAND4_X1 port map( A1 => n10844, A2 => n10845, A3 => n10846, A4 => 
                           n10847, ZN => n10816);
   U7578 : NAND4_X1 port map( A1 => n10836, A2 => n10837, A3 => n10838, A4 => 
                           n10839, ZN => n10817);
   U7579 : AOI21_X1 port map( B1 => n16666, B2 => net226959, A => n10772, ZN =>
                           n10771);
   U7580 : NOR4_X1 port map( A1 => n10773, A2 => n10774, A3 => n10775, A4 => 
                           n10776, ZN => n10772);
   U7581 : NAND4_X1 port map( A1 => n10801, A2 => n10802, A3 => n10803, A4 => 
                           n10804, ZN => n10773);
   U7582 : NAND4_X1 port map( A1 => n10793, A2 => n10794, A3 => n10795, A4 => 
                           n10796, ZN => n10774);
   U7583 : AOI21_X1 port map( B1 => n16667, B2 => net226961, A => n10729, ZN =>
                           n10728);
   U7584 : NOR4_X1 port map( A1 => n10730, A2 => n10731, A3 => n10732, A4 => 
                           n10733, ZN => n10729);
   U7585 : NAND4_X1 port map( A1 => n10758, A2 => n10759, A3 => n10760, A4 => 
                           n10761, ZN => n10730);
   U7586 : NAND4_X1 port map( A1 => n10750, A2 => n10751, A3 => n10752, A4 => 
                           n10753, ZN => n10731);
   U7587 : AOI21_X1 port map( B1 => n16666, B2 => net226963, A => n10670, ZN =>
                           n10669);
   U7588 : NOR4_X1 port map( A1 => n10671, A2 => n10672, A3 => n10673, A4 => 
                           n10674, ZN => n10670);
   U7589 : NAND4_X1 port map( A1 => n10713, A2 => n10714, A3 => n10715, A4 => 
                           n10716, ZN => n10671);
   U7590 : NAND4_X1 port map( A1 => n10700, A2 => n10701, A3 => n10702, A4 => 
                           n10703, ZN => n10672);
   U7591 : AOI21_X1 port map( B1 => n16667, B2 => net226965, A => n10526, ZN =>
                           n10524);
   U7592 : NOR4_X1 port map( A1 => n10527, A2 => n10528, A3 => n10529, A4 => 
                           n10530, ZN => n10526);
   U7593 : NAND4_X1 port map( A1 => n10628, A2 => n10629, A3 => n10630, A4 => 
                           n10631, ZN => n10527);
   U7594 : NAND4_X1 port map( A1 => n10596, A2 => n10597, A3 => n10598, A4 => 
                           n10599, ZN => n10528);
   U7595 : NAND2_X1 port map( A1 => call, A2 => n14133, ZN => n14122);
   U7596 : NAND4_X1 port map( A1 => n12907, A2 => n12908, A3 => n12909, A4 => 
                           n12910, ZN => n12897);
   U7597 : AOI221_X1 port map( B1 => net227339, B2 => n16351, C1 => 
                           registers_30_24_port, C2 => n16348, A => n12912, ZN 
                           => n12909);
   U7598 : AOI221_X1 port map( B1 => registers_10_24_port, B2 => n16327, C1 => 
                           registers_0_24_port, C2 => n16324, A => n12914, ZN 
                           => n12907);
   U7599 : AOI221_X1 port map( B1 => net227338, B2 => n16339, C1 => 
                           registers_34_24_port, C2 => n16336, A => n12913, ZN 
                           => n12908);
   U7600 : NAND4_X1 port map( A1 => n12865, A2 => n12866, A3 => n12867, A4 => 
                           n12868, ZN => n12855);
   U7601 : AOI221_X1 port map( B1 => net227357, B2 => n16351, C1 => 
                           registers_30_25_port, C2 => n16348, A => n12870, ZN 
                           => n12867);
   U7602 : AOI221_X1 port map( B1 => registers_10_25_port, B2 => n16327, C1 => 
                           registers_0_25_port, C2 => n16324, A => n12872, ZN 
                           => n12865);
   U7603 : AOI221_X1 port map( B1 => net227356, B2 => n16339, C1 => 
                           registers_34_25_port, C2 => n16336, A => n12871, ZN 
                           => n12866);
   U7604 : NAND4_X1 port map( A1 => n12823, A2 => n12824, A3 => n12825, A4 => 
                           n12826, ZN => n12813);
   U7605 : AOI221_X1 port map( B1 => net227375, B2 => n16351, C1 => 
                           registers_30_26_port, C2 => n16348, A => n12828, ZN 
                           => n12825);
   U7606 : AOI221_X1 port map( B1 => registers_10_26_port, B2 => n16327, C1 => 
                           registers_0_26_port, C2 => n16324, A => n12830, ZN 
                           => n12823);
   U7607 : AOI221_X1 port map( B1 => net227374, B2 => n16339, C1 => 
                           registers_34_26_port, C2 => n16336, A => n12829, ZN 
                           => n12824);
   U7608 : NAND4_X1 port map( A1 => n12781, A2 => n12782, A3 => n12783, A4 => 
                           n12784, ZN => n12771);
   U7609 : AOI221_X1 port map( B1 => net227393, B2 => n16351, C1 => 
                           registers_30_27_port, C2 => n16348, A => n12786, ZN 
                           => n12783);
   U7610 : AOI221_X1 port map( B1 => registers_10_27_port, B2 => n16327, C1 => 
                           registers_0_27_port, C2 => n16324, A => n12788, ZN 
                           => n12781);
   U7611 : AOI221_X1 port map( B1 => net227392, B2 => n16339, C1 => 
                           registers_34_27_port, C2 => n16336, A => n12787, ZN 
                           => n12782);
   U7612 : NAND4_X1 port map( A1 => n12739, A2 => n12740, A3 => n12741, A4 => 
                           n12742, ZN => n12729);
   U7613 : AOI221_X1 port map( B1 => net227411, B2 => n16351, C1 => 
                           registers_30_28_port, C2 => n16348, A => n12744, ZN 
                           => n12741);
   U7614 : AOI221_X1 port map( B1 => registers_10_28_port, B2 => n16327, C1 => 
                           registers_0_28_port, C2 => n16324, A => n12746, ZN 
                           => n12739);
   U7615 : AOI221_X1 port map( B1 => net227410, B2 => n16339, C1 => 
                           registers_34_28_port, C2 => n16336, A => n12745, ZN 
                           => n12740);
   U7616 : NAND4_X1 port map( A1 => n12697, A2 => n12698, A3 => n12699, A4 => 
                           n12700, ZN => n12687);
   U7617 : AOI221_X1 port map( B1 => net227429, B2 => n16351, C1 => 
                           registers_30_29_port, C2 => n16348, A => n12702, ZN 
                           => n12699);
   U7618 : AOI221_X1 port map( B1 => registers_10_29_port, B2 => n16327, C1 => 
                           registers_0_29_port, C2 => n16324, A => n12704, ZN 
                           => n12697);
   U7619 : AOI221_X1 port map( B1 => net227428, B2 => n16339, C1 => 
                           registers_34_29_port, C2 => n16336, A => n12703, ZN 
                           => n12698);
   U7620 : NAND4_X1 port map( A1 => n12654, A2 => n12655, A3 => n12656, A4 => 
                           n12657, ZN => n12643);
   U7621 : AOI221_X1 port map( B1 => net227447, B2 => n16351, C1 => 
                           registers_30_30_port, C2 => n16348, A => n12659, ZN 
                           => n12656);
   U7622 : AOI221_X1 port map( B1 => registers_10_30_port, B2 => n16327, C1 => 
                           registers_0_30_port, C2 => n16324, A => n12661, ZN 
                           => n12654);
   U7623 : AOI221_X1 port map( B1 => net227446, B2 => n16339, C1 => 
                           registers_34_30_port, C2 => n16336, A => n12660, ZN 
                           => n12655);
   U7624 : NAND4_X1 port map( A1 => n12557, A2 => n12558, A3 => n12559, A4 => 
                           n12560, ZN => n12531);
   U7625 : AOI221_X1 port map( B1 => net227465, B2 => n16351, C1 => 
                           registers_30_31_port, C2 => n16348, A => n12569, ZN 
                           => n12559);
   U7626 : AOI221_X1 port map( B1 => registers_10_31_port, B2 => n16327, C1 => 
                           registers_0_31_port, C2 => n16324, A => n12579, ZN 
                           => n12557);
   U7627 : AOI221_X1 port map( B1 => net227464, B2 => n16339, C1 => 
                           registers_34_31_port, C2 => n16336, A => n12574, ZN 
                           => n12558);
   U7628 : NAND4_X1 port map( A1 => n10957, A2 => n10958, A3 => n10959, A4 => 
                           n10960, ZN => n10947);
   U7629 : AOI221_X1 port map( B1 => net227339, B2 => n16603, C1 => 
                           registers_30_24_port, C2 => n16600, A => n10962, ZN 
                           => n10959);
   U7630 : AOI221_X1 port map( B1 => registers_10_24_port, B2 => n16579, C1 => 
                           registers_0_24_port, C2 => n16576, A => n10964, ZN 
                           => n10957);
   U7631 : AOI221_X1 port map( B1 => net227338, B2 => n16591, C1 => 
                           registers_34_24_port, C2 => n16588, A => n10963, ZN 
                           => n10958);
   U7632 : NAND4_X1 port map( A1 => n10914, A2 => n10915, A3 => n10916, A4 => 
                           n10917, ZN => n10904);
   U7633 : AOI221_X1 port map( B1 => net227357, B2 => n16603, C1 => 
                           registers_30_25_port, C2 => n16600, A => n10919, ZN 
                           => n10916);
   U7634 : AOI221_X1 port map( B1 => registers_10_25_port, B2 => n16579, C1 => 
                           registers_0_25_port, C2 => n16576, A => n10921, ZN 
                           => n10914);
   U7635 : AOI221_X1 port map( B1 => net227356, B2 => n16591, C1 => 
                           registers_34_25_port, C2 => n16588, A => n10920, ZN 
                           => n10915);
   U7636 : NAND4_X1 port map( A1 => n10871, A2 => n10872, A3 => n10873, A4 => 
                           n10874, ZN => n10861);
   U7637 : AOI221_X1 port map( B1 => net227375, B2 => n16603, C1 => 
                           registers_30_26_port, C2 => n16600, A => n10876, ZN 
                           => n10873);
   U7638 : AOI221_X1 port map( B1 => registers_10_26_port, B2 => n16579, C1 => 
                           registers_0_26_port, C2 => n16576, A => n10878, ZN 
                           => n10871);
   U7639 : AOI221_X1 port map( B1 => net227374, B2 => n16591, C1 => 
                           registers_34_26_port, C2 => n16588, A => n10877, ZN 
                           => n10872);
   U7640 : NAND4_X1 port map( A1 => n10828, A2 => n10829, A3 => n10830, A4 => 
                           n10831, ZN => n10818);
   U7641 : AOI221_X1 port map( B1 => net227393, B2 => n16603, C1 => 
                           registers_30_27_port, C2 => n16600, A => n10833, ZN 
                           => n10830);
   U7642 : AOI221_X1 port map( B1 => registers_10_27_port, B2 => n16579, C1 => 
                           registers_0_27_port, C2 => n16576, A => n10835, ZN 
                           => n10828);
   U7643 : AOI221_X1 port map( B1 => net227392, B2 => n16591, C1 => 
                           registers_34_27_port, C2 => n16588, A => n10834, ZN 
                           => n10829);
   U7644 : NAND4_X1 port map( A1 => n10785, A2 => n10786, A3 => n10787, A4 => 
                           n10788, ZN => n10775);
   U7645 : AOI221_X1 port map( B1 => net227411, B2 => n16603, C1 => 
                           registers_30_28_port, C2 => n16600, A => n10790, ZN 
                           => n10787);
   U7646 : AOI221_X1 port map( B1 => registers_10_28_port, B2 => n16579, C1 => 
                           registers_0_28_port, C2 => n16576, A => n10792, ZN 
                           => n10785);
   U7647 : AOI221_X1 port map( B1 => net227410, B2 => n16591, C1 => 
                           registers_34_28_port, C2 => n16588, A => n10791, ZN 
                           => n10786);
   U7648 : NAND4_X1 port map( A1 => n10742, A2 => n10743, A3 => n10744, A4 => 
                           n10745, ZN => n10732);
   U7649 : AOI221_X1 port map( B1 => net227429, B2 => n16603, C1 => 
                           registers_30_29_port, C2 => n16600, A => n10747, ZN 
                           => n10744);
   U7650 : AOI221_X1 port map( B1 => registers_10_29_port, B2 => n16579, C1 => 
                           registers_0_29_port, C2 => n16576, A => n10749, ZN 
                           => n10742);
   U7651 : AOI221_X1 port map( B1 => net227428, B2 => n16591, C1 => 
                           registers_34_29_port, C2 => n16588, A => n10748, ZN 
                           => n10743);
   U7652 : NAND4_X1 port map( A1 => n10687, A2 => n10688, A3 => n10689, A4 => 
                           n10690, ZN => n10673);
   U7653 : AOI221_X1 port map( B1 => net227447, B2 => n16603, C1 => 
                           registers_30_30_port, C2 => n16600, A => n10694, ZN 
                           => n10689);
   U7654 : AOI221_X1 port map( B1 => registers_10_30_port, B2 => n16579, C1 => 
                           registers_0_30_port, C2 => n16576, A => n10698, ZN 
                           => n10687);
   U7655 : AOI221_X1 port map( B1 => net227446, B2 => n16591, C1 => 
                           registers_34_30_port, C2 => n16588, A => n10695, ZN 
                           => n10688);
   U7656 : NAND4_X1 port map( A1 => n10562, A2 => n10563, A3 => n10564, A4 => 
                           n10565, ZN => n10529);
   U7657 : AOI221_X1 port map( B1 => net227465, B2 => n16603, C1 => 
                           registers_30_31_port, C2 => n16600, A => n10577, ZN 
                           => n10564);
   U7658 : AOI221_X1 port map( B1 => registers_10_31_port, B2 => n16579, C1 => 
                           registers_0_31_port, C2 => n16576, A => n10591, ZN 
                           => n10562);
   U7659 : AOI221_X1 port map( B1 => net227464, B2 => n16591, C1 => 
                           registers_34_31_port, C2 => n16588, A => n10584, ZN 
                           => n10563);
   U7660 : NAND4_X1 port map( A1 => n5286, A2 => n5288, A3 => n5290, A4 => 
                           n5291, ZN => n5275);
   U7661 : AOI221_X1 port map( B1 => net227323, B2 => n17759, C1 => 
                           registers_25_23_port, C2 => n17756, A => n5293, ZN 
                           => n5290);
   U7662 : AOI221_X1 port map( B1 => registers_36_23_port, B2 => n17735, C1 => 
                           registers_38_23_port, C2 => n17732, A => n5295, ZN 
                           => n5286);
   U7663 : AOI221_X1 port map( B1 => net227318, B2 => n17771, C1 => 
                           registers_50_23_port, C2 => n17768, A => n5292, ZN 
                           => n5291);
   U7664 : NAND4_X1 port map( A1 => n5120, A2 => n5121, A3 => n5122, A4 => 
                           n5123, ZN => n5109);
   U7665 : AOI221_X1 port map( B1 => net227341, B2 => n17759, C1 => 
                           registers_25_24_port, C2 => n17756, A => n5125, ZN 
                           => n5122);
   U7666 : AOI221_X1 port map( B1 => registers_36_24_port, B2 => n17735, C1 => 
                           registers_38_24_port, C2 => n17732, A => n5129, ZN 
                           => n5120);
   U7667 : AOI221_X1 port map( B1 => net227336, B2 => n17771, C1 => 
                           registers_50_24_port, C2 => n17768, A => n5124, ZN 
                           => n5123);
   U7668 : NAND4_X1 port map( A1 => n5006, A2 => n5007, A3 => n5008, A4 => 
                           n5009, ZN => n4996);
   U7669 : AOI221_X1 port map( B1 => net227359, B2 => n17759, C1 => 
                           registers_25_25_port, C2 => n17756, A => n5011, ZN 
                           => n5008);
   U7670 : AOI221_X1 port map( B1 => registers_36_25_port, B2 => n17735, C1 => 
                           registers_38_25_port, C2 => n17732, A => n5013, ZN 
                           => n5006);
   U7671 : AOI221_X1 port map( B1 => net227354, B2 => n17771, C1 => 
                           registers_50_25_port, C2 => n17768, A => n5010, ZN 
                           => n5009);
   U7672 : NAND4_X1 port map( A1 => n4884, A2 => n4885, A3 => n4886, A4 => 
                           n4887, ZN => n4874);
   U7673 : AOI221_X1 port map( B1 => net227377, B2 => n17759, C1 => 
                           registers_25_26_port, C2 => n17756, A => n4889, ZN 
                           => n4886);
   U7674 : AOI221_X1 port map( B1 => registers_36_26_port, B2 => n17735, C1 => 
                           registers_38_26_port, C2 => n17732, A => n4891, ZN 
                           => n4884);
   U7675 : AOI221_X1 port map( B1 => net227372, B2 => n17771, C1 => 
                           registers_50_26_port, C2 => n17768, A => n4888, ZN 
                           => n4887);
   U7676 : NAND4_X1 port map( A1 => n4757, A2 => n4758, A3 => n4759, A4 => 
                           n4760, ZN => n4741);
   U7677 : AOI221_X1 port map( B1 => net227395, B2 => n17759, C1 => 
                           registers_25_27_port, C2 => n17756, A => n4762, ZN 
                           => n4759);
   U7678 : AOI221_X1 port map( B1 => registers_36_27_port, B2 => n17735, C1 => 
                           registers_38_27_port, C2 => n17732, A => n4764, ZN 
                           => n4757);
   U7679 : AOI221_X1 port map( B1 => net227390, B2 => n17771, C1 => 
                           registers_50_27_port, C2 => n17768, A => n4761, ZN 
                           => n4760);
   U7680 : NAND4_X1 port map( A1 => n4626, A2 => n4627, A3 => n4628, A4 => 
                           n4629, ZN => n4614);
   U7681 : AOI221_X1 port map( B1 => net227413, B2 => n17759, C1 => 
                           registers_25_28_port, C2 => n17756, A => n4631, ZN 
                           => n4628);
   U7682 : AOI221_X1 port map( B1 => registers_36_28_port, B2 => n17735, C1 => 
                           registers_38_28_port, C2 => n17732, A => n4633, ZN 
                           => n4626);
   U7683 : AOI221_X1 port map( B1 => net227408, B2 => n17771, C1 => 
                           registers_50_28_port, C2 => n17768, A => n4630, ZN 
                           => n4629);
   U7684 : NAND4_X1 port map( A1 => n4495, A2 => n4498, A3 => n4499, A4 => 
                           n4500, ZN => n4483);
   U7685 : AOI221_X1 port map( B1 => net227431, B2 => n17759, C1 => 
                           registers_25_29_port, C2 => n17756, A => n4502, ZN 
                           => n4499);
   U7686 : AOI221_X1 port map( B1 => registers_36_29_port, B2 => n17735, C1 => 
                           registers_38_29_port, C2 => n17732, A => n4506, ZN 
                           => n4495);
   U7687 : AOI221_X1 port map( B1 => net227426, B2 => n17771, C1 => 
                           registers_50_29_port, C2 => n17768, A => n4501, ZN 
                           => n4500);
   U7688 : NAND4_X1 port map( A1 => n4137, A2 => n4138, A3 => n4139, A4 => 
                           n4140, ZN => n4099);
   U7689 : AOI221_X1 port map( B1 => net227449, B2 => n17759, C1 => 
                           registers_25_30_port, C2 => n17756, A => n4156, ZN 
                           => n4139);
   U7690 : AOI221_X1 port map( B1 => registers_36_30_port, B2 => n17735, C1 => 
                           registers_38_30_port, C2 => n17732, A => n4172, ZN 
                           => n4137);
   U7691 : AOI221_X1 port map( B1 => net227444, B2 => n17771, C1 => 
                           registers_50_30_port, C2 => n17768, A => n4145, ZN 
                           => n4140);
   U7692 : NAND4_X1 port map( A1 => n13938, A2 => n13939, A3 => n13940, A4 => 
                           n13941, ZN => n13910);
   U7693 : AOI221_X1 port map( B1 => net226848, B2 => n16349, C1 => 
                           registers_30_0_port, C2 => n16346, A => n13943, ZN 
                           => n13940);
   U7694 : AOI221_X1 port map( B1 => registers_10_0_port, B2 => n16325, C1 => 
                           registers_0_0_port, C2 => n16322, A => n13947, ZN =>
                           n13938);
   U7695 : AOI221_X1 port map( B1 => net226847, B2 => n16337, C1 => 
                           registers_34_0_port, C2 => n16334, A => n13945, ZN 
                           => n13939);
   U7696 : NAND4_X1 port map( A1 => n13873, A2 => n13874, A3 => n13875, A4 => 
                           n13876, ZN => n13863);
   U7697 : AOI221_X1 port map( B1 => net226869, B2 => n16349, C1 => 
                           registers_30_1_port, C2 => n16346, A => n13878, ZN 
                           => n13875);
   U7698 : AOI221_X1 port map( B1 => registers_10_1_port, B2 => n16325, C1 => 
                           registers_0_1_port, C2 => n16322, A => n13880, ZN =>
                           n13873);
   U7699 : AOI221_X1 port map( B1 => net226868, B2 => n16337, C1 => 
                           registers_34_1_port, C2 => n16334, A => n13879, ZN 
                           => n13874);
   U7700 : NAND4_X1 port map( A1 => n13831, A2 => n13832, A3 => n13833, A4 => 
                           n13834, ZN => n13821);
   U7701 : AOI221_X1 port map( B1 => net226888, B2 => n16349, C1 => 
                           registers_30_2_port, C2 => n16346, A => n13836, ZN 
                           => n13833);
   U7702 : AOI221_X1 port map( B1 => registers_10_2_port, B2 => n16325, C1 => 
                           registers_0_2_port, C2 => n16322, A => n13838, ZN =>
                           n13831);
   U7703 : AOI221_X1 port map( B1 => net226880, B2 => n16337, C1 => 
                           registers_34_2_port, C2 => n16334, A => n13837, ZN 
                           => n13832);
   U7704 : NAND4_X1 port map( A1 => n13789, A2 => n13790, A3 => n13791, A4 => 
                           n13792, ZN => n13779);
   U7705 : AOI221_X1 port map( B1 => net226908, B2 => n16349, C1 => 
                           registers_30_3_port, C2 => n16346, A => n13794, ZN 
                           => n13791);
   U7706 : AOI221_X1 port map( B1 => registers_10_3_port, B2 => n16325, C1 => 
                           registers_0_3_port, C2 => n16322, A => n13796, ZN =>
                           n13789);
   U7707 : AOI221_X1 port map( B1 => net226900, B2 => n16337, C1 => 
                           registers_34_3_port, C2 => n16334, A => n13795, ZN 
                           => n13790);
   U7708 : NAND4_X1 port map( A1 => n13747, A2 => n13748, A3 => n13749, A4 => 
                           n13750, ZN => n13737);
   U7709 : AOI221_X1 port map( B1 => net226982, B2 => n16349, C1 => 
                           registers_30_4_port, C2 => n16346, A => n13752, ZN 
                           => n13749);
   U7710 : AOI221_X1 port map( B1 => registers_10_4_port, B2 => n16325, C1 => 
                           registers_0_4_port, C2 => n16322, A => n13754, ZN =>
                           n13747);
   U7711 : AOI221_X1 port map( B1 => net226973, B2 => n16337, C1 => 
                           registers_34_4_port, C2 => n16334, A => n13753, ZN 
                           => n13748);
   U7712 : NAND4_X1 port map( A1 => n13705, A2 => n13706, A3 => n13707, A4 => 
                           n13708, ZN => n13695);
   U7713 : AOI221_X1 port map( B1 => net226991, B2 => n16349, C1 => 
                           registers_30_5_port, C2 => n16346, A => n13710, ZN 
                           => n13707);
   U7714 : AOI221_X1 port map( B1 => registers_10_5_port, B2 => n16325, C1 => 
                           registers_0_5_port, C2 => n16322, A => n13712, ZN =>
                           n13705);
   U7715 : AOI221_X1 port map( B1 => net226990, B2 => n16337, C1 => 
                           registers_34_5_port, C2 => n16334, A => n13711, ZN 
                           => n13706);
   U7716 : NAND4_X1 port map( A1 => n13663, A2 => n13664, A3 => n13665, A4 => 
                           n13666, ZN => n13653);
   U7717 : AOI221_X1 port map( B1 => net227015, B2 => n16349, C1 => 
                           registers_30_6_port, C2 => n16346, A => n13668, ZN 
                           => n13665);
   U7718 : AOI221_X1 port map( B1 => registers_10_6_port, B2 => n16325, C1 => 
                           registers_0_6_port, C2 => n16322, A => n13670, ZN =>
                           n13663);
   U7719 : AOI221_X1 port map( B1 => net227014, B2 => n16337, C1 => 
                           registers_34_6_port, C2 => n16334, A => n13669, ZN 
                           => n13664);
   U7720 : NAND4_X1 port map( A1 => n13621, A2 => n13622, A3 => n13623, A4 => 
                           n13624, ZN => n13611);
   U7721 : AOI221_X1 port map( B1 => net227033, B2 => n16349, C1 => 
                           registers_30_7_port, C2 => n16346, A => n13626, ZN 
                           => n13623);
   U7722 : AOI221_X1 port map( B1 => registers_10_7_port, B2 => n16325, C1 => 
                           registers_0_7_port, C2 => n16322, A => n13628, ZN =>
                           n13621);
   U7723 : AOI221_X1 port map( B1 => net227032, B2 => n16337, C1 => 
                           registers_34_7_port, C2 => n16334, A => n13627, ZN 
                           => n13622);
   U7724 : NAND4_X1 port map( A1 => n13579, A2 => n13580, A3 => n13581, A4 => 
                           n13582, ZN => n13569);
   U7725 : AOI221_X1 port map( B1 => net227051, B2 => n16349, C1 => 
                           registers_30_8_port, C2 => n16346, A => n13584, ZN 
                           => n13581);
   U7726 : AOI221_X1 port map( B1 => registers_10_8_port, B2 => n16325, C1 => 
                           registers_0_8_port, C2 => n16322, A => n13586, ZN =>
                           n13579);
   U7727 : AOI221_X1 port map( B1 => net227050, B2 => n16337, C1 => 
                           registers_34_8_port, C2 => n16334, A => n13585, ZN 
                           => n13580);
   U7728 : NAND4_X1 port map( A1 => n13537, A2 => n13538, A3 => n13539, A4 => 
                           n13540, ZN => n13527);
   U7729 : AOI221_X1 port map( B1 => net227069, B2 => n16349, C1 => 
                           registers_30_9_port, C2 => n16346, A => n13542, ZN 
                           => n13539);
   U7730 : AOI221_X1 port map( B1 => registers_10_9_port, B2 => n16325, C1 => 
                           registers_0_9_port, C2 => n16322, A => n13544, ZN =>
                           n13537);
   U7731 : AOI221_X1 port map( B1 => net227068, B2 => n16337, C1 => 
                           registers_34_9_port, C2 => n16334, A => n13543, ZN 
                           => n13538);
   U7732 : NAND4_X1 port map( A1 => n13495, A2 => n13496, A3 => n13497, A4 => 
                           n13498, ZN => n13485);
   U7733 : AOI221_X1 port map( B1 => net227087, B2 => n16349, C1 => 
                           registers_30_10_port, C2 => n16346, A => n13500, ZN 
                           => n13497);
   U7734 : AOI221_X1 port map( B1 => registers_10_10_port, B2 => n16325, C1 => 
                           registers_0_10_port, C2 => n16322, A => n13502, ZN 
                           => n13495);
   U7735 : AOI221_X1 port map( B1 => net227086, B2 => n16337, C1 => 
                           registers_34_10_port, C2 => n16334, A => n13501, ZN 
                           => n13496);
   U7736 : NAND4_X1 port map( A1 => n13453, A2 => n13454, A3 => n13455, A4 => 
                           n13456, ZN => n13443);
   U7737 : AOI221_X1 port map( B1 => net227105, B2 => n16349, C1 => 
                           registers_30_11_port, C2 => n16346, A => n13458, ZN 
                           => n13455);
   U7738 : AOI221_X1 port map( B1 => registers_10_11_port, B2 => n16325, C1 => 
                           registers_0_11_port, C2 => n16322, A => n13460, ZN 
                           => n13453);
   U7739 : AOI221_X1 port map( B1 => net227104, B2 => n16337, C1 => 
                           registers_34_11_port, C2 => n16334, A => n13459, ZN 
                           => n13454);
   U7740 : NAND4_X1 port map( A1 => n13411, A2 => n13412, A3 => n13413, A4 => 
                           n13414, ZN => n13401);
   U7741 : AOI221_X1 port map( B1 => net227123, B2 => n16350, C1 => 
                           registers_30_12_port, C2 => n16347, A => n13416, ZN 
                           => n13413);
   U7742 : AOI221_X1 port map( B1 => registers_10_12_port, B2 => n16326, C1 => 
                           registers_0_12_port, C2 => n16323, A => n13418, ZN 
                           => n13411);
   U7743 : AOI221_X1 port map( B1 => net227122, B2 => n16338, C1 => 
                           registers_34_12_port, C2 => n16335, A => n13417, ZN 
                           => n13412);
   U7744 : NAND4_X1 port map( A1 => n13369, A2 => n13370, A3 => n13371, A4 => 
                           n13372, ZN => n13359);
   U7745 : AOI221_X1 port map( B1 => net227141, B2 => n16350, C1 => 
                           registers_30_13_port, C2 => n16347, A => n13374, ZN 
                           => n13371);
   U7746 : AOI221_X1 port map( B1 => registers_10_13_port, B2 => n16326, C1 => 
                           registers_0_13_port, C2 => n16323, A => n13376, ZN 
                           => n13369);
   U7747 : AOI221_X1 port map( B1 => net227140, B2 => n16338, C1 => 
                           registers_34_13_port, C2 => n16335, A => n13375, ZN 
                           => n13370);
   U7748 : NAND4_X1 port map( A1 => n13327, A2 => n13328, A3 => n13329, A4 => 
                           n13330, ZN => n13317);
   U7749 : AOI221_X1 port map( B1 => net227159, B2 => n16350, C1 => 
                           registers_30_14_port, C2 => n16347, A => n13332, ZN 
                           => n13329);
   U7750 : AOI221_X1 port map( B1 => registers_10_14_port, B2 => n16326, C1 => 
                           registers_0_14_port, C2 => n16323, A => n13334, ZN 
                           => n13327);
   U7751 : AOI221_X1 port map( B1 => net227158, B2 => n16338, C1 => 
                           registers_34_14_port, C2 => n16335, A => n13333, ZN 
                           => n13328);
   U7752 : NAND4_X1 port map( A1 => n13285, A2 => n13286, A3 => n13287, A4 => 
                           n13288, ZN => n13275);
   U7753 : AOI221_X1 port map( B1 => net227177, B2 => n16350, C1 => 
                           registers_30_15_port, C2 => n16347, A => n13290, ZN 
                           => n13287);
   U7754 : AOI221_X1 port map( B1 => registers_10_15_port, B2 => n16326, C1 => 
                           registers_0_15_port, C2 => n16323, A => n13292, ZN 
                           => n13285);
   U7755 : AOI221_X1 port map( B1 => net227176, B2 => n16338, C1 => 
                           registers_34_15_port, C2 => n16335, A => n13291, ZN 
                           => n13286);
   U7756 : NAND4_X1 port map( A1 => n13243, A2 => n13244, A3 => n13245, A4 => 
                           n13246, ZN => n13233);
   U7757 : AOI221_X1 port map( B1 => net227195, B2 => n16350, C1 => 
                           registers_30_16_port, C2 => n16347, A => n13248, ZN 
                           => n13245);
   U7758 : AOI221_X1 port map( B1 => registers_10_16_port, B2 => n16326, C1 => 
                           registers_0_16_port, C2 => n16323, A => n13250, ZN 
                           => n13243);
   U7759 : AOI221_X1 port map( B1 => net227194, B2 => n16338, C1 => 
                           registers_34_16_port, C2 => n16335, A => n13249, ZN 
                           => n13244);
   U7760 : NAND4_X1 port map( A1 => n13201, A2 => n13202, A3 => n13203, A4 => 
                           n13204, ZN => n13191);
   U7761 : AOI221_X1 port map( B1 => net227213, B2 => n16350, C1 => 
                           registers_30_17_port, C2 => n16347, A => n13206, ZN 
                           => n13203);
   U7762 : AOI221_X1 port map( B1 => registers_10_17_port, B2 => n16326, C1 => 
                           registers_0_17_port, C2 => n16323, A => n13208, ZN 
                           => n13201);
   U7763 : AOI221_X1 port map( B1 => net227212, B2 => n16338, C1 => 
                           registers_34_17_port, C2 => n16335, A => n13207, ZN 
                           => n13202);
   U7764 : NAND4_X1 port map( A1 => n13159, A2 => n13160, A3 => n13161, A4 => 
                           n13162, ZN => n13149);
   U7765 : AOI221_X1 port map( B1 => net227231, B2 => n16350, C1 => 
                           registers_30_18_port, C2 => n16347, A => n13164, ZN 
                           => n13161);
   U7766 : AOI221_X1 port map( B1 => registers_10_18_port, B2 => n16326, C1 => 
                           registers_0_18_port, C2 => n16323, A => n13166, ZN 
                           => n13159);
   U7767 : AOI221_X1 port map( B1 => net227230, B2 => n16338, C1 => 
                           registers_34_18_port, C2 => n16335, A => n13165, ZN 
                           => n13160);
   U7768 : NAND4_X1 port map( A1 => n13117, A2 => n13118, A3 => n13119, A4 => 
                           n13120, ZN => n13107);
   U7769 : AOI221_X1 port map( B1 => net227249, B2 => n16350, C1 => 
                           registers_30_19_port, C2 => n16347, A => n13122, ZN 
                           => n13119);
   U7770 : AOI221_X1 port map( B1 => registers_10_19_port, B2 => n16326, C1 => 
                           registers_0_19_port, C2 => n16323, A => n13124, ZN 
                           => n13117);
   U7771 : AOI221_X1 port map( B1 => net227248, B2 => n16338, C1 => 
                           registers_34_19_port, C2 => n16335, A => n13123, ZN 
                           => n13118);
   U7772 : NAND4_X1 port map( A1 => n13075, A2 => n13076, A3 => n13077, A4 => 
                           n13078, ZN => n13065);
   U7773 : AOI221_X1 port map( B1 => net227267, B2 => n16350, C1 => 
                           registers_30_20_port, C2 => n16347, A => n13080, ZN 
                           => n13077);
   U7774 : AOI221_X1 port map( B1 => registers_10_20_port, B2 => n16326, C1 => 
                           registers_0_20_port, C2 => n16323, A => n13082, ZN 
                           => n13075);
   U7775 : AOI221_X1 port map( B1 => net227266, B2 => n16338, C1 => 
                           registers_34_20_port, C2 => n16335, A => n13081, ZN 
                           => n13076);
   U7776 : NAND4_X1 port map( A1 => n13033, A2 => n13034, A3 => n13035, A4 => 
                           n13036, ZN => n13023);
   U7777 : AOI221_X1 port map( B1 => net227285, B2 => n16350, C1 => 
                           registers_30_21_port, C2 => n16347, A => n13038, ZN 
                           => n13035);
   U7778 : AOI221_X1 port map( B1 => registers_10_21_port, B2 => n16326, C1 => 
                           registers_0_21_port, C2 => n16323, A => n13040, ZN 
                           => n13033);
   U7779 : AOI221_X1 port map( B1 => net227284, B2 => n16338, C1 => 
                           registers_34_21_port, C2 => n16335, A => n13039, ZN 
                           => n13034);
   U7780 : NAND4_X1 port map( A1 => n12991, A2 => n12992, A3 => n12993, A4 => 
                           n12994, ZN => n12981);
   U7781 : AOI221_X1 port map( B1 => net227303, B2 => n16350, C1 => 
                           registers_30_22_port, C2 => n16347, A => n12996, ZN 
                           => n12993);
   U7782 : AOI221_X1 port map( B1 => registers_10_22_port, B2 => n16326, C1 => 
                           registers_0_22_port, C2 => n16323, A => n12998, ZN 
                           => n12991);
   U7783 : AOI221_X1 port map( B1 => net227302, B2 => n16338, C1 => 
                           registers_34_22_port, C2 => n16335, A => n12997, ZN 
                           => n12992);
   U7784 : NAND4_X1 port map( A1 => n12949, A2 => n12950, A3 => n12951, A4 => 
                           n12952, ZN => n12939);
   U7785 : AOI221_X1 port map( B1 => net227321, B2 => n16350, C1 => 
                           registers_30_23_port, C2 => n16347, A => n12954, ZN 
                           => n12951);
   U7786 : AOI221_X1 port map( B1 => registers_10_23_port, B2 => n16326, C1 => 
                           registers_0_23_port, C2 => n16323, A => n12956, ZN 
                           => n12949);
   U7787 : AOI221_X1 port map( B1 => net227320, B2 => n16338, C1 => 
                           registers_34_23_port, C2 => n16335, A => n12955, ZN 
                           => n12950);
   U7788 : NAND4_X1 port map( A1 => n12457, A2 => n12458, A3 => n12459, A4 => 
                           n12460, ZN => n12429);
   U7789 : AOI221_X1 port map( B1 => net226848, B2 => n16601, C1 => 
                           registers_30_0_port, C2 => n16598, A => n12462, ZN 
                           => n12459);
   U7790 : AOI221_X1 port map( B1 => registers_10_0_port, B2 => n16577, C1 => 
                           registers_0_0_port, C2 => n16574, A => n12466, ZN =>
                           n12457);
   U7791 : AOI221_X1 port map( B1 => net226847, B2 => n16589, C1 => 
                           registers_34_0_port, C2 => n16586, A => n12464, ZN 
                           => n12458);
   U7792 : NAND4_X1 port map( A1 => n12277, A2 => n12278, A3 => n12279, A4 => 
                           n12280, ZN => n12267);
   U7793 : AOI221_X1 port map( B1 => net226869, B2 => n16601, C1 => 
                           registers_30_1_port, C2 => n16598, A => n12282, ZN 
                           => n12279);
   U7794 : AOI221_X1 port map( B1 => registers_10_1_port, B2 => n16577, C1 => 
                           registers_0_1_port, C2 => n16574, A => n12284, ZN =>
                           n12277);
   U7795 : AOI221_X1 port map( B1 => net226868, B2 => n16589, C1 => 
                           registers_34_1_port, C2 => n16586, A => n12283, ZN 
                           => n12278);
   U7796 : NAND4_X1 port map( A1 => n12124, A2 => n12125, A3 => n12126, A4 => 
                           n12127, ZN => n12114);
   U7797 : AOI221_X1 port map( B1 => net226888, B2 => n16601, C1 => 
                           registers_30_2_port, C2 => n16598, A => n12129, ZN 
                           => n12126);
   U7798 : AOI221_X1 port map( B1 => registers_10_2_port, B2 => n16577, C1 => 
                           registers_0_2_port, C2 => n16574, A => n12131, ZN =>
                           n12124);
   U7799 : AOI221_X1 port map( B1 => net226880, B2 => n16589, C1 => 
                           registers_34_2_port, C2 => n16586, A => n12130, ZN 
                           => n12125);
   U7800 : NAND4_X1 port map( A1 => n11971, A2 => n11972, A3 => n11973, A4 => 
                           n11974, ZN => n11961);
   U7801 : AOI221_X1 port map( B1 => net226908, B2 => n16601, C1 => 
                           registers_30_3_port, C2 => n16598, A => n11976, ZN 
                           => n11973);
   U7802 : AOI221_X1 port map( B1 => registers_10_3_port, B2 => n16577, C1 => 
                           registers_0_3_port, C2 => n16574, A => n11978, ZN =>
                           n11971);
   U7803 : AOI221_X1 port map( B1 => net226900, B2 => n16589, C1 => 
                           registers_34_3_port, C2 => n16586, A => n11977, ZN 
                           => n11972);
   U7804 : NAND4_X1 port map( A1 => n11818, A2 => n11819, A3 => n11820, A4 => 
                           n11821, ZN => n11808);
   U7805 : AOI221_X1 port map( B1 => net226982, B2 => n16601, C1 => 
                           registers_30_4_port, C2 => n16598, A => n11823, ZN 
                           => n11820);
   U7806 : AOI221_X1 port map( B1 => registers_10_4_port, B2 => n16577, C1 => 
                           registers_0_4_port, C2 => n16574, A => n11825, ZN =>
                           n11818);
   U7807 : AOI221_X1 port map( B1 => net226973, B2 => n16589, C1 => 
                           registers_34_4_port, C2 => n16586, A => n11824, ZN 
                           => n11819);
   U7808 : NAND4_X1 port map( A1 => n11775, A2 => n11776, A3 => n11777, A4 => 
                           n11778, ZN => n11765);
   U7809 : AOI221_X1 port map( B1 => net226991, B2 => n16601, C1 => 
                           registers_30_5_port, C2 => n16598, A => n11780, ZN 
                           => n11777);
   U7810 : AOI221_X1 port map( B1 => registers_10_5_port, B2 => n16577, C1 => 
                           registers_0_5_port, C2 => n16574, A => n11782, ZN =>
                           n11775);
   U7811 : AOI221_X1 port map( B1 => net226990, B2 => n16589, C1 => 
                           registers_34_5_port, C2 => n16586, A => n11781, ZN 
                           => n11776);
   U7812 : NAND4_X1 port map( A1 => n11732, A2 => n11733, A3 => n11734, A4 => 
                           n11735, ZN => n11722);
   U7813 : AOI221_X1 port map( B1 => net227015, B2 => n16601, C1 => 
                           registers_30_6_port, C2 => n16598, A => n11737, ZN 
                           => n11734);
   U7814 : AOI221_X1 port map( B1 => registers_10_6_port, B2 => n16577, C1 => 
                           registers_0_6_port, C2 => n16574, A => n11739, ZN =>
                           n11732);
   U7815 : AOI221_X1 port map( B1 => net227014, B2 => n16589, C1 => 
                           registers_34_6_port, C2 => n16586, A => n11738, ZN 
                           => n11733);
   U7816 : NAND4_X1 port map( A1 => n11689, A2 => n11690, A3 => n11691, A4 => 
                           n11692, ZN => n11679);
   U7817 : AOI221_X1 port map( B1 => net227033, B2 => n16601, C1 => 
                           registers_30_7_port, C2 => n16598, A => n11694, ZN 
                           => n11691);
   U7818 : AOI221_X1 port map( B1 => registers_10_7_port, B2 => n16577, C1 => 
                           registers_0_7_port, C2 => n16574, A => n11696, ZN =>
                           n11689);
   U7819 : AOI221_X1 port map( B1 => net227032, B2 => n16589, C1 => 
                           registers_34_7_port, C2 => n16586, A => n11695, ZN 
                           => n11690);
   U7820 : NAND4_X1 port map( A1 => n11646, A2 => n11647, A3 => n11648, A4 => 
                           n11649, ZN => n11636);
   U7821 : AOI221_X1 port map( B1 => net227051, B2 => n16601, C1 => 
                           registers_30_8_port, C2 => n16598, A => n11651, ZN 
                           => n11648);
   U7822 : AOI221_X1 port map( B1 => registers_10_8_port, B2 => n16577, C1 => 
                           registers_0_8_port, C2 => n16574, A => n11653, ZN =>
                           n11646);
   U7823 : AOI221_X1 port map( B1 => net227050, B2 => n16589, C1 => 
                           registers_34_8_port, C2 => n16586, A => n11652, ZN 
                           => n11647);
   U7824 : NAND4_X1 port map( A1 => n11603, A2 => n11604, A3 => n11605, A4 => 
                           n11606, ZN => n11593);
   U7825 : AOI221_X1 port map( B1 => net227069, B2 => n16601, C1 => 
                           registers_30_9_port, C2 => n16598, A => n11608, ZN 
                           => n11605);
   U7826 : AOI221_X1 port map( B1 => registers_10_9_port, B2 => n16577, C1 => 
                           registers_0_9_port, C2 => n16574, A => n11610, ZN =>
                           n11603);
   U7827 : AOI221_X1 port map( B1 => net227068, B2 => n16589, C1 => 
                           registers_34_9_port, C2 => n16586, A => n11609, ZN 
                           => n11604);
   U7828 : NAND4_X1 port map( A1 => n11560, A2 => n11561, A3 => n11562, A4 => 
                           n11563, ZN => n11550);
   U7829 : AOI221_X1 port map( B1 => net227087, B2 => n16601, C1 => 
                           registers_30_10_port, C2 => n16598, A => n11565, ZN 
                           => n11562);
   U7830 : AOI221_X1 port map( B1 => registers_10_10_port, B2 => n16577, C1 => 
                           registers_0_10_port, C2 => n16574, A => n11567, ZN 
                           => n11560);
   U7831 : AOI221_X1 port map( B1 => net227086, B2 => n16589, C1 => 
                           registers_34_10_port, C2 => n16586, A => n11566, ZN 
                           => n11561);
   U7832 : NAND4_X1 port map( A1 => n11517, A2 => n11518, A3 => n11519, A4 => 
                           n11520, ZN => n11507);
   U7833 : AOI221_X1 port map( B1 => net227105, B2 => n16601, C1 => 
                           registers_30_11_port, C2 => n16598, A => n11522, ZN 
                           => n11519);
   U7834 : AOI221_X1 port map( B1 => registers_10_11_port, B2 => n16577, C1 => 
                           registers_0_11_port, C2 => n16574, A => n11524, ZN 
                           => n11517);
   U7835 : AOI221_X1 port map( B1 => net227104, B2 => n16589, C1 => 
                           registers_34_11_port, C2 => n16586, A => n11523, ZN 
                           => n11518);
   U7836 : NAND4_X1 port map( A1 => n11474, A2 => n11475, A3 => n11476, A4 => 
                           n11477, ZN => n11464);
   U7837 : AOI221_X1 port map( B1 => net227123, B2 => n16602, C1 => 
                           registers_30_12_port, C2 => n16599, A => n11479, ZN 
                           => n11476);
   U7838 : AOI221_X1 port map( B1 => registers_10_12_port, B2 => n16578, C1 => 
                           registers_0_12_port, C2 => n16575, A => n11481, ZN 
                           => n11474);
   U7839 : AOI221_X1 port map( B1 => net227122, B2 => n16590, C1 => 
                           registers_34_12_port, C2 => n16587, A => n11480, ZN 
                           => n11475);
   U7840 : NAND4_X1 port map( A1 => n11430, A2 => n11431, A3 => n11432, A4 => 
                           n11433, ZN => n11420);
   U7841 : AOI221_X1 port map( B1 => net227141, B2 => n16602, C1 => 
                           registers_30_13_port, C2 => n16599, A => n11435, ZN 
                           => n11432);
   U7842 : AOI221_X1 port map( B1 => registers_10_13_port, B2 => n16578, C1 => 
                           registers_0_13_port, C2 => n16575, A => n11437, ZN 
                           => n11430);
   U7843 : AOI221_X1 port map( B1 => net227140, B2 => n16590, C1 => 
                           registers_34_13_port, C2 => n16587, A => n11436, ZN 
                           => n11431);
   U7844 : NAND4_X1 port map( A1 => n11387, A2 => n11388, A3 => n11389, A4 => 
                           n11390, ZN => n11377);
   U7845 : AOI221_X1 port map( B1 => net227159, B2 => n16602, C1 => 
                           registers_30_14_port, C2 => n16599, A => n11392, ZN 
                           => n11389);
   U7846 : AOI221_X1 port map( B1 => registers_10_14_port, B2 => n16578, C1 => 
                           registers_0_14_port, C2 => n16575, A => n11394, ZN 
                           => n11387);
   U7847 : AOI221_X1 port map( B1 => net227158, B2 => n16590, C1 => 
                           registers_34_14_port, C2 => n16587, A => n11393, ZN 
                           => n11388);
   U7848 : NAND4_X1 port map( A1 => n11344, A2 => n11345, A3 => n11346, A4 => 
                           n11347, ZN => n11334);
   U7849 : AOI221_X1 port map( B1 => net227177, B2 => n16602, C1 => 
                           registers_30_15_port, C2 => n16599, A => n11349, ZN 
                           => n11346);
   U7850 : AOI221_X1 port map( B1 => registers_10_15_port, B2 => n16578, C1 => 
                           registers_0_15_port, C2 => n16575, A => n11351, ZN 
                           => n11344);
   U7851 : AOI221_X1 port map( B1 => net227176, B2 => n16590, C1 => 
                           registers_34_15_port, C2 => n16587, A => n11350, ZN 
                           => n11345);
   U7852 : NAND4_X1 port map( A1 => n11301, A2 => n11302, A3 => n11303, A4 => 
                           n11304, ZN => n11291);
   U7853 : AOI221_X1 port map( B1 => net227195, B2 => n16602, C1 => 
                           registers_30_16_port, C2 => n16599, A => n11306, ZN 
                           => n11303);
   U7854 : AOI221_X1 port map( B1 => registers_10_16_port, B2 => n16578, C1 => 
                           registers_0_16_port, C2 => n16575, A => n11308, ZN 
                           => n11301);
   U7855 : AOI221_X1 port map( B1 => net227194, B2 => n16590, C1 => 
                           registers_34_16_port, C2 => n16587, A => n11307, ZN 
                           => n11302);
   U7856 : NAND4_X1 port map( A1 => n11258, A2 => n11259, A3 => n11260, A4 => 
                           n11261, ZN => n11248);
   U7857 : AOI221_X1 port map( B1 => net227213, B2 => n16602, C1 => 
                           registers_30_17_port, C2 => n16599, A => n11263, ZN 
                           => n11260);
   U7858 : AOI221_X1 port map( B1 => registers_10_17_port, B2 => n16578, C1 => 
                           registers_0_17_port, C2 => n16575, A => n11265, ZN 
                           => n11258);
   U7859 : AOI221_X1 port map( B1 => net227212, B2 => n16590, C1 => 
                           registers_34_17_port, C2 => n16587, A => n11264, ZN 
                           => n11259);
   U7860 : NAND4_X1 port map( A1 => n11215, A2 => n11216, A3 => n11217, A4 => 
                           n11218, ZN => n11205);
   U7861 : AOI221_X1 port map( B1 => net227231, B2 => n16602, C1 => 
                           registers_30_18_port, C2 => n16599, A => n11220, ZN 
                           => n11217);
   U7862 : AOI221_X1 port map( B1 => registers_10_18_port, B2 => n16578, C1 => 
                           registers_0_18_port, C2 => n16575, A => n11222, ZN 
                           => n11215);
   U7863 : AOI221_X1 port map( B1 => net227230, B2 => n16590, C1 => 
                           registers_34_18_port, C2 => n16587, A => n11221, ZN 
                           => n11216);
   U7864 : NAND4_X1 port map( A1 => n11172, A2 => n11173, A3 => n11174, A4 => 
                           n11175, ZN => n11162);
   U7865 : AOI221_X1 port map( B1 => net227249, B2 => n16602, C1 => 
                           registers_30_19_port, C2 => n16599, A => n11177, ZN 
                           => n11174);
   U7866 : AOI221_X1 port map( B1 => registers_10_19_port, B2 => n16578, C1 => 
                           registers_0_19_port, C2 => n16575, A => n11179, ZN 
                           => n11172);
   U7867 : AOI221_X1 port map( B1 => net227248, B2 => n16590, C1 => 
                           registers_34_19_port, C2 => n16587, A => n11178, ZN 
                           => n11173);
   U7868 : NAND4_X1 port map( A1 => n11129, A2 => n11130, A3 => n11131, A4 => 
                           n11132, ZN => n11119);
   U7869 : AOI221_X1 port map( B1 => net227267, B2 => n16602, C1 => 
                           registers_30_20_port, C2 => n16599, A => n11134, ZN 
                           => n11131);
   U7870 : AOI221_X1 port map( B1 => registers_10_20_port, B2 => n16578, C1 => 
                           registers_0_20_port, C2 => n16575, A => n11136, ZN 
                           => n11129);
   U7871 : AOI221_X1 port map( B1 => net227266, B2 => n16590, C1 => 
                           registers_34_20_port, C2 => n16587, A => n11135, ZN 
                           => n11130);
   U7872 : NAND4_X1 port map( A1 => n11086, A2 => n11087, A3 => n11088, A4 => 
                           n11089, ZN => n11076);
   U7873 : AOI221_X1 port map( B1 => net227285, B2 => n16602, C1 => 
                           registers_30_21_port, C2 => n16599, A => n11091, ZN 
                           => n11088);
   U7874 : AOI221_X1 port map( B1 => registers_10_21_port, B2 => n16578, C1 => 
                           registers_0_21_port, C2 => n16575, A => n11093, ZN 
                           => n11086);
   U7875 : AOI221_X1 port map( B1 => net227284, B2 => n16590, C1 => 
                           registers_34_21_port, C2 => n16587, A => n11092, ZN 
                           => n11087);
   U7876 : NAND4_X1 port map( A1 => n11043, A2 => n11044, A3 => n11045, A4 => 
                           n11046, ZN => n11033);
   U7877 : AOI221_X1 port map( B1 => net227303, B2 => n16602, C1 => 
                           registers_30_22_port, C2 => n16599, A => n11048, ZN 
                           => n11045);
   U7878 : AOI221_X1 port map( B1 => registers_10_22_port, B2 => n16578, C1 => 
                           registers_0_22_port, C2 => n16575, A => n11050, ZN 
                           => n11043);
   U7879 : AOI221_X1 port map( B1 => net227302, B2 => n16590, C1 => 
                           registers_34_22_port, C2 => n16587, A => n11049, ZN 
                           => n11044);
   U7880 : NAND4_X1 port map( A1 => n11000, A2 => n11001, A3 => n11002, A4 => 
                           n11003, ZN => n10990);
   U7881 : AOI221_X1 port map( B1 => net227321, B2 => n16602, C1 => 
                           registers_30_23_port, C2 => n16599, A => n11005, ZN 
                           => n11002);
   U7882 : AOI221_X1 port map( B1 => registers_10_23_port, B2 => n16578, C1 => 
                           registers_0_23_port, C2 => n16575, A => n11007, ZN 
                           => n11000);
   U7883 : AOI221_X1 port map( B1 => net227320, B2 => n16590, C1 => 
                           registers_34_23_port, C2 => n16587, A => n11006, ZN 
                           => n11001);
   U7884 : NAND4_X1 port map( A1 => n12383, A2 => n12384, A3 => n12385, A4 => 
                           n12386, ZN => n12373);
   U7885 : AOI221_X1 port map( B1 => net226840, B2 => n17757, C1 => 
                           registers_25_0_port, C2 => n17754, A => n12388, ZN 
                           => n12385);
   U7886 : AOI221_X1 port map( B1 => net226837, B2 => n17769, C1 => 
                           registers_50_0_port, C2 => n17766, A => n12387, ZN 
                           => n12386);
   U7887 : AOI221_X1 port map( B1 => registers_36_0_port, B2 => n17733, C1 => 
                           registers_38_0_port, C2 => n17730, A => n12390, ZN 
                           => n12383);
   U7888 : NAND4_X1 port map( A1 => n12229, A2 => n12230, A3 => n12231, A4 => 
                           n12232, ZN => n12219);
   U7889 : AOI221_X1 port map( B1 => net226862, B2 => n17757, C1 => 
                           registers_25_1_port, C2 => n17754, A => n12234, ZN 
                           => n12231);
   U7890 : AOI221_X1 port map( B1 => net226860, B2 => n17769, C1 => 
                           registers_50_1_port, C2 => n17766, A => n12233, ZN 
                           => n12232);
   U7891 : AOI221_X1 port map( B1 => registers_36_1_port, B2 => n17733, C1 => 
                           registers_38_1_port, C2 => n17730, A => n12236, ZN 
                           => n12229);
   U7892 : NAND4_X1 port map( A1 => n12074, A2 => n12075, A3 => n12076, A4 => 
                           n12077, ZN => n12064);
   U7893 : AOI221_X1 port map( B1 => net226881, B2 => n17757, C1 => 
                           registers_25_2_port, C2 => n17754, A => n12079, ZN 
                           => n12076);
   U7894 : AOI221_X1 port map( B1 => net226886, B2 => n17769, C1 => 
                           registers_50_2_port, C2 => n17766, A => n12078, ZN 
                           => n12077);
   U7895 : AOI221_X1 port map( B1 => registers_36_2_port, B2 => n17733, C1 => 
                           registers_38_2_port, C2 => n17730, A => n12081, ZN 
                           => n12074);
   U7896 : NAND4_X1 port map( A1 => n11921, A2 => n11922, A3 => n11923, A4 => 
                           n11924, ZN => n11911);
   U7897 : AOI221_X1 port map( B1 => net226910, B2 => n17757, C1 => 
                           registers_25_3_port, C2 => n17754, A => n11926, ZN 
                           => n11923);
   U7898 : AOI221_X1 port map( B1 => net226899, B2 => n17769, C1 => 
                           registers_50_3_port, C2 => n17766, A => n11925, ZN 
                           => n11924);
   U7899 : AOI221_X1 port map( B1 => registers_36_3_port, B2 => n17733, C1 => 
                           registers_38_3_port, C2 => n17730, A => n11928, ZN 
                           => n11921);
   U7900 : NAND4_X1 port map( A1 => n10478, A2 => n10479, A3 => n10480, A4 => 
                           n10481, ZN => n10468);
   U7901 : AOI221_X1 port map( B1 => net226984, B2 => n17757, C1 => 
                           registers_25_4_port, C2 => n17754, A => n10483, ZN 
                           => n10480);
   U7902 : AOI221_X1 port map( B1 => net226981, B2 => n17769, C1 => 
                           registers_50_4_port, C2 => n17766, A => n10482, ZN 
                           => n10481);
   U7903 : AOI221_X1 port map( B1 => registers_36_4_port, B2 => n17733, C1 => 
                           registers_38_4_port, C2 => n17730, A => n10485, ZN 
                           => n10478);
   U7904 : NAND4_X1 port map( A1 => n10368, A2 => n10369, A3 => n10370, A4 => 
                           n10371, ZN => n10358);
   U7905 : AOI221_X1 port map( B1 => net226993, B2 => n17757, C1 => 
                           registers_25_5_port, C2 => n17754, A => n10373, ZN 
                           => n10370);
   U7906 : AOI221_X1 port map( B1 => net227001, B2 => n17769, C1 => 
                           registers_50_5_port, C2 => n17766, A => n10372, ZN 
                           => n10371);
   U7907 : AOI221_X1 port map( B1 => registers_36_5_port, B2 => n17733, C1 => 
                           registers_38_5_port, C2 => n17730, A => n10375, ZN 
                           => n10368);
   U7908 : NAND4_X1 port map( A1 => n10256, A2 => n10257, A3 => n10258, A4 => 
                           n10259, ZN => n10246);
   U7909 : AOI221_X1 port map( B1 => net227017, B2 => n17757, C1 => 
                           registers_25_6_port, C2 => n17754, A => n10261, ZN 
                           => n10258);
   U7910 : AOI221_X1 port map( B1 => net227012, B2 => n17769, C1 => 
                           registers_50_6_port, C2 => n17766, A => n10260, ZN 
                           => n10259);
   U7911 : AOI221_X1 port map( B1 => registers_36_6_port, B2 => n17733, C1 => 
                           registers_38_6_port, C2 => n17730, A => n10263, ZN 
                           => n10256);
   U7912 : NAND4_X1 port map( A1 => n7620, A2 => n7621, A3 => n7622, A4 => 
                           n7623, ZN => n7610);
   U7913 : AOI221_X1 port map( B1 => net227035, B2 => n17757, C1 => 
                           registers_25_7_port, C2 => n17754, A => n7625, ZN =>
                           n7622);
   U7914 : AOI221_X1 port map( B1 => net227030, B2 => n17769, C1 => 
                           registers_50_7_port, C2 => n17766, A => n7624, ZN =>
                           n7623);
   U7915 : AOI221_X1 port map( B1 => registers_36_7_port, B2 => n17733, C1 => 
                           registers_38_7_port, C2 => n17730, A => n7627, ZN =>
                           n7620);
   U7916 : NAND4_X1 port map( A1 => n7505, A2 => n7506, A3 => n7507, A4 => 
                           n7508, ZN => n7495);
   U7917 : AOI221_X1 port map( B1 => net227053, B2 => n17757, C1 => 
                           registers_25_8_port, C2 => n17754, A => n7510, ZN =>
                           n7507);
   U7918 : AOI221_X1 port map( B1 => net227048, B2 => n17769, C1 => 
                           registers_50_8_port, C2 => n17766, A => n7509, ZN =>
                           n7508);
   U7919 : AOI221_X1 port map( B1 => registers_36_8_port, B2 => n17733, C1 => 
                           registers_38_8_port, C2 => n17730, A => n7512, ZN =>
                           n7505);
   U7920 : NAND4_X1 port map( A1 => n7396, A2 => n7397, A3 => n7398, A4 => 
                           n7399, ZN => n7386);
   U7921 : AOI221_X1 port map( B1 => net227071, B2 => n17757, C1 => 
                           registers_25_9_port, C2 => n17754, A => n7401, ZN =>
                           n7398);
   U7922 : AOI221_X1 port map( B1 => net227066, B2 => n17769, C1 => 
                           registers_50_9_port, C2 => n17766, A => n7400, ZN =>
                           n7399);
   U7923 : AOI221_X1 port map( B1 => registers_36_9_port, B2 => n17733, C1 => 
                           registers_38_9_port, C2 => n17730, A => n7403, ZN =>
                           n7396);
   U7924 : NAND4_X1 port map( A1 => n7287, A2 => n7288, A3 => n7289, A4 => 
                           n7290, ZN => n7277);
   U7925 : AOI221_X1 port map( B1 => net227089, B2 => n17757, C1 => 
                           registers_25_10_port, C2 => n17754, A => n7292, ZN 
                           => n7289);
   U7926 : AOI221_X1 port map( B1 => net227084, B2 => n17769, C1 => 
                           registers_50_10_port, C2 => n17766, A => n7291, ZN 
                           => n7290);
   U7927 : AOI221_X1 port map( B1 => registers_36_10_port, B2 => n17733, C1 => 
                           registers_38_10_port, C2 => n17730, A => n7294, ZN 
                           => n7287);
   U7928 : NAND4_X1 port map( A1 => n7173, A2 => n7174, A3 => n7175, A4 => 
                           n7176, ZN => n7163);
   U7929 : AOI221_X1 port map( B1 => net227107, B2 => n17758, C1 => 
                           registers_25_11_port, C2 => n17755, A => n7178, ZN 
                           => n7175);
   U7930 : AOI221_X1 port map( B1 => net227102, B2 => n17770, C1 => 
                           registers_50_11_port, C2 => n17767, A => n7177, ZN 
                           => n7176);
   U7931 : AOI221_X1 port map( B1 => registers_36_11_port, B2 => n17734, C1 => 
                           registers_38_11_port, C2 => n17731, A => n7180, ZN 
                           => n7173);
   U7932 : NAND4_X1 port map( A1 => n7064, A2 => n7065, A3 => n7066, A4 => 
                           n7067, ZN => n7054);
   U7933 : AOI221_X1 port map( B1 => net227125, B2 => n17758, C1 => 
                           registers_25_12_port, C2 => n17755, A => n7069, ZN 
                           => n7066);
   U7934 : AOI221_X1 port map( B1 => net227120, B2 => n17770, C1 => 
                           registers_50_12_port, C2 => n17767, A => n7068, ZN 
                           => n7067);
   U7935 : AOI221_X1 port map( B1 => registers_36_12_port, B2 => n17734, C1 => 
                           registers_38_12_port, C2 => n17731, A => n7071, ZN 
                           => n7064);
   U7936 : NAND4_X1 port map( A1 => n6955, A2 => n6956, A3 => n6957, A4 => 
                           n6958, ZN => n6945);
   U7937 : AOI221_X1 port map( B1 => net227143, B2 => n17758, C1 => 
                           registers_25_13_port, C2 => n17755, A => n6960, ZN 
                           => n6957);
   U7938 : AOI221_X1 port map( B1 => net227138, B2 => n17770, C1 => 
                           registers_50_13_port, C2 => n17767, A => n6959, ZN 
                           => n6958);
   U7939 : AOI221_X1 port map( B1 => registers_36_13_port, B2 => n17734, C1 => 
                           registers_38_13_port, C2 => n17731, A => n6962, ZN 
                           => n6955);
   U7940 : NAND4_X1 port map( A1 => n6846, A2 => n6847, A3 => n6848, A4 => 
                           n6849, ZN => n6836);
   U7941 : AOI221_X1 port map( B1 => net227161, B2 => n17758, C1 => 
                           registers_25_14_port, C2 => n17755, A => n6851, ZN 
                           => n6848);
   U7942 : AOI221_X1 port map( B1 => net227156, B2 => n17770, C1 => 
                           registers_50_14_port, C2 => n17767, A => n6850, ZN 
                           => n6849);
   U7943 : AOI221_X1 port map( B1 => registers_36_14_port, B2 => n17734, C1 => 
                           registers_38_14_port, C2 => n17731, A => n6853, ZN 
                           => n6846);
   U7944 : NAND4_X1 port map( A1 => n6737, A2 => n6738, A3 => n6739, A4 => 
                           n6740, ZN => n6727);
   U7945 : AOI221_X1 port map( B1 => net227179, B2 => n17758, C1 => 
                           registers_25_15_port, C2 => n17755, A => n6742, ZN 
                           => n6739);
   U7946 : AOI221_X1 port map( B1 => net227174, B2 => n17770, C1 => 
                           registers_50_15_port, C2 => n17767, A => n6741, ZN 
                           => n6740);
   U7947 : AOI221_X1 port map( B1 => registers_36_15_port, B2 => n17734, C1 => 
                           registers_38_15_port, C2 => n17731, A => n6744, ZN 
                           => n6737);
   U7948 : NAND4_X1 port map( A1 => n6577, A2 => n6580, A3 => n6581, A4 => 
                           n6582, ZN => n6564);
   U7949 : AOI221_X1 port map( B1 => net227197, B2 => n17758, C1 => 
                           registers_25_16_port, C2 => n17755, A => n6599, ZN 
                           => n6581);
   U7950 : AOI221_X1 port map( B1 => net227192, B2 => n17770, C1 => 
                           registers_50_16_port, C2 => n17767, A => n6598, ZN 
                           => n6582);
   U7951 : AOI221_X1 port map( B1 => registers_36_16_port, B2 => n17734, C1 => 
                           registers_38_16_port, C2 => n17731, A => n6601, ZN 
                           => n6577);
   U7952 : NAND4_X1 port map( A1 => n6392, A2 => n6393, A3 => n6409, A4 => 
                           n6410, ZN => n6377);
   U7953 : AOI221_X1 port map( B1 => net227215, B2 => n17758, C1 => 
                           registers_25_17_port, C2 => n17755, A => n6412, ZN 
                           => n6409);
   U7954 : AOI221_X1 port map( B1 => net227210, B2 => n17770, C1 => 
                           registers_50_17_port, C2 => n17767, A => n6411, ZN 
                           => n6410);
   U7955 : AOI221_X1 port map( B1 => registers_36_17_port, B2 => n17734, C1 => 
                           registers_38_17_port, C2 => n17731, A => n6414, ZN 
                           => n6392);
   U7956 : NAND4_X1 port map( A1 => n6220, A2 => n6221, A3 => n6222, A4 => 
                           n6223, ZN => n6192);
   U7957 : AOI221_X1 port map( B1 => net227233, B2 => n17758, C1 => 
                           registers_25_18_port, C2 => n17755, A => n6225, ZN 
                           => n6222);
   U7958 : AOI221_X1 port map( B1 => net227228, B2 => n17770, C1 => 
                           registers_50_18_port, C2 => n17767, A => n6224, ZN 
                           => n6223);
   U7959 : AOI221_X1 port map( B1 => registers_36_18_port, B2 => n17734, C1 => 
                           registers_38_18_port, C2 => n17731, A => n6227, ZN 
                           => n6220);
   U7960 : NAND4_X1 port map( A1 => n6033, A2 => n6034, A3 => n6035, A4 => 
                           n6036, ZN => n6006);
   U7961 : AOI221_X1 port map( B1 => net227251, B2 => n17758, C1 => 
                           registers_25_19_port, C2 => n17755, A => n6038, ZN 
                           => n6035);
   U7962 : AOI221_X1 port map( B1 => net227246, B2 => n17770, C1 => 
                           registers_50_19_port, C2 => n17767, A => n6037, ZN 
                           => n6036);
   U7963 : AOI221_X1 port map( B1 => registers_36_19_port, B2 => n17734, C1 => 
                           registers_38_19_port, C2 => n17731, A => n6040, ZN 
                           => n6033);
   U7964 : NAND4_X1 port map( A1 => n5846, A2 => n5847, A3 => n5848, A4 => 
                           n5849, ZN => n5819);
   U7965 : AOI221_X1 port map( B1 => net227269, B2 => n17758, C1 => 
                           registers_25_20_port, C2 => n17755, A => n5851, ZN 
                           => n5848);
   U7966 : AOI221_X1 port map( B1 => net227264, B2 => n17770, C1 => 
                           registers_50_20_port, C2 => n17767, A => n5850, ZN 
                           => n5849);
   U7967 : AOI221_X1 port map( B1 => registers_36_20_port, B2 => n17734, C1 => 
                           registers_38_20_port, C2 => n17731, A => n5854, ZN 
                           => n5846);
   U7968 : NAND4_X1 port map( A1 => n5659, A2 => n5660, A3 => n5661, A4 => 
                           n5662, ZN => n5632);
   U7969 : AOI221_X1 port map( B1 => net227287, B2 => n17758, C1 => 
                           registers_25_21_port, C2 => n17755, A => n5665, ZN 
                           => n5661);
   U7970 : AOI221_X1 port map( B1 => net227282, B2 => n17770, C1 => 
                           registers_50_21_port, C2 => n17767, A => n5664, ZN 
                           => n5662);
   U7971 : AOI221_X1 port map( B1 => registers_36_21_port, B2 => n17734, C1 => 
                           registers_38_21_port, C2 => n17731, A => n5669, ZN 
                           => n5659);
   U7972 : NAND4_X1 port map( A1 => n5472, A2 => n5473, A3 => n5475, A4 => 
                           n5476, ZN => n5447);
   U7973 : AOI221_X1 port map( B1 => net227305, B2 => n17758, C1 => 
                           registers_25_22_port, C2 => n17755, A => n5480, ZN 
                           => n5475);
   U7974 : AOI221_X1 port map( B1 => net227300, B2 => n17770, C1 => 
                           registers_50_22_port, C2 => n17767, A => n5478, ZN 
                           => n5476);
   U7975 : AOI221_X1 port map( B1 => registers_36_22_port, B2 => n17734, C1 => 
                           registers_38_22_port, C2 => n17731, A => n5482, ZN 
                           => n5472);
   U7976 : NAND4_X1 port map( A1 => n14109, A2 => n14110, A3 => n14111, A4 => 
                           n14112, ZN => n14078);
   U7977 : AOI221_X1 port map( B1 => net227467, B2 => n17757, C1 => 
                           registers_25_31_port, C2 => n17754, A => n14126, ZN 
                           => n14111);
   U7978 : AOI221_X1 port map( B1 => net227462, B2 => n17769, C1 => 
                           registers_50_31_port, C2 => n17766, A => n14113, ZN 
                           => n14112);
   U7979 : AOI221_X1 port map( B1 => registers_36_31_port, B2 => n17733, C1 => 
                           registers_38_31_port, C2 => n17730, A => n14148, ZN 
                           => n14109);
   U7980 : NAND2_X1 port map( A1 => n14129, A2 => call, ZN => n14115);
   U7981 : NAND4_X1 port map( A1 => n5298, A2 => n5299, A3 => n5301, A4 => 
                           n5302, ZN => n5274);
   U7982 : AOI221_X1 port map( B1 => net227316, B2 => n17711, C1 => net227315, 
                           C2 => n17708, A => n5304, ZN => n5301);
   U7983 : AOI221_X1 port map( B1 => net227317, B2 => n17723, C1 => 
                           registers_54_23_port, C2 => n17720, A => n5303, ZN 
                           => n5302);
   U7984 : AOI221_X1 port map( B1 => registers_42_23_port, B2 => n17687, C1 => 
                           registers_43_23_port, C2 => n17684, A => n5307, ZN 
                           => n5298);
   U7985 : NAND4_X1 port map( A1 => n5130, A2 => n5131, A3 => n5132, A4 => 
                           n5133, ZN => n5108);
   U7986 : AOI221_X1 port map( B1 => net227334, B2 => n17711, C1 => net227333, 
                           C2 => n17708, A => n5135, ZN => n5132);
   U7987 : AOI221_X1 port map( B1 => net227335, B2 => n17723, C1 => 
                           registers_54_24_port, C2 => n17720, A => n5134, ZN 
                           => n5133);
   U7988 : AOI221_X1 port map( B1 => registers_42_24_port, B2 => n17687, C1 => 
                           registers_43_24_port, C2 => n17684, A => n5137, ZN 
                           => n5130);
   U7989 : NAND4_X1 port map( A1 => n5014, A2 => n5015, A3 => n5016, A4 => 
                           n5017, ZN => n4995);
   U7990 : AOI221_X1 port map( B1 => net227352, B2 => n17711, C1 => net227351, 
                           C2 => n17708, A => n5021, ZN => n5016);
   U7991 : AOI221_X1 port map( B1 => net227353, B2 => n17723, C1 => 
                           registers_54_25_port, C2 => n17720, A => n5020, ZN 
                           => n5017);
   U7992 : AOI221_X1 port map( B1 => registers_42_25_port, B2 => n17687, C1 => 
                           registers_43_25_port, C2 => n17684, A => n5023, ZN 
                           => n5014);
   U7993 : NAND4_X1 port map( A1 => n4892, A2 => n4895, A3 => n4898, A4 => 
                           n4899, ZN => n4873);
   U7994 : AOI221_X1 port map( B1 => net227370, B2 => n17711, C1 => net227369, 
                           C2 => n17708, A => n4901, ZN => n4898);
   U7995 : AOI221_X1 port map( B1 => net227371, B2 => n17723, C1 => 
                           registers_54_26_port, C2 => n17720, A => n4900, ZN 
                           => n4899);
   U7996 : AOI221_X1 port map( B1 => registers_42_26_port, B2 => n17687, C1 => 
                           registers_43_26_port, C2 => n17684, A => n4903, ZN 
                           => n4892);
   U7997 : NAND4_X1 port map( A1 => n4767, A2 => n4768, A3 => n4769, A4 => 
                           n4770, ZN => n4740);
   U7998 : AOI221_X1 port map( B1 => net227388, B2 => n17711, C1 => net227387, 
                           C2 => n17708, A => n4772, ZN => n4769);
   U7999 : AOI221_X1 port map( B1 => net227389, B2 => n17723, C1 => 
                           registers_54_27_port, C2 => n17720, A => n4771, ZN 
                           => n4770);
   U8000 : AOI221_X1 port map( B1 => registers_42_27_port, B2 => n17687, C1 => 
                           registers_43_27_port, C2 => n17684, A => n4774, ZN 
                           => n4767);
   U8001 : NAND4_X1 port map( A1 => n4634, A2 => n4635, A3 => n4636, A4 => 
                           n4637, ZN => n4613);
   U8002 : AOI221_X1 port map( B1 => net227406, B2 => n17711, C1 => net227405, 
                           C2 => n17708, A => n4639, ZN => n4636);
   U8003 : AOI221_X1 port map( B1 => net227407, B2 => n17723, C1 => 
                           registers_54_28_port, C2 => n17720, A => n4638, ZN 
                           => n4637);
   U8004 : AOI221_X1 port map( B1 => registers_42_28_port, B2 => n17687, C1 => 
                           registers_43_28_port, C2 => n17684, A => n4641, ZN 
                           => n4634);
   U8005 : NAND4_X1 port map( A1 => n4507, A2 => n4508, A3 => n4509, A4 => 
                           n4510, ZN => n4482);
   U8006 : AOI221_X1 port map( B1 => net227424, B2 => n17711, C1 => net227423, 
                           C2 => n17708, A => n4512, ZN => n4509);
   U8007 : AOI221_X1 port map( B1 => net227425, B2 => n17723, C1 => 
                           registers_54_29_port, C2 => n17720, A => n4511, ZN 
                           => n4510);
   U8008 : AOI221_X1 port map( B1 => registers_42_29_port, B2 => n17687, C1 => 
                           registers_43_29_port, C2 => n17684, A => n4514, ZN 
                           => n4507);
   U8009 : NAND4_X1 port map( A1 => n4177, A2 => n4178, A3 => n4179, A4 => 
                           n4180, ZN => n4098);
   U8010 : AOI221_X1 port map( B1 => net227442, B2 => n17711, C1 => net227441, 
                           C2 => n17708, A => n4190, ZN => n4179);
   U8011 : AOI221_X1 port map( B1 => net227443, B2 => n17723, C1 => 
                           registers_54_30_port, C2 => n17720, A => n4183, ZN 
                           => n4180);
   U8012 : AOI221_X1 port map( B1 => registers_42_30_port, B2 => n17687, C1 => 
                           registers_43_30_port, C2 => n17684, A => n4208, ZN 
                           => n4177);
   U8013 : NAND4_X1 port map( A1 => n12391, A2 => n12392, A3 => n12393, A4 => 
                           n12394, ZN => n12372);
   U8014 : AOI221_X1 port map( B1 => net226845, B2 => n17709, C1 => net226836, 
                           C2 => n17706, A => n12396, ZN => n12393);
   U8015 : AOI221_X1 port map( B1 => net226846, B2 => n17721, C1 => 
                           registers_54_0_port, C2 => n17718, A => n12395, ZN 
                           => n12394);
   U8016 : AOI221_X1 port map( B1 => registers_42_0_port, B2 => n17685, C1 => 
                           registers_43_0_port, C2 => n17682, A => n12398, ZN 
                           => n12391);
   U8017 : NAND4_X1 port map( A1 => n12237, A2 => n12238, A3 => n12239, A4 => 
                           n12240, ZN => n12218);
   U8018 : AOI221_X1 port map( B1 => net226858, B2 => n17709, C1 => net226866, 
                           C2 => n17706, A => n12242, ZN => n12239);
   U8019 : AOI221_X1 port map( B1 => net226859, B2 => n17721, C1 => 
                           registers_54_1_port, C2 => n17718, A => n12241, ZN 
                           => n12240);
   U8020 : AOI221_X1 port map( B1 => registers_42_1_port, B2 => n17685, C1 => 
                           registers_43_1_port, C2 => n17682, A => n12244, ZN 
                           => n12237);
   U8021 : NAND4_X1 port map( A1 => n12082, A2 => n12083, A3 => n12084, A4 => 
                           n12085, ZN => n12063);
   U8022 : AOI221_X1 port map( B1 => net226879, B2 => n17709, C1 => net226878, 
                           C2 => n17706, A => n12087, ZN => n12084);
   U8023 : AOI221_X1 port map( B1 => net226885, B2 => n17721, C1 => 
                           registers_54_2_port, C2 => n17718, A => n12086, ZN 
                           => n12085);
   U8024 : AOI221_X1 port map( B1 => registers_42_2_port, B2 => n17685, C1 => 
                           registers_43_2_port, C2 => n17682, A => n12089, ZN 
                           => n12082);
   U8025 : NAND4_X1 port map( A1 => n11929, A2 => n11930, A3 => n11931, A4 => 
                           n11932, ZN => n11910);
   U8026 : AOI221_X1 port map( B1 => net226906, B2 => n17709, C1 => net226905, 
                           C2 => n17706, A => n11934, ZN => n11931);
   U8027 : AOI221_X1 port map( B1 => net226898, B2 => n17721, C1 => 
                           registers_54_3_port, C2 => n17718, A => n11933, ZN 
                           => n11932);
   U8028 : AOI221_X1 port map( B1 => registers_42_3_port, B2 => n17685, C1 => 
                           registers_43_3_port, C2 => n17682, A => n11936, ZN 
                           => n11929);
   U8029 : NAND4_X1 port map( A1 => n10486, A2 => n10487, A3 => n10488, A4 => 
                           n10489, ZN => n10467);
   U8030 : AOI221_X1 port map( B1 => net226979, B2 => n17709, C1 => net226978, 
                           C2 => n17706, A => n10491, ZN => n10488);
   U8031 : AOI221_X1 port map( B1 => net226980, B2 => n17721, C1 => 
                           registers_54_4_port, C2 => n17718, A => n10490, ZN 
                           => n10489);
   U8032 : AOI221_X1 port map( B1 => registers_42_4_port, B2 => n17685, C1 => 
                           registers_43_4_port, C2 => n17682, A => n10493, ZN 
                           => n10486);
   U8033 : NAND4_X1 port map( A1 => n10376, A2 => n10377, A3 => n10378, A4 => 
                           n10379, ZN => n10357);
   U8034 : AOI221_X1 port map( B1 => net226999, B2 => n17709, C1 => net226998, 
                           C2 => n17706, A => n10381, ZN => n10378);
   U8035 : AOI221_X1 port map( B1 => net227000, B2 => n17721, C1 => 
                           registers_54_5_port, C2 => n17718, A => n10380, ZN 
                           => n10379);
   U8036 : AOI221_X1 port map( B1 => registers_42_5_port, B2 => n17685, C1 => 
                           registers_43_5_port, C2 => n17682, A => n10383, ZN 
                           => n10376);
   U8037 : NAND4_X1 port map( A1 => n10264, A2 => n10265, A3 => n10266, A4 => 
                           n10267, ZN => n10245);
   U8038 : AOI221_X1 port map( B1 => net227010, B2 => n17709, C1 => net227009, 
                           C2 => n17706, A => n10269, ZN => n10266);
   U8039 : AOI221_X1 port map( B1 => net227011, B2 => n17721, C1 => 
                           registers_54_6_port, C2 => n17718, A => n10268, ZN 
                           => n10267);
   U8040 : AOI221_X1 port map( B1 => registers_42_6_port, B2 => n17685, C1 => 
                           registers_43_6_port, C2 => n17682, A => n10271, ZN 
                           => n10264);
   U8041 : NAND4_X1 port map( A1 => n7628, A2 => n7629, A3 => n7630, A4 => 
                           n7631, ZN => n7609);
   U8042 : AOI221_X1 port map( B1 => net227028, B2 => n17709, C1 => net227027, 
                           C2 => n17706, A => n7633, ZN => n7630);
   U8043 : AOI221_X1 port map( B1 => net227029, B2 => n17721, C1 => 
                           registers_54_7_port, C2 => n17718, A => n7632, ZN =>
                           n7631);
   U8044 : AOI221_X1 port map( B1 => registers_42_7_port, B2 => n17685, C1 => 
                           registers_43_7_port, C2 => n17682, A => n7635, ZN =>
                           n7628);
   U8045 : NAND4_X1 port map( A1 => n7513, A2 => n7514, A3 => n7515, A4 => 
                           n7516, ZN => n7494);
   U8046 : AOI221_X1 port map( B1 => net227046, B2 => n17709, C1 => net227045, 
                           C2 => n17706, A => n7518, ZN => n7515);
   U8047 : AOI221_X1 port map( B1 => net227047, B2 => n17721, C1 => 
                           registers_54_8_port, C2 => n17718, A => n7517, ZN =>
                           n7516);
   U8048 : AOI221_X1 port map( B1 => registers_42_8_port, B2 => n17685, C1 => 
                           registers_43_8_port, C2 => n17682, A => n7520, ZN =>
                           n7513);
   U8049 : NAND4_X1 port map( A1 => n7404, A2 => n7405, A3 => n7406, A4 => 
                           n7407, ZN => n7385);
   U8050 : AOI221_X1 port map( B1 => net227064, B2 => n17709, C1 => net227063, 
                           C2 => n17706, A => n7409, ZN => n7406);
   U8051 : AOI221_X1 port map( B1 => net227065, B2 => n17721, C1 => 
                           registers_54_9_port, C2 => n17718, A => n7408, ZN =>
                           n7407);
   U8052 : AOI221_X1 port map( B1 => registers_42_9_port, B2 => n17685, C1 => 
                           registers_43_9_port, C2 => n17682, A => n7411, ZN =>
                           n7404);
   U8053 : NAND4_X1 port map( A1 => n7295, A2 => n7296, A3 => n7297, A4 => 
                           n7298, ZN => n7276);
   U8054 : AOI221_X1 port map( B1 => net227082, B2 => n17709, C1 => net227081, 
                           C2 => n17706, A => n7300, ZN => n7297);
   U8055 : AOI221_X1 port map( B1 => net227083, B2 => n17721, C1 => 
                           registers_54_10_port, C2 => n17718, A => n7299, ZN 
                           => n7298);
   U8056 : AOI221_X1 port map( B1 => registers_42_10_port, B2 => n17685, C1 => 
                           registers_43_10_port, C2 => n17682, A => n7302, ZN 
                           => n7295);
   U8057 : NAND4_X1 port map( A1 => n7181, A2 => n7182, A3 => n7183, A4 => 
                           n7184, ZN => n7162);
   U8058 : AOI221_X1 port map( B1 => net227100, B2 => n17710, C1 => net227099, 
                           C2 => n17707, A => n7186, ZN => n7183);
   U8059 : AOI221_X1 port map( B1 => net227101, B2 => n17722, C1 => 
                           registers_54_11_port, C2 => n17719, A => n7185, ZN 
                           => n7184);
   U8060 : AOI221_X1 port map( B1 => registers_42_11_port, B2 => n17686, C1 => 
                           registers_43_11_port, C2 => n17683, A => n7188, ZN 
                           => n7181);
   U8061 : NAND4_X1 port map( A1 => n7072, A2 => n7073, A3 => n7074, A4 => 
                           n7075, ZN => n7053);
   U8062 : AOI221_X1 port map( B1 => net227118, B2 => n17710, C1 => net227117, 
                           C2 => n17707, A => n7077, ZN => n7074);
   U8063 : AOI221_X1 port map( B1 => net227119, B2 => n17722, C1 => 
                           registers_54_12_port, C2 => n17719, A => n7076, ZN 
                           => n7075);
   U8064 : AOI221_X1 port map( B1 => registers_42_12_port, B2 => n17686, C1 => 
                           registers_43_12_port, C2 => n17683, A => n7079, ZN 
                           => n7072);
   U8065 : NAND4_X1 port map( A1 => n6963, A2 => n6964, A3 => n6965, A4 => 
                           n6966, ZN => n6944);
   U8066 : AOI221_X1 port map( B1 => net227136, B2 => n17710, C1 => net227135, 
                           C2 => n17707, A => n6968, ZN => n6965);
   U8067 : AOI221_X1 port map( B1 => net227137, B2 => n17722, C1 => 
                           registers_54_13_port, C2 => n17719, A => n6967, ZN 
                           => n6966);
   U8068 : AOI221_X1 port map( B1 => registers_42_13_port, B2 => n17686, C1 => 
                           registers_43_13_port, C2 => n17683, A => n6970, ZN 
                           => n6963);
   U8069 : NAND4_X1 port map( A1 => n6854, A2 => n6855, A3 => n6856, A4 => 
                           n6857, ZN => n6835);
   U8070 : AOI221_X1 port map( B1 => net227154, B2 => n17710, C1 => net227153, 
                           C2 => n17707, A => n6859, ZN => n6856);
   U8071 : AOI221_X1 port map( B1 => net227155, B2 => n17722, C1 => 
                           registers_54_14_port, C2 => n17719, A => n6858, ZN 
                           => n6857);
   U8072 : AOI221_X1 port map( B1 => registers_42_14_port, B2 => n17686, C1 => 
                           registers_43_14_port, C2 => n17683, A => n6861, ZN 
                           => n6854);
   U8073 : NAND4_X1 port map( A1 => n6745, A2 => n6746, A3 => n6747, A4 => 
                           n6748, ZN => n6726);
   U8074 : AOI221_X1 port map( B1 => net227172, B2 => n17710, C1 => net227171, 
                           C2 => n17707, A => n6750, ZN => n6747);
   U8075 : AOI221_X1 port map( B1 => net227173, B2 => n17722, C1 => 
                           registers_54_15_port, C2 => n17719, A => n6749, ZN 
                           => n6748);
   U8076 : AOI221_X1 port map( B1 => registers_42_15_port, B2 => n17686, C1 => 
                           registers_43_15_port, C2 => n17683, A => n6752, ZN 
                           => n6745);
   U8077 : NAND4_X1 port map( A1 => n6602, A2 => n6603, A3 => n6604, A4 => 
                           n6605, ZN => n6563);
   U8078 : AOI221_X1 port map( B1 => net227190, B2 => n17710, C1 => net227189, 
                           C2 => n17707, A => n6607, ZN => n6604);
   U8079 : AOI221_X1 port map( B1 => net227191, B2 => n17722, C1 => 
                           registers_54_16_port, C2 => n17719, A => n6606, ZN 
                           => n6605);
   U8080 : AOI221_X1 port map( B1 => registers_42_16_port, B2 => n17686, C1 => 
                           registers_43_16_port, C2 => n17683, A => n6610, ZN 
                           => n6602);
   U8081 : NAND4_X1 port map( A1 => n6415, A2 => n6416, A3 => n6417, A4 => 
                           n6418, ZN => n6376);
   U8082 : AOI221_X1 port map( B1 => net227208, B2 => n17710, C1 => net227207, 
                           C2 => n17707, A => n6421, ZN => n6417);
   U8083 : AOI221_X1 port map( B1 => net227209, B2 => n17722, C1 => 
                           registers_54_17_port, C2 => n17719, A => n6420, ZN 
                           => n6418);
   U8084 : AOI221_X1 port map( B1 => registers_42_17_port, B2 => n17686, C1 => 
                           registers_43_17_port, C2 => n17683, A => n6425, ZN 
                           => n6415);
   U8085 : NAND4_X1 port map( A1 => n6228, A2 => n6229, A3 => n6231, A4 => 
                           n6232, ZN => n6190);
   U8086 : AOI221_X1 port map( B1 => net227226, B2 => n17710, C1 => net227225, 
                           C2 => n17707, A => n6236, ZN => n6231);
   U8087 : AOI221_X1 port map( B1 => net227227, B2 => n17722, C1 => 
                           registers_54_18_port, C2 => n17719, A => n6234, ZN 
                           => n6232);
   U8088 : AOI221_X1 port map( B1 => registers_42_18_port, B2 => n17686, C1 => 
                           registers_43_18_port, C2 => n17683, A => n6238, ZN 
                           => n6228);
   U8089 : NAND4_X1 port map( A1 => n6042, A2 => n6043, A3 => n6045, A4 => 
                           n6047, ZN => n6005);
   U8090 : AOI221_X1 port map( B1 => net227244, B2 => n17710, C1 => net227243, 
                           C2 => n17707, A => n6049, ZN => n6045);
   U8091 : AOI221_X1 port map( B1 => net227245, B2 => n17722, C1 => 
                           registers_54_19_port, C2 => n17719, A => n6048, ZN 
                           => n6047);
   U8092 : AOI221_X1 port map( B1 => registers_42_19_port, B2 => n17686, C1 => 
                           registers_43_19_port, C2 => n17683, A => n6051, ZN 
                           => n6042);
   U8093 : NAND4_X1 port map( A1 => n5856, A2 => n5858, A3 => n5859, A4 => 
                           n5860, ZN => n5818);
   U8094 : AOI221_X1 port map( B1 => net227262, B2 => n17710, C1 => net227261, 
                           C2 => n17707, A => n5862, ZN => n5859);
   U8095 : AOI221_X1 port map( B1 => net227263, B2 => n17722, C1 => 
                           registers_54_20_port, C2 => n17719, A => n5861, ZN 
                           => n5860);
   U8096 : AOI221_X1 port map( B1 => registers_42_20_port, B2 => n17686, C1 => 
                           registers_43_20_port, C2 => n17683, A => n5866, ZN 
                           => n5856);
   U8097 : NAND4_X1 port map( A1 => n5670, A2 => n5671, A3 => n5672, A4 => 
                           n5673, ZN => n5631);
   U8098 : AOI221_X1 port map( B1 => net227280, B2 => n17710, C1 => net227279, 
                           C2 => n17707, A => n5677, ZN => n5672);
   U8099 : AOI221_X1 port map( B1 => net227281, B2 => n17722, C1 => 
                           registers_54_21_port, C2 => n17719, A => n5674, ZN 
                           => n5673);
   U8100 : AOI221_X1 port map( B1 => registers_42_21_port, B2 => n17686, C1 => 
                           registers_43_21_port, C2 => n17683, A => n5680, ZN 
                           => n5670);
   U8101 : NAND4_X1 port map( A1 => n5483, A2 => n5484, A3 => n5485, A4 => 
                           n5488, ZN => n5446);
   U8102 : AOI221_X1 port map( B1 => net227298, B2 => n17710, C1 => net227297, 
                           C2 => n17707, A => n5491, ZN => n5485);
   U8103 : AOI221_X1 port map( B1 => net227299, B2 => n17722, C1 => 
                           registers_54_22_port, C2 => n17719, A => n5489, ZN 
                           => n5488);
   U8104 : AOI221_X1 port map( B1 => registers_42_22_port, B2 => n17686, C1 => 
                           registers_43_22_port, C2 => n17683, A => n5493, ZN 
                           => n5483);
   U8105 : NAND4_X1 port map( A1 => n14153, A2 => n14154, A3 => n14155, A4 => 
                           n14156, ZN => n14077);
   U8106 : AOI221_X1 port map( B1 => net227460, B2 => n17709, C1 => net227459, 
                           C2 => n17706, A => n14161, ZN => n14155);
   U8107 : AOI221_X1 port map( B1 => net227461, B2 => n17721, C1 => 
                           registers_54_31_port, C2 => n17718, A => n14157, ZN 
                           => n14156);
   U8108 : AOI221_X1 port map( B1 => registers_42_31_port, B2 => n17685, C1 => 
                           registers_43_31_port, C2 => n17682, A => n14175, ZN 
                           => n14153);
   U8109 : NAND4_X1 port map( A1 => n13912, A2 => n13913, A3 => n13914, A4 => 
                           n13915, ZN => n13911);
   U8110 : AOI211_X1 port map( C1 => registers_23_0_port, C2 => n16373, A => 
                           n13934, B => n16412, ZN => n13912);
   U8111 : AOI221_X1 port map( B1 => registers_1_0_port, B2 => n16385, C1 => 
                           registers_19_0_port, C2 => n16382, A => n13930, ZN 
                           => n13913);
   U8112 : AOI221_X1 port map( B1 => registers_16_0_port, B2 => n16397, C1 => 
                           registers_15_0_port, C2 => n16394, A => n13924, ZN 
                           => n13914);
   U8113 : NAND4_X1 port map( A1 => n13865, A2 => n13866, A3 => n13867, A4 => 
                           n13868, ZN => n13864);
   U8114 : AOI211_X1 port map( C1 => registers_23_1_port, C2 => n16373, A => 
                           n13872, B => n16412, ZN => n13865);
   U8115 : AOI221_X1 port map( B1 => registers_1_1_port, B2 => n16385, C1 => 
                           registers_19_1_port, C2 => n16382, A => n13871, ZN 
                           => n13866);
   U8116 : AOI221_X1 port map( B1 => registers_16_1_port, B2 => n16397, C1 => 
                           registers_15_1_port, C2 => n16394, A => n13870, ZN 
                           => n13867);
   U8117 : NAND4_X1 port map( A1 => n13823, A2 => n13824, A3 => n13825, A4 => 
                           n13826, ZN => n13822);
   U8118 : AOI211_X1 port map( C1 => registers_23_2_port, C2 => n16373, A => 
                           n13830, B => n16412, ZN => n13823);
   U8119 : AOI221_X1 port map( B1 => registers_1_2_port, B2 => n16385, C1 => 
                           registers_19_2_port, C2 => n16382, A => n13829, ZN 
                           => n13824);
   U8120 : AOI221_X1 port map( B1 => registers_16_2_port, B2 => n16397, C1 => 
                           registers_15_2_port, C2 => n16394, A => n13828, ZN 
                           => n13825);
   U8121 : NAND4_X1 port map( A1 => n13781, A2 => n13782, A3 => n13783, A4 => 
                           n13784, ZN => n13780);
   U8122 : AOI211_X1 port map( C1 => registers_23_3_port, C2 => n16373, A => 
                           n13788, B => n16412, ZN => n13781);
   U8123 : AOI221_X1 port map( B1 => registers_1_3_port, B2 => n16385, C1 => 
                           registers_19_3_port, C2 => n16382, A => n13787, ZN 
                           => n13782);
   U8124 : AOI221_X1 port map( B1 => registers_16_3_port, B2 => n16397, C1 => 
                           registers_15_3_port, C2 => n16394, A => n13786, ZN 
                           => n13783);
   U8125 : NAND4_X1 port map( A1 => n13739, A2 => n13740, A3 => n13741, A4 => 
                           n13742, ZN => n13738);
   U8126 : AOI211_X1 port map( C1 => registers_23_4_port, C2 => n16373, A => 
                           n13746, B => n16412, ZN => n13739);
   U8127 : AOI221_X1 port map( B1 => registers_1_4_port, B2 => n16385, C1 => 
                           registers_19_4_port, C2 => n16382, A => n13745, ZN 
                           => n13740);
   U8128 : AOI221_X1 port map( B1 => registers_16_4_port, B2 => n16397, C1 => 
                           registers_15_4_port, C2 => n16394, A => n13744, ZN 
                           => n13741);
   U8129 : NAND4_X1 port map( A1 => n13697, A2 => n13698, A3 => n13699, A4 => 
                           n13700, ZN => n13696);
   U8130 : AOI211_X1 port map( C1 => registers_23_5_port, C2 => n16373, A => 
                           n13704, B => n16412, ZN => n13697);
   U8131 : AOI221_X1 port map( B1 => registers_1_5_port, B2 => n16385, C1 => 
                           registers_19_5_port, C2 => n16382, A => n13703, ZN 
                           => n13698);
   U8132 : AOI221_X1 port map( B1 => registers_16_5_port, B2 => n16397, C1 => 
                           registers_15_5_port, C2 => n16394, A => n13702, ZN 
                           => n13699);
   U8133 : NAND4_X1 port map( A1 => n13655, A2 => n13656, A3 => n13657, A4 => 
                           n13658, ZN => n13654);
   U8134 : AOI211_X1 port map( C1 => registers_23_6_port, C2 => n16373, A => 
                           n13662, B => n16412, ZN => n13655);
   U8135 : AOI221_X1 port map( B1 => registers_1_6_port, B2 => n16385, C1 => 
                           registers_19_6_port, C2 => n16382, A => n13661, ZN 
                           => n13656);
   U8136 : AOI221_X1 port map( B1 => registers_16_6_port, B2 => n16397, C1 => 
                           registers_15_6_port, C2 => n16394, A => n13660, ZN 
                           => n13657);
   U8137 : NAND4_X1 port map( A1 => n13613, A2 => n13614, A3 => n13615, A4 => 
                           n13616, ZN => n13612);
   U8138 : AOI211_X1 port map( C1 => registers_23_7_port, C2 => n16373, A => 
                           n13620, B => n16412, ZN => n13613);
   U8139 : AOI221_X1 port map( B1 => registers_1_7_port, B2 => n16385, C1 => 
                           registers_19_7_port, C2 => n16382, A => n13619, ZN 
                           => n13614);
   U8140 : AOI221_X1 port map( B1 => registers_16_7_port, B2 => n16397, C1 => 
                           registers_15_7_port, C2 => n16394, A => n13618, ZN 
                           => n13615);
   U8141 : NAND4_X1 port map( A1 => n13571, A2 => n13572, A3 => n13573, A4 => 
                           n13574, ZN => n13570);
   U8142 : AOI211_X1 port map( C1 => registers_23_8_port, C2 => n16373, A => 
                           n13578, B => n16413, ZN => n13571);
   U8143 : AOI221_X1 port map( B1 => registers_1_8_port, B2 => n16385, C1 => 
                           registers_19_8_port, C2 => n16382, A => n13577, ZN 
                           => n13572);
   U8144 : AOI221_X1 port map( B1 => registers_16_8_port, B2 => n16397, C1 => 
                           registers_15_8_port, C2 => n16394, A => n13576, ZN 
                           => n13573);
   U8145 : NAND4_X1 port map( A1 => n13529, A2 => n13530, A3 => n13531, A4 => 
                           n13532, ZN => n13528);
   U8146 : AOI211_X1 port map( C1 => registers_23_9_port, C2 => n16373, A => 
                           n13536, B => n16413, ZN => n13529);
   U8147 : AOI221_X1 port map( B1 => registers_1_9_port, B2 => n16385, C1 => 
                           registers_19_9_port, C2 => n16382, A => n13535, ZN 
                           => n13530);
   U8148 : AOI221_X1 port map( B1 => registers_16_9_port, B2 => n16397, C1 => 
                           registers_15_9_port, C2 => n16394, A => n13534, ZN 
                           => n13531);
   U8149 : NAND4_X1 port map( A1 => n13487, A2 => n13488, A3 => n13489, A4 => 
                           n13490, ZN => n13486);
   U8150 : AOI211_X1 port map( C1 => registers_23_10_port, C2 => n16373, A => 
                           n13494, B => n16413, ZN => n13487);
   U8151 : AOI221_X1 port map( B1 => registers_1_10_port, B2 => n16385, C1 => 
                           registers_19_10_port, C2 => n16382, A => n13493, ZN 
                           => n13488);
   U8152 : AOI221_X1 port map( B1 => registers_16_10_port, B2 => n16397, C1 => 
                           registers_15_10_port, C2 => n16394, A => n13492, ZN 
                           => n13489);
   U8153 : NAND4_X1 port map( A1 => n13445, A2 => n13446, A3 => n13447, A4 => 
                           n13448, ZN => n13444);
   U8154 : AOI211_X1 port map( C1 => registers_23_11_port, C2 => n16373, A => 
                           n13452, B => n16413, ZN => n13445);
   U8155 : AOI221_X1 port map( B1 => registers_1_11_port, B2 => n16385, C1 => 
                           registers_19_11_port, C2 => n16382, A => n13451, ZN 
                           => n13446);
   U8156 : AOI221_X1 port map( B1 => registers_16_11_port, B2 => n16397, C1 => 
                           registers_15_11_port, C2 => n16394, A => n13450, ZN 
                           => n13447);
   U8157 : NAND4_X1 port map( A1 => n13403, A2 => n13404, A3 => n13405, A4 => 
                           n13406, ZN => n13402);
   U8158 : AOI211_X1 port map( C1 => registers_23_12_port, C2 => n16374, A => 
                           n13410, B => n16413, ZN => n13403);
   U8159 : AOI221_X1 port map( B1 => registers_1_12_port, B2 => n16386, C1 => 
                           registers_19_12_port, C2 => n16383, A => n13409, ZN 
                           => n13404);
   U8160 : AOI221_X1 port map( B1 => registers_16_12_port, B2 => n16398, C1 => 
                           registers_15_12_port, C2 => n16395, A => n13408, ZN 
                           => n13405);
   U8161 : NAND4_X1 port map( A1 => n13361, A2 => n13362, A3 => n13363, A4 => 
                           n13364, ZN => n13360);
   U8162 : AOI211_X1 port map( C1 => registers_23_13_port, C2 => n16374, A => 
                           n13368, B => n16413, ZN => n13361);
   U8163 : AOI221_X1 port map( B1 => registers_1_13_port, B2 => n16386, C1 => 
                           registers_19_13_port, C2 => n16383, A => n13367, ZN 
                           => n13362);
   U8164 : AOI221_X1 port map( B1 => registers_16_13_port, B2 => n16398, C1 => 
                           registers_15_13_port, C2 => n16395, A => n13366, ZN 
                           => n13363);
   U8165 : NAND4_X1 port map( A1 => n13319, A2 => n13320, A3 => n13321, A4 => 
                           n13322, ZN => n13318);
   U8166 : AOI211_X1 port map( C1 => registers_23_14_port, C2 => n16374, A => 
                           n13326, B => n16413, ZN => n13319);
   U8167 : AOI221_X1 port map( B1 => registers_1_14_port, B2 => n16386, C1 => 
                           registers_19_14_port, C2 => n16383, A => n13325, ZN 
                           => n13320);
   U8168 : AOI221_X1 port map( B1 => registers_16_14_port, B2 => n16398, C1 => 
                           registers_15_14_port, C2 => n16395, A => n13324, ZN 
                           => n13321);
   U8169 : NAND4_X1 port map( A1 => n13277, A2 => n13278, A3 => n13279, A4 => 
                           n13280, ZN => n13276);
   U8170 : AOI211_X1 port map( C1 => registers_23_15_port, C2 => n16374, A => 
                           n13284, B => n16413, ZN => n13277);
   U8171 : AOI221_X1 port map( B1 => registers_1_15_port, B2 => n16386, C1 => 
                           registers_19_15_port, C2 => n16383, A => n13283, ZN 
                           => n13278);
   U8172 : AOI221_X1 port map( B1 => registers_16_15_port, B2 => n16398, C1 => 
                           registers_15_15_port, C2 => n16395, A => n13282, ZN 
                           => n13279);
   U8173 : NAND4_X1 port map( A1 => n13151, A2 => n13152, A3 => n13153, A4 => 
                           n13154, ZN => n13150);
   U8174 : AOI211_X1 port map( C1 => registers_23_18_port, C2 => n16374, A => 
                           n13158, B => n16413, ZN => n13151);
   U8175 : AOI221_X1 port map( B1 => registers_1_18_port, B2 => n16386, C1 => 
                           registers_19_18_port, C2 => n16383, A => n13157, ZN 
                           => n13152);
   U8176 : AOI221_X1 port map( B1 => registers_16_18_port, B2 => n16398, C1 => 
                           registers_15_18_port, C2 => n16395, A => n13156, ZN 
                           => n13153);
   U8177 : NAND4_X1 port map( A1 => n12857, A2 => n12858, A3 => n12859, A4 => 
                           n12860, ZN => n12856);
   U8178 : AOI211_X1 port map( C1 => registers_23_25_port, C2 => n16375, A => 
                           n12864, B => n16413, ZN => n12857);
   U8179 : AOI221_X1 port map( B1 => registers_1_25_port, B2 => n16387, C1 => 
                           registers_19_25_port, C2 => n16384, A => n12863, ZN 
                           => n12858);
   U8180 : AOI221_X1 port map( B1 => registers_16_25_port, B2 => n16399, C1 => 
                           registers_15_25_port, C2 => n16396, A => n12862, ZN 
                           => n12859);
   U8181 : NAND4_X1 port map( A1 => n12815, A2 => n12816, A3 => n12817, A4 => 
                           n12818, ZN => n12814);
   U8182 : AOI211_X1 port map( C1 => registers_23_26_port, C2 => n16375, A => 
                           n12822, B => n16413, ZN => n12815);
   U8183 : AOI221_X1 port map( B1 => registers_1_26_port, B2 => n16387, C1 => 
                           registers_19_26_port, C2 => n16384, A => n12821, ZN 
                           => n12816);
   U8184 : AOI221_X1 port map( B1 => registers_16_26_port, B2 => n16399, C1 => 
                           registers_15_26_port, C2 => n16396, A => n12820, ZN 
                           => n12817);
   U8185 : NAND4_X1 port map( A1 => n12773, A2 => n12774, A3 => n12775, A4 => 
                           n12776, ZN => n12772);
   U8186 : AOI211_X1 port map( C1 => registers_23_27_port, C2 => n16375, A => 
                           n12780, B => n16413, ZN => n12773);
   U8187 : AOI221_X1 port map( B1 => registers_1_27_port, B2 => n16387, C1 => 
                           registers_19_27_port, C2 => n16384, A => n12779, ZN 
                           => n12774);
   U8188 : AOI221_X1 port map( B1 => registers_16_27_port, B2 => n16399, C1 => 
                           registers_15_27_port, C2 => n16396, A => n12778, ZN 
                           => n12775);
   U8189 : NAND4_X1 port map( A1 => n12731, A2 => n12732, A3 => n12733, A4 => 
                           n12734, ZN => n12730);
   U8190 : AOI211_X1 port map( C1 => registers_23_28_port, C2 => n16375, A => 
                           n12738, B => n16412, ZN => n12731);
   U8191 : AOI221_X1 port map( B1 => registers_1_28_port, B2 => n16387, C1 => 
                           registers_19_28_port, C2 => n16384, A => n12737, ZN 
                           => n12732);
   U8192 : AOI221_X1 port map( B1 => registers_16_28_port, B2 => n16399, C1 => 
                           registers_15_28_port, C2 => n16396, A => n12736, ZN 
                           => n12733);
   U8193 : NAND4_X1 port map( A1 => n12689, A2 => n12690, A3 => n12691, A4 => 
                           n12692, ZN => n12688);
   U8194 : AOI211_X1 port map( C1 => registers_23_29_port, C2 => n16375, A => 
                           n12696, B => n16412, ZN => n12689);
   U8195 : AOI221_X1 port map( B1 => registers_1_29_port, B2 => n16387, C1 => 
                           registers_19_29_port, C2 => n16384, A => n12695, ZN 
                           => n12690);
   U8196 : AOI221_X1 port map( B1 => registers_16_29_port, B2 => n16399, C1 => 
                           registers_15_29_port, C2 => n16396, A => n12694, ZN 
                           => n12691);
   U8197 : NAND4_X1 port map( A1 => n12645, A2 => n12646, A3 => n12647, A4 => 
                           n12648, ZN => n12644);
   U8198 : AOI211_X1 port map( C1 => registers_23_30_port, C2 => n16375, A => 
                           n12653, B => n16412, ZN => n12645);
   U8199 : AOI221_X1 port map( B1 => registers_1_30_port, B2 => n16387, C1 => 
                           registers_19_30_port, C2 => n16384, A => n12651, ZN 
                           => n12646);
   U8200 : AOI221_X1 port map( B1 => registers_16_30_port, B2 => n16399, C1 => 
                           registers_15_30_port, C2 => n16396, A => n12650, ZN 
                           => n12647);
   U8201 : NAND4_X1 port map( A1 => n12533, A2 => n12534, A3 => n12535, A4 => 
                           n12536, ZN => n12532);
   U8202 : AOI211_X1 port map( C1 => registers_23_31_port, C2 => n16375, A => 
                           n12554, B => n16412, ZN => n12533);
   U8203 : AOI221_X1 port map( B1 => registers_1_31_port, B2 => n16387, C1 => 
                           registers_19_31_port, C2 => n16384, A => n12549, ZN 
                           => n12534);
   U8204 : AOI221_X1 port map( B1 => registers_16_31_port, B2 => n16399, C1 => 
                           registers_15_31_port, C2 => n16396, A => n12544, ZN 
                           => n12535);
   U8205 : NAND4_X1 port map( A1 => n12431, A2 => n12432, A3 => n12433, A4 => 
                           n12434, ZN => n12430);
   U8206 : AOI221_X1 port map( B1 => registers_16_0_port, B2 => n16649, C1 => 
                           registers_19_0_port, C2 => n16646, A => n12442, ZN 
                           => n12433);
   U8207 : AOI211_X1 port map( C1 => registers_23_0_port, C2 => n16625, A => 
                           n12453, B => n16664, ZN => n12431);
   U8208 : AOI221_X1 port map( B1 => registers_1_0_port, B2 => n16637, C1 => 
                           registers_22_0_port, C2 => n16634, A => n12448, ZN 
                           => n12432);
   U8209 : NAND4_X1 port map( A1 => n12269, A2 => n12270, A3 => n12271, A4 => 
                           n12272, ZN => n12268);
   U8210 : AOI221_X1 port map( B1 => registers_16_1_port, B2 => n16649, C1 => 
                           registers_19_1_port, C2 => n16646, A => n12274, ZN 
                           => n12271);
   U8211 : AOI211_X1 port map( C1 => registers_23_1_port, C2 => n16625, A => 
                           n12276, B => n16664, ZN => n12269);
   U8212 : AOI221_X1 port map( B1 => registers_1_1_port, B2 => n16637, C1 => 
                           registers_22_1_port, C2 => n16634, A => n12275, ZN 
                           => n12270);
   U8213 : NAND4_X1 port map( A1 => n12116, A2 => n12117, A3 => n12118, A4 => 
                           n12119, ZN => n12115);
   U8214 : AOI221_X1 port map( B1 => registers_16_2_port, B2 => n16649, C1 => 
                           registers_19_2_port, C2 => n16646, A => n12121, ZN 
                           => n12118);
   U8215 : AOI211_X1 port map( C1 => registers_23_2_port, C2 => n16625, A => 
                           n12123, B => n16664, ZN => n12116);
   U8216 : AOI221_X1 port map( B1 => registers_1_2_port, B2 => n16637, C1 => 
                           registers_22_2_port, C2 => n16634, A => n12122, ZN 
                           => n12117);
   U8217 : NAND4_X1 port map( A1 => n11963, A2 => n11964, A3 => n11965, A4 => 
                           n11966, ZN => n11962);
   U8218 : AOI221_X1 port map( B1 => registers_16_3_port, B2 => n16649, C1 => 
                           registers_19_3_port, C2 => n16646, A => n11968, ZN 
                           => n11965);
   U8219 : AOI211_X1 port map( C1 => registers_23_3_port, C2 => n16625, A => 
                           n11970, B => n16664, ZN => n11963);
   U8220 : AOI221_X1 port map( B1 => registers_1_3_port, B2 => n16637, C1 => 
                           registers_22_3_port, C2 => n16634, A => n11969, ZN 
                           => n11964);
   U8221 : NAND4_X1 port map( A1 => n11810, A2 => n11811, A3 => n11812, A4 => 
                           n11813, ZN => n11809);
   U8222 : AOI221_X1 port map( B1 => registers_16_4_port, B2 => n16649, C1 => 
                           registers_19_4_port, C2 => n16646, A => n11815, ZN 
                           => n11812);
   U8223 : AOI211_X1 port map( C1 => registers_23_4_port, C2 => n16625, A => 
                           n11817, B => n16664, ZN => n11810);
   U8224 : AOI221_X1 port map( B1 => registers_1_4_port, B2 => n16637, C1 => 
                           registers_22_4_port, C2 => n16634, A => n11816, ZN 
                           => n11811);
   U8225 : NAND4_X1 port map( A1 => n11767, A2 => n11768, A3 => n11769, A4 => 
                           n11770, ZN => n11766);
   U8226 : AOI221_X1 port map( B1 => registers_16_5_port, B2 => n16649, C1 => 
                           registers_19_5_port, C2 => n16646, A => n11772, ZN 
                           => n11769);
   U8227 : AOI211_X1 port map( C1 => registers_23_5_port, C2 => n16625, A => 
                           n11774, B => n16664, ZN => n11767);
   U8228 : AOI221_X1 port map( B1 => registers_1_5_port, B2 => n16637, C1 => 
                           registers_22_5_port, C2 => n16634, A => n11773, ZN 
                           => n11768);
   U8229 : NAND4_X1 port map( A1 => n11724, A2 => n11725, A3 => n11726, A4 => 
                           n11727, ZN => n11723);
   U8230 : AOI221_X1 port map( B1 => registers_16_6_port, B2 => n16649, C1 => 
                           registers_19_6_port, C2 => n16646, A => n11729, ZN 
                           => n11726);
   U8231 : AOI211_X1 port map( C1 => registers_23_6_port, C2 => n16625, A => 
                           n11731, B => n16664, ZN => n11724);
   U8232 : AOI221_X1 port map( B1 => registers_1_6_port, B2 => n16637, C1 => 
                           registers_22_6_port, C2 => n16634, A => n11730, ZN 
                           => n11725);
   U8233 : NAND4_X1 port map( A1 => n11681, A2 => n11682, A3 => n11683, A4 => 
                           n11684, ZN => n11680);
   U8234 : AOI221_X1 port map( B1 => registers_16_7_port, B2 => n16649, C1 => 
                           registers_19_7_port, C2 => n16646, A => n11686, ZN 
                           => n11683);
   U8235 : AOI211_X1 port map( C1 => registers_23_7_port, C2 => n16625, A => 
                           n11688, B => n16664, ZN => n11681);
   U8236 : AOI221_X1 port map( B1 => registers_1_7_port, B2 => n16637, C1 => 
                           registers_22_7_port, C2 => n16634, A => n11687, ZN 
                           => n11682);
   U8237 : NAND4_X1 port map( A1 => n11638, A2 => n11639, A3 => n11640, A4 => 
                           n11641, ZN => n11637);
   U8238 : AOI221_X1 port map( B1 => registers_16_8_port, B2 => n16649, C1 => 
                           registers_19_8_port, C2 => n16646, A => n11643, ZN 
                           => n11640);
   U8239 : AOI211_X1 port map( C1 => registers_23_8_port, C2 => n16625, A => 
                           n11645, B => n16665, ZN => n11638);
   U8240 : AOI221_X1 port map( B1 => registers_1_8_port, B2 => n16637, C1 => 
                           registers_22_8_port, C2 => n16634, A => n11644, ZN 
                           => n11639);
   U8241 : NAND4_X1 port map( A1 => n11595, A2 => n11596, A3 => n11597, A4 => 
                           n11598, ZN => n11594);
   U8242 : AOI221_X1 port map( B1 => registers_16_9_port, B2 => n16649, C1 => 
                           registers_19_9_port, C2 => n16646, A => n11600, ZN 
                           => n11597);
   U8243 : AOI211_X1 port map( C1 => registers_23_9_port, C2 => n16625, A => 
                           n11602, B => n16665, ZN => n11595);
   U8244 : AOI221_X1 port map( B1 => registers_1_9_port, B2 => n16637, C1 => 
                           registers_22_9_port, C2 => n16634, A => n11601, ZN 
                           => n11596);
   U8245 : NAND4_X1 port map( A1 => n11552, A2 => n11553, A3 => n11554, A4 => 
                           n11555, ZN => n11551);
   U8246 : AOI221_X1 port map( B1 => registers_16_10_port, B2 => n16649, C1 => 
                           registers_19_10_port, C2 => n16646, A => n11557, ZN 
                           => n11554);
   U8247 : AOI211_X1 port map( C1 => registers_23_10_port, C2 => n16625, A => 
                           n11559, B => n16665, ZN => n11552);
   U8248 : AOI221_X1 port map( B1 => registers_1_10_port, B2 => n16637, C1 => 
                           registers_22_10_port, C2 => n16634, A => n11558, ZN 
                           => n11553);
   U8249 : NAND4_X1 port map( A1 => n11509, A2 => n11510, A3 => n11511, A4 => 
                           n11512, ZN => n11508);
   U8250 : AOI221_X1 port map( B1 => registers_16_11_port, B2 => n16649, C1 => 
                           registers_19_11_port, C2 => n16646, A => n11514, ZN 
                           => n11511);
   U8251 : AOI211_X1 port map( C1 => registers_23_11_port, C2 => n16625, A => 
                           n11516, B => n16665, ZN => n11509);
   U8252 : AOI221_X1 port map( B1 => registers_1_11_port, B2 => n16637, C1 => 
                           registers_22_11_port, C2 => n16634, A => n11515, ZN 
                           => n11510);
   U8253 : NAND4_X1 port map( A1 => n11466, A2 => n11467, A3 => n11468, A4 => 
                           n11469, ZN => n11465);
   U8254 : AOI221_X1 port map( B1 => registers_16_12_port, B2 => n16650, C1 => 
                           registers_19_12_port, C2 => n16647, A => n11471, ZN 
                           => n11468);
   U8255 : AOI211_X1 port map( C1 => registers_23_12_port, C2 => n16626, A => 
                           n11473, B => n16665, ZN => n11466);
   U8256 : AOI221_X1 port map( B1 => registers_1_12_port, B2 => n16638, C1 => 
                           registers_22_12_port, C2 => n16635, A => n11472, ZN 
                           => n11467);
   U8257 : NAND4_X1 port map( A1 => n11422, A2 => n11423, A3 => n11424, A4 => 
                           n11425, ZN => n11421);
   U8258 : AOI221_X1 port map( B1 => registers_16_13_port, B2 => n16650, C1 => 
                           registers_19_13_port, C2 => n16647, A => n11427, ZN 
                           => n11424);
   U8259 : AOI211_X1 port map( C1 => registers_23_13_port, C2 => n16626, A => 
                           n11429, B => n16665, ZN => n11422);
   U8260 : AOI221_X1 port map( B1 => registers_1_13_port, B2 => n16638, C1 => 
                           registers_22_13_port, C2 => n16635, A => n11428, ZN 
                           => n11423);
   U8261 : NAND4_X1 port map( A1 => n11379, A2 => n11380, A3 => n11381, A4 => 
                           n11382, ZN => n11378);
   U8262 : AOI221_X1 port map( B1 => registers_16_14_port, B2 => n16650, C1 => 
                           registers_19_14_port, C2 => n16647, A => n11384, ZN 
                           => n11381);
   U8263 : AOI211_X1 port map( C1 => registers_23_14_port, C2 => n16626, A => 
                           n11386, B => n16665, ZN => n11379);
   U8264 : AOI221_X1 port map( B1 => registers_1_14_port, B2 => n16638, C1 => 
                           registers_22_14_port, C2 => n16635, A => n11385, ZN 
                           => n11380);
   U8265 : NAND4_X1 port map( A1 => n11336, A2 => n11337, A3 => n11338, A4 => 
                           n11339, ZN => n11335);
   U8266 : AOI221_X1 port map( B1 => registers_16_15_port, B2 => n16650, C1 => 
                           registers_19_15_port, C2 => n16647, A => n11341, ZN 
                           => n11338);
   U8267 : AOI211_X1 port map( C1 => registers_23_15_port, C2 => n16626, A => 
                           n11343, B => n16665, ZN => n11336);
   U8268 : AOI221_X1 port map( B1 => registers_1_15_port, B2 => n16638, C1 => 
                           registers_22_15_port, C2 => n16635, A => n11342, ZN 
                           => n11337);
   U8269 : NAND4_X1 port map( A1 => n11207, A2 => n11208, A3 => n11209, A4 => 
                           n11210, ZN => n11206);
   U8270 : AOI221_X1 port map( B1 => registers_16_18_port, B2 => n16650, C1 => 
                           registers_19_18_port, C2 => n16647, A => n11212, ZN 
                           => n11209);
   U8271 : AOI211_X1 port map( C1 => registers_23_18_port, C2 => n16626, A => 
                           n11214, B => n16665, ZN => n11207);
   U8272 : AOI221_X1 port map( B1 => registers_1_18_port, B2 => n16638, C1 => 
                           registers_22_18_port, C2 => n16635, A => n11213, ZN 
                           => n11208);
   U8273 : NAND4_X1 port map( A1 => n10906, A2 => n10907, A3 => n10908, A4 => 
                           n10909, ZN => n10905);
   U8274 : AOI221_X1 port map( B1 => registers_16_25_port, B2 => n16651, C1 => 
                           registers_19_25_port, C2 => n16648, A => n10911, ZN 
                           => n10908);
   U8275 : AOI211_X1 port map( C1 => registers_23_25_port, C2 => n16627, A => 
                           n10913, B => n16665, ZN => n10906);
   U8276 : AOI221_X1 port map( B1 => registers_1_25_port, B2 => n16639, C1 => 
                           registers_22_25_port, C2 => n16636, A => n10912, ZN 
                           => n10907);
   U8277 : NAND4_X1 port map( A1 => n10863, A2 => n10864, A3 => n10865, A4 => 
                           n10866, ZN => n10862);
   U8278 : AOI221_X1 port map( B1 => registers_16_26_port, B2 => n16651, C1 => 
                           registers_19_26_port, C2 => n16648, A => n10868, ZN 
                           => n10865);
   U8279 : AOI211_X1 port map( C1 => registers_23_26_port, C2 => n16627, A => 
                           n10870, B => n16665, ZN => n10863);
   U8280 : AOI221_X1 port map( B1 => registers_1_26_port, B2 => n16639, C1 => 
                           registers_22_26_port, C2 => n16636, A => n10869, ZN 
                           => n10864);
   U8281 : NAND4_X1 port map( A1 => n10820, A2 => n10821, A3 => n10822, A4 => 
                           n10823, ZN => n10819);
   U8282 : AOI221_X1 port map( B1 => registers_16_27_port, B2 => n16651, C1 => 
                           registers_19_27_port, C2 => n16648, A => n10825, ZN 
                           => n10822);
   U8283 : AOI211_X1 port map( C1 => registers_23_27_port, C2 => n16627, A => 
                           n10827, B => n16665, ZN => n10820);
   U8284 : AOI221_X1 port map( B1 => registers_1_27_port, B2 => n16639, C1 => 
                           registers_22_27_port, C2 => n16636, A => n10826, ZN 
                           => n10821);
   U8285 : NAND4_X1 port map( A1 => n10777, A2 => n10778, A3 => n10779, A4 => 
                           n10780, ZN => n10776);
   U8286 : AOI221_X1 port map( B1 => registers_16_28_port, B2 => n16651, C1 => 
                           registers_19_28_port, C2 => n16648, A => n10782, ZN 
                           => n10779);
   U8287 : AOI211_X1 port map( C1 => registers_23_28_port, C2 => n16627, A => 
                           n10784, B => n16664, ZN => n10777);
   U8288 : AOI221_X1 port map( B1 => registers_1_28_port, B2 => n16639, C1 => 
                           registers_22_28_port, C2 => n16636, A => n10783, ZN 
                           => n10778);
   U8289 : NAND4_X1 port map( A1 => n10734, A2 => n10735, A3 => n10736, A4 => 
                           n10737, ZN => n10733);
   U8290 : AOI221_X1 port map( B1 => registers_16_29_port, B2 => n16651, C1 => 
                           registers_19_29_port, C2 => n16648, A => n10739, ZN 
                           => n10736);
   U8291 : AOI211_X1 port map( C1 => registers_23_29_port, C2 => n16627, A => 
                           n10741, B => n16664, ZN => n10734);
   U8292 : AOI221_X1 port map( B1 => registers_1_29_port, B2 => n16639, C1 => 
                           registers_22_29_port, C2 => n16636, A => n10740, ZN 
                           => n10735);
   U8293 : NAND4_X1 port map( A1 => n10675, A2 => n10676, A3 => n10677, A4 => 
                           n10678, ZN => n10674);
   U8294 : AOI221_X1 port map( B1 => registers_16_30_port, B2 => n16651, C1 => 
                           registers_19_30_port, C2 => n16648, A => n10682, ZN 
                           => n10677);
   U8295 : AOI211_X1 port map( C1 => registers_23_30_port, C2 => n16627, A => 
                           n10685, B => n16664, ZN => n10675);
   U8296 : AOI221_X1 port map( B1 => registers_1_30_port, B2 => n16639, C1 => 
                           registers_22_30_port, C2 => n16636, A => n10683, ZN 
                           => n10676);
   U8297 : NAND4_X1 port map( A1 => n10531, A2 => n10532, A3 => n10533, A4 => 
                           n10534, ZN => n10530);
   U8298 : AOI221_X1 port map( B1 => registers_16_31_port, B2 => n16651, C1 => 
                           registers_19_31_port, C2 => n16648, A => n10544, ZN 
                           => n10533);
   U8299 : AOI211_X1 port map( C1 => registers_23_31_port, C2 => n16627, A => 
                           n10557, B => n16664, ZN => n10531);
   U8300 : AOI221_X1 port map( B1 => registers_1_31_port, B2 => n16639, C1 => 
                           registers_22_31_port, C2 => n16636, A => n10551, ZN 
                           => n10532);
   U8301 : NAND4_X1 port map( A1 => n13235, A2 => n13236, A3 => n13237, A4 => 
                           n13238, ZN => n13234);
   U8302 : AOI211_X1 port map( C1 => registers_23_16_port, C2 => n16374, A => 
                           n13242, B => n16414, ZN => n13235);
   U8303 : AOI221_X1 port map( B1 => registers_1_16_port, B2 => n16386, C1 => 
                           registers_19_16_port, C2 => n16383, A => n13241, ZN 
                           => n13236);
   U8304 : AOI221_X1 port map( B1 => registers_16_16_port, B2 => n16398, C1 => 
                           registers_15_16_port, C2 => n16395, A => n13240, ZN 
                           => n13237);
   U8305 : NAND4_X1 port map( A1 => n13193, A2 => n13194, A3 => n13195, A4 => 
                           n13196, ZN => n13192);
   U8306 : AOI211_X1 port map( C1 => registers_23_17_port, C2 => n16374, A => 
                           n13200, B => n16414, ZN => n13193);
   U8307 : AOI221_X1 port map( B1 => registers_1_17_port, B2 => n16386, C1 => 
                           registers_19_17_port, C2 => n16383, A => n13199, ZN 
                           => n13194);
   U8308 : AOI221_X1 port map( B1 => registers_16_17_port, B2 => n16398, C1 => 
                           registers_15_17_port, C2 => n16395, A => n13198, ZN 
                           => n13195);
   U8309 : NAND4_X1 port map( A1 => n13109, A2 => n13110, A3 => n13111, A4 => 
                           n13112, ZN => n13108);
   U8310 : AOI211_X1 port map( C1 => registers_23_19_port, C2 => n16374, A => 
                           n13116, B => n16414, ZN => n13109);
   U8311 : AOI221_X1 port map( B1 => registers_1_19_port, B2 => n16386, C1 => 
                           registers_19_19_port, C2 => n16383, A => n13115, ZN 
                           => n13110);
   U8312 : AOI221_X1 port map( B1 => registers_16_19_port, B2 => n16398, C1 => 
                           registers_15_19_port, C2 => n16395, A => n13114, ZN 
                           => n13111);
   U8313 : NAND4_X1 port map( A1 => n13067, A2 => n13068, A3 => n13069, A4 => 
                           n13070, ZN => n13066);
   U8314 : AOI211_X1 port map( C1 => registers_23_20_port, C2 => n16374, A => 
                           n13074, B => n16414, ZN => n13067);
   U8315 : AOI221_X1 port map( B1 => registers_1_20_port, B2 => n16386, C1 => 
                           registers_19_20_port, C2 => n16383, A => n13073, ZN 
                           => n13068);
   U8316 : AOI221_X1 port map( B1 => registers_16_20_port, B2 => n16398, C1 => 
                           registers_15_20_port, C2 => n16395, A => n13072, ZN 
                           => n13069);
   U8317 : NAND4_X1 port map( A1 => n13025, A2 => n13026, A3 => n13027, A4 => 
                           n13028, ZN => n13024);
   U8318 : AOI211_X1 port map( C1 => registers_23_21_port, C2 => n16374, A => 
                           n13032, B => n16414, ZN => n13025);
   U8319 : AOI221_X1 port map( B1 => registers_1_21_port, B2 => n16386, C1 => 
                           registers_19_21_port, C2 => n16383, A => n13031, ZN 
                           => n13026);
   U8320 : AOI221_X1 port map( B1 => registers_16_21_port, B2 => n16398, C1 => 
                           registers_15_21_port, C2 => n16395, A => n13030, ZN 
                           => n13027);
   U8321 : NAND4_X1 port map( A1 => n12983, A2 => n12984, A3 => n12985, A4 => 
                           n12986, ZN => n12982);
   U8322 : AOI211_X1 port map( C1 => registers_23_22_port, C2 => n16374, A => 
                           n12990, B => n16414, ZN => n12983);
   U8323 : AOI221_X1 port map( B1 => registers_1_22_port, B2 => n16386, C1 => 
                           registers_19_22_port, C2 => n16383, A => n12989, ZN 
                           => n12984);
   U8324 : AOI221_X1 port map( B1 => registers_16_22_port, B2 => n16398, C1 => 
                           registers_15_22_port, C2 => n16395, A => n12988, ZN 
                           => n12985);
   U8325 : NAND4_X1 port map( A1 => n12941, A2 => n12942, A3 => n12943, A4 => 
                           n12944, ZN => n12940);
   U8326 : AOI211_X1 port map( C1 => registers_23_23_port, C2 => n16374, A => 
                           n12948, B => n16414, ZN => n12941);
   U8327 : AOI221_X1 port map( B1 => registers_1_23_port, B2 => n16386, C1 => 
                           registers_19_23_port, C2 => n16383, A => n12947, ZN 
                           => n12942);
   U8328 : AOI221_X1 port map( B1 => registers_16_23_port, B2 => n16398, C1 => 
                           registers_15_23_port, C2 => n16395, A => n12946, ZN 
                           => n12943);
   U8329 : NAND4_X1 port map( A1 => n12899, A2 => n12900, A3 => n12901, A4 => 
                           n12902, ZN => n12898);
   U8330 : AOI211_X1 port map( C1 => registers_23_24_port, C2 => n16375, A => 
                           n12906, B => n16414, ZN => n12899);
   U8331 : AOI221_X1 port map( B1 => registers_1_24_port, B2 => n16387, C1 => 
                           registers_19_24_port, C2 => n16384, A => n12905, ZN 
                           => n12900);
   U8332 : AOI221_X1 port map( B1 => registers_16_24_port, B2 => n16399, C1 => 
                           registers_15_24_port, C2 => n16396, A => n12904, ZN 
                           => n12901);
   U8333 : NAND4_X1 port map( A1 => n11293, A2 => n11294, A3 => n11295, A4 => 
                           n11296, ZN => n11292);
   U8334 : AOI221_X1 port map( B1 => registers_16_16_port, B2 => n16650, C1 => 
                           registers_19_16_port, C2 => n16647, A => n11298, ZN 
                           => n11295);
   U8335 : AOI211_X1 port map( C1 => registers_23_16_port, C2 => n16626, A => 
                           n11300, B => n16666, ZN => n11293);
   U8336 : AOI221_X1 port map( B1 => registers_1_16_port, B2 => n16638, C1 => 
                           registers_22_16_port, C2 => n16635, A => n11299, ZN 
                           => n11294);
   U8337 : NAND4_X1 port map( A1 => n11250, A2 => n11251, A3 => n11252, A4 => 
                           n11253, ZN => n11249);
   U8338 : AOI221_X1 port map( B1 => registers_16_17_port, B2 => n16650, C1 => 
                           registers_19_17_port, C2 => n16647, A => n11255, ZN 
                           => n11252);
   U8339 : AOI211_X1 port map( C1 => registers_23_17_port, C2 => n16626, A => 
                           n11257, B => n16666, ZN => n11250);
   U8340 : AOI221_X1 port map( B1 => registers_1_17_port, B2 => n16638, C1 => 
                           registers_22_17_port, C2 => n16635, A => n11256, ZN 
                           => n11251);
   U8341 : NAND4_X1 port map( A1 => n11164, A2 => n11165, A3 => n11166, A4 => 
                           n11167, ZN => n11163);
   U8342 : AOI221_X1 port map( B1 => registers_16_19_port, B2 => n16650, C1 => 
                           registers_19_19_port, C2 => n16647, A => n11169, ZN 
                           => n11166);
   U8343 : AOI211_X1 port map( C1 => registers_23_19_port, C2 => n16626, A => 
                           n11171, B => n16666, ZN => n11164);
   U8344 : AOI221_X1 port map( B1 => registers_1_19_port, B2 => n16638, C1 => 
                           registers_22_19_port, C2 => n16635, A => n11170, ZN 
                           => n11165);
   U8345 : NAND4_X1 port map( A1 => n11121, A2 => n11122, A3 => n11123, A4 => 
                           n11124, ZN => n11120);
   U8346 : AOI221_X1 port map( B1 => registers_16_20_port, B2 => n16650, C1 => 
                           registers_19_20_port, C2 => n16647, A => n11126, ZN 
                           => n11123);
   U8347 : AOI211_X1 port map( C1 => registers_23_20_port, C2 => n16626, A => 
                           n11128, B => n16666, ZN => n11121);
   U8348 : AOI221_X1 port map( B1 => registers_1_20_port, B2 => n16638, C1 => 
                           registers_22_20_port, C2 => n16635, A => n11127, ZN 
                           => n11122);
   U8349 : NAND4_X1 port map( A1 => n11078, A2 => n11079, A3 => n11080, A4 => 
                           n11081, ZN => n11077);
   U8350 : AOI221_X1 port map( B1 => registers_16_21_port, B2 => n16650, C1 => 
                           registers_19_21_port, C2 => n16647, A => n11083, ZN 
                           => n11080);
   U8351 : AOI211_X1 port map( C1 => registers_23_21_port, C2 => n16626, A => 
                           n11085, B => n16666, ZN => n11078);
   U8352 : AOI221_X1 port map( B1 => registers_1_21_port, B2 => n16638, C1 => 
                           registers_22_21_port, C2 => n16635, A => n11084, ZN 
                           => n11079);
   U8353 : NAND4_X1 port map( A1 => n11035, A2 => n11036, A3 => n11037, A4 => 
                           n11038, ZN => n11034);
   U8354 : AOI221_X1 port map( B1 => registers_16_22_port, B2 => n16650, C1 => 
                           registers_19_22_port, C2 => n16647, A => n11040, ZN 
                           => n11037);
   U8355 : AOI211_X1 port map( C1 => registers_23_22_port, C2 => n16626, A => 
                           n11042, B => n16666, ZN => n11035);
   U8356 : AOI221_X1 port map( B1 => registers_1_22_port, B2 => n16638, C1 => 
                           registers_22_22_port, C2 => n16635, A => n11041, ZN 
                           => n11036);
   U8357 : NAND4_X1 port map( A1 => n10992, A2 => n10993, A3 => n10994, A4 => 
                           n10995, ZN => n10991);
   U8358 : AOI221_X1 port map( B1 => registers_16_23_port, B2 => n16650, C1 => 
                           registers_19_23_port, C2 => n16647, A => n10997, ZN 
                           => n10994);
   U8359 : AOI211_X1 port map( C1 => registers_23_23_port, C2 => n16626, A => 
                           n10999, B => n16666, ZN => n10992);
   U8360 : AOI221_X1 port map( B1 => registers_1_23_port, B2 => n16638, C1 => 
                           registers_22_23_port, C2 => n16635, A => n10998, ZN 
                           => n10993);
   U8361 : NAND4_X1 port map( A1 => n10949, A2 => n10950, A3 => n10951, A4 => 
                           n10952, ZN => n10948);
   U8362 : AOI221_X1 port map( B1 => registers_16_24_port, B2 => n16651, C1 => 
                           registers_19_24_port, C2 => n16648, A => n10954, ZN 
                           => n10951);
   U8363 : AOI211_X1 port map( C1 => registers_23_24_port, C2 => n16627, A => 
                           n10956, B => n16666, ZN => n10949);
   U8364 : AOI221_X1 port map( B1 => registers_1_24_port, B2 => n16639, C1 => 
                           registers_22_24_port, C2 => n16636, A => n10955, ZN 
                           => n10950);
   U8365 : NAND2_X1 port map( A1 => n14016, A2 => call, ZN => n14159);
   U8366 : NAND2_X1 port map( A1 => n10190, A2 => N9909, ZN => n14144);
   U8367 : INV_X1 port map( A => add_rd2(2), ZN => n13984);
   U8368 : INV_X1 port map( A => add_wr(0), ZN => n14229);
   U8369 : INV_X1 port map( A => add_rd1(2), ZN => n12503);
   U8370 : AND2_X1 port map( A1 => n13987, A2 => add_rd2(0), ZN => n13901);
   U8371 : AND2_X1 port map( A1 => n12506, A2 => add_rd1(0), ZN => n12420);
   U8372 : NAND2_X1 port map( A1 => n7592, A2 => n14265, ZN => n14247);
   U8373 : OR2_X1 port map( A1 => add_wr(0), A2 => add_wr(1), ZN => n14213);
   U8374 : NOR2_X1 port map( A1 => n10189, A2 => n14004, ZN => n10179);
   U8375 : NOR2_X1 port map( A1 => n10187, A2 => n14004, ZN => n10175);
   U8376 : NOR2_X1 port map( A1 => n7587, A2 => n14229, ZN => 
                           add_73_carry_1_port);
   U8377 : NOR2_X1 port map( A1 => n10190, A2 => n14004, ZN => n10180);
   U8378 : OAI21_X1 port map( B1 => n5522, B2 => n18049, A => n13998, ZN => 
                           n10183);
   U8379 : NOR2_X1 port map( A1 => n10188, A2 => n14004, ZN => n10177);
   U8380 : AOI22_X1 port map( A1 => net226855, A2 => n16466, B1 => 
                           registers_68_1_port, B2 => n16463, ZN => n12259);
   U8381 : AOI221_X1 port map( B1 => net226854, B2 => n16687, C1 => net226853, 
                           C2 => n16682, A => n12262, ZN => n12261);
   U8382 : AOI221_X1 port map( B1 => net226856, B2 => n16675, C1 => net226865, 
                           C2 => n16670, A => n12263, ZN => n12260);
   U8383 : AOI22_X1 port map( A1 => net226876, A2 => n16466, B1 => 
                           registers_68_2_port, B2 => n16463, ZN => n12106);
   U8384 : AOI221_X1 port map( B1 => net226874, B2 => n16687, C1 => net226873, 
                           C2 => n16682, A => n12109, ZN => n12108);
   U8385 : AOI221_X1 port map( B1 => net226877, B2 => n16675, C1 => net226875, 
                           C2 => n16670, A => n12110, ZN => n12107);
   U8386 : AOI22_X1 port map( A1 => net226896, A2 => n16466, B1 => 
                           registers_68_3_port, B2 => n16463, ZN => n11953);
   U8387 : AOI221_X1 port map( B1 => net226894, B2 => n16687, C1 => net226893, 
                           C2 => n16682, A => n11956, ZN => n11955);
   U8388 : AOI221_X1 port map( B1 => net226897, B2 => n16675, C1 => net226895, 
                           C2 => n16670, A => n11957, ZN => n11954);
   U8389 : AOI22_X1 port map( A1 => n16214, A2 => net226843, B1 => n16213, B2 
                           => registers_68_0_port, ZN => n13897);
   U8390 : AOI221_X1 port map( B1 => n16433, B2 => net226842, C1 => n16430, C2 
                           => net226833, A => n13900, ZN => n13899);
   U8391 : AOI221_X1 port map( B1 => n16421, B2 => net226835, C1 => n16418, C2 
                           => net226834, A => n13906, ZN => n13898);
   U8392 : AOI22_X1 port map( A1 => n16214, A2 => net226855, B1 => n16213, B2 
                           => registers_68_1_port, ZN => n13855);
   U8393 : AOI221_X1 port map( B1 => n16433, B2 => net226854, C1 => n16430, C2 
                           => net226853, A => n13858, ZN => n13857);
   U8394 : AOI221_X1 port map( B1 => n16421, B2 => net226856, C1 => n16418, C2 
                           => net226865, A => n13859, ZN => n13856);
   U8395 : AOI22_X1 port map( A1 => n16214, A2 => net226876, B1 => n16213, B2 
                           => registers_68_2_port, ZN => n13813);
   U8396 : AOI221_X1 port map( B1 => n16433, B2 => net226874, C1 => n16430, C2 
                           => net226873, A => n13816, ZN => n13815);
   U8397 : AOI221_X1 port map( B1 => n16421, B2 => net226877, C1 => n16418, C2 
                           => net226875, A => n13817, ZN => n13814);
   U8398 : AOI22_X1 port map( A1 => n16214, A2 => net226896, B1 => n16213, B2 
                           => registers_68_3_port, ZN => n13771);
   U8399 : AOI221_X1 port map( B1 => n16433, B2 => net226894, C1 => n16430, C2 
                           => net226893, A => n13774, ZN => n13773);
   U8400 : AOI221_X1 port map( B1 => n16421, B2 => net226897, C1 => n16418, C2 
                           => net226895, A => n13775, ZN => n13772);
   U8401 : AOI22_X1 port map( A1 => n16214, A2 => net226970, B1 => n16213, B2 
                           => registers_68_4_port, ZN => n13729);
   U8402 : AOI221_X1 port map( B1 => n16433, B2 => net226968, C1 => n16430, C2 
                           => net226967, A => n13732, ZN => n13731);
   U8403 : AOI221_X1 port map( B1 => n16421, B2 => net226971, C1 => n16418, C2 
                           => net226969, A => n13733, ZN => n13730);
   U8404 : AOI22_X1 port map( A1 => n16214, A2 => net226988, B1 => n16213, B2 
                           => registers_68_5_port, ZN => n13687);
   U8405 : AOI221_X1 port map( B1 => n16433, B2 => net226986, C1 => n16430, C2 
                           => net226985, A => n13690, ZN => n13689);
   U8406 : AOI221_X1 port map( B1 => n16421, B2 => net226989, C1 => n16418, C2 
                           => net226987, A => n13691, ZN => n13688);
   U8407 : AOI22_X1 port map( A1 => n16214, A2 => net227006, B1 => n16213, B2 
                           => registers_68_6_port, ZN => n13645);
   U8408 : AOI221_X1 port map( B1 => n16433, B2 => net227004, C1 => n16430, C2 
                           => net227003, A => n13648, ZN => n13647);
   U8409 : AOI221_X1 port map( B1 => n16421, B2 => net227007, C1 => n16418, C2 
                           => net227005, A => n13649, ZN => n13646);
   U8410 : AOI22_X1 port map( A1 => n16214, A2 => net227024, B1 => n16213, B2 
                           => registers_68_7_port, ZN => n13603);
   U8411 : AOI221_X1 port map( B1 => n16433, B2 => net227022, C1 => n16430, C2 
                           => net227021, A => n13606, ZN => n13605);
   U8412 : AOI221_X1 port map( B1 => n16421, B2 => net227025, C1 => n16418, C2 
                           => net227023, A => n13607, ZN => n13604);
   U8413 : AOI22_X1 port map( A1 => n16214, A2 => net227042, B1 => n16212, B2 
                           => registers_68_8_port, ZN => n13561);
   U8414 : AOI221_X1 port map( B1 => n16433, B2 => net227040, C1 => n16430, C2 
                           => net227039, A => n13564, ZN => n13563);
   U8415 : AOI221_X1 port map( B1 => n16421, B2 => net227043, C1 => n16418, C2 
                           => net227041, A => n13565, ZN => n13562);
   U8416 : AOI22_X1 port map( A1 => n16214, A2 => net227060, B1 => n16212, B2 
                           => registers_68_9_port, ZN => n13519);
   U8417 : AOI221_X1 port map( B1 => n16433, B2 => net227058, C1 => n16430, C2 
                           => net227057, A => n13522, ZN => n13521);
   U8418 : AOI221_X1 port map( B1 => n16421, B2 => net227061, C1 => n16418, C2 
                           => net227059, A => n13523, ZN => n13520);
   U8419 : AOI22_X1 port map( A1 => n16214, A2 => net227078, B1 => n16212, B2 
                           => registers_68_10_port, ZN => n13477);
   U8420 : AOI221_X1 port map( B1 => n16433, B2 => net227076, C1 => n16430, C2 
                           => net227075, A => n13480, ZN => n13479);
   U8421 : AOI221_X1 port map( B1 => n16421, B2 => net227079, C1 => n16418, C2 
                           => net227077, A => n13481, ZN => n13478);
   U8422 : AOI22_X1 port map( A1 => n16214, A2 => net227096, B1 => n16212, B2 
                           => registers_68_11_port, ZN => n13435);
   U8423 : AOI221_X1 port map( B1 => n16433, B2 => net227094, C1 => n16430, C2 
                           => net227093, A => n13438, ZN => n13437);
   U8424 : AOI221_X1 port map( B1 => n16421, B2 => net227097, C1 => n16418, C2 
                           => net227095, A => n13439, ZN => n13436);
   U8425 : AOI22_X1 port map( A1 => n16215, A2 => net227114, B1 => n16212, B2 
                           => registers_68_12_port, ZN => n13393);
   U8426 : AOI221_X1 port map( B1 => n16434, B2 => net227112, C1 => n16431, C2 
                           => net227111, A => n13396, ZN => n13395);
   U8427 : AOI221_X1 port map( B1 => n16422, B2 => net227115, C1 => n16419, C2 
                           => net227113, A => n13397, ZN => n13394);
   U8428 : AOI22_X1 port map( A1 => n16215, A2 => net227132, B1 => n16212, B2 
                           => registers_68_13_port, ZN => n13351);
   U8429 : AOI221_X1 port map( B1 => n16434, B2 => net227130, C1 => n16431, C2 
                           => net227129, A => n13354, ZN => n13353);
   U8430 : AOI221_X1 port map( B1 => n16422, B2 => net227133, C1 => n16419, C2 
                           => net227131, A => n13355, ZN => n13352);
   U8431 : AOI22_X1 port map( A1 => n16215, A2 => net227150, B1 => n16212, B2 
                           => registers_68_14_port, ZN => n13309);
   U8432 : AOI221_X1 port map( B1 => n16434, B2 => net227148, C1 => n16431, C2 
                           => net227147, A => n13312, ZN => n13311);
   U8433 : AOI221_X1 port map( B1 => n16422, B2 => net227151, C1 => n16419, C2 
                           => net227149, A => n13313, ZN => n13310);
   U8434 : AOI22_X1 port map( A1 => n16215, A2 => net227168, B1 => n16212, B2 
                           => registers_68_15_port, ZN => n13267);
   U8435 : AOI221_X1 port map( B1 => n16434, B2 => net227166, C1 => n16431, C2 
                           => net227165, A => n13270, ZN => n13269);
   U8436 : AOI221_X1 port map( B1 => n16422, B2 => net227169, C1 => n16419, C2 
                           => net227167, A => n13271, ZN => n13268);
   U8437 : AOI22_X1 port map( A1 => n16215, A2 => net227186, B1 => n16212, B2 
                           => registers_68_16_port, ZN => n13225);
   U8438 : AOI221_X1 port map( B1 => n16434, B2 => net227184, C1 => n16431, C2 
                           => net227183, A => n13228, ZN => n13227);
   U8439 : AOI221_X1 port map( B1 => n16422, B2 => net227187, C1 => n16419, C2 
                           => net227185, A => n13229, ZN => n13226);
   U8440 : AOI22_X1 port map( A1 => n16215, A2 => net227204, B1 => n16212, B2 
                           => registers_68_17_port, ZN => n13183);
   U8441 : AOI221_X1 port map( B1 => n16434, B2 => net227202, C1 => n16431, C2 
                           => net227201, A => n13186, ZN => n13185);
   U8442 : AOI221_X1 port map( B1 => n16422, B2 => net227205, C1 => n16419, C2 
                           => net227203, A => n13187, ZN => n13184);
   U8443 : AOI22_X1 port map( A1 => n16215, A2 => net227222, B1 => n16212, B2 
                           => registers_68_18_port, ZN => n13141);
   U8444 : AOI221_X1 port map( B1 => n16434, B2 => net227220, C1 => n16431, C2 
                           => net227219, A => n13144, ZN => n13143);
   U8445 : AOI221_X1 port map( B1 => n16422, B2 => net227223, C1 => n16419, C2 
                           => net227221, A => n13145, ZN => n13142);
   U8446 : AOI22_X1 port map( A1 => n16215, A2 => net227240, B1 => n16212, B2 
                           => registers_68_19_port, ZN => n13099);
   U8447 : AOI221_X1 port map( B1 => n16434, B2 => net227238, C1 => n16431, C2 
                           => net227237, A => n13102, ZN => n13101);
   U8448 : AOI221_X1 port map( B1 => n16422, B2 => net227241, C1 => n16419, C2 
                           => net227239, A => n13103, ZN => n13100);
   U8449 : AOI22_X1 port map( A1 => n16215, A2 => net227258, B1 => n16211, B2 
                           => registers_68_20_port, ZN => n13057);
   U8450 : AOI221_X1 port map( B1 => n16434, B2 => net227256, C1 => n16431, C2 
                           => net227255, A => n13060, ZN => n13059);
   U8451 : AOI221_X1 port map( B1 => n16422, B2 => net227259, C1 => n16419, C2 
                           => net227257, A => n13061, ZN => n13058);
   U8452 : AOI22_X1 port map( A1 => n16215, A2 => net227276, B1 => n16211, B2 
                           => registers_68_21_port, ZN => n13015);
   U8453 : AOI221_X1 port map( B1 => n16434, B2 => net227274, C1 => n16431, C2 
                           => net227273, A => n13018, ZN => n13017);
   U8454 : AOI221_X1 port map( B1 => n16422, B2 => net227277, C1 => n16419, C2 
                           => net227275, A => n13019, ZN => n13016);
   U8455 : AOI22_X1 port map( A1 => n16215, A2 => net227294, B1 => n16211, B2 
                           => registers_68_22_port, ZN => n12973);
   U8456 : AOI221_X1 port map( B1 => n16434, B2 => net227292, C1 => n16431, C2 
                           => net227291, A => n12976, ZN => n12975);
   U8457 : AOI221_X1 port map( B1 => n16422, B2 => net227295, C1 => n16419, C2 
                           => net227293, A => n12977, ZN => n12974);
   U8458 : AOI22_X1 port map( A1 => n16215, A2 => net227312, B1 => n16211, B2 
                           => registers_68_23_port, ZN => n12931);
   U8459 : AOI221_X1 port map( B1 => n16434, B2 => net227310, C1 => n16431, C2 
                           => net227309, A => n12934, ZN => n12933);
   U8460 : AOI221_X1 port map( B1 => n16422, B2 => net227313, C1 => n16419, C2 
                           => net227311, A => n12935, ZN => n12932);
   U8461 : AOI22_X1 port map( A1 => n16466, A2 => net226970, B1 => n16463, B2 
                           => registers_68_4_port, ZN => n11800);
   U8462 : AOI221_X1 port map( B1 => n16687, B2 => net226968, C1 => n16682, C2 
                           => net226967, A => n11803, ZN => n11802);
   U8463 : AOI221_X1 port map( B1 => n16675, B2 => net226971, C1 => n16670, C2 
                           => net226969, A => n11804, ZN => n11801);
   U8464 : AOI22_X1 port map( A1 => n16468, A2 => net227024, B1 => n16465, B2 
                           => registers_68_7_port, ZN => n11671);
   U8465 : AOI221_X1 port map( B1 => n16686, B2 => net227022, C1 => n16684, C2 
                           => net227021, A => n11674, ZN => n11673);
   U8466 : AOI221_X1 port map( B1 => n16674, B2 => net227025, C1 => n16672, C2 
                           => net227023, A => n11675, ZN => n11672);
   U8467 : AOI22_X1 port map( A1 => n16468, A2 => net227042, B1 => n16465, B2 
                           => registers_68_8_port, ZN => n11628);
   U8468 : AOI221_X1 port map( B1 => n16686, B2 => net227040, C1 => n16684, C2 
                           => net227039, A => n11631, ZN => n11630);
   U8469 : AOI221_X1 port map( B1 => n16674, B2 => net227043, C1 => n16672, C2 
                           => net227041, A => n11632, ZN => n11629);
   U8470 : AOI22_X1 port map( A1 => n16468, A2 => net227060, B1 => n16465, B2 
                           => registers_68_9_port, ZN => n11585);
   U8471 : AOI221_X1 port map( B1 => n16686, B2 => net227058, C1 => n16684, C2 
                           => net227057, A => n11588, ZN => n11587);
   U8472 : AOI221_X1 port map( B1 => n16674, B2 => net227061, C1 => n16672, C2 
                           => net227059, A => n11589, ZN => n11586);
   U8473 : AOI22_X1 port map( A1 => n16468, A2 => net227078, B1 => n16465, B2 
                           => registers_68_10_port, ZN => n11542);
   U8474 : AOI221_X1 port map( B1 => n16686, B2 => net227076, C1 => n16684, C2 
                           => net227075, A => n11545, ZN => n11544);
   U8475 : AOI221_X1 port map( B1 => n16674, B2 => net227079, C1 => n16672, C2 
                           => net227077, A => n11546, ZN => n11543);
   U8476 : AOI22_X1 port map( A1 => n16467, A2 => net227096, B1 => n16464, B2 
                           => registers_68_11_port, ZN => n11499);
   U8477 : AOI221_X1 port map( B1 => n16686, B2 => net227094, C1 => n16683, C2 
                           => net227093, A => n11502, ZN => n11501);
   U8478 : AOI221_X1 port map( B1 => n16674, B2 => net227097, C1 => n16671, C2 
                           => net227095, A => n11503, ZN => n11500);
   U8479 : AOI22_X1 port map( A1 => n16467, A2 => net227114, B1 => n16464, B2 
                           => registers_68_12_port, ZN => n11455);
   U8480 : AOI221_X1 port map( B1 => n16686, B2 => net227112, C1 => n16683, C2 
                           => net227111, A => n11458, ZN => n11457);
   U8481 : AOI221_X1 port map( B1 => n16674, B2 => net227115, C1 => n16671, C2 
                           => net227113, A => n11459, ZN => n11456);
   U8482 : AOI22_X1 port map( A1 => n16467, A2 => net227132, B1 => n16464, B2 
                           => registers_68_13_port, ZN => n11412);
   U8483 : AOI221_X1 port map( B1 => n16686, B2 => net227130, C1 => n16683, C2 
                           => net227129, A => n11415, ZN => n11414);
   U8484 : AOI221_X1 port map( B1 => n16674, B2 => net227133, C1 => n16671, C2 
                           => net227131, A => n11416, ZN => n11413);
   U8485 : AOI22_X1 port map( A1 => n16467, A2 => net227150, B1 => n16464, B2 
                           => registers_68_14_port, ZN => n11369);
   U8486 : AOI221_X1 port map( B1 => n16686, B2 => net227148, C1 => n16683, C2 
                           => net227147, A => n11372, ZN => n11371);
   U8487 : AOI221_X1 port map( B1 => n16674, B2 => net227151, C1 => n16671, C2 
                           => net227149, A => n11373, ZN => n11370);
   U8488 : AOI22_X1 port map( A1 => n16467, A2 => net227168, B1 => n16464, B2 
                           => registers_68_15_port, ZN => n11326);
   U8489 : AOI221_X1 port map( B1 => n16686, B2 => net227166, C1 => n16683, C2 
                           => net227165, A => n11329, ZN => n11328);
   U8490 : AOI221_X1 port map( B1 => n16674, B2 => net227169, C1 => n16671, C2 
                           => net227167, A => n11330, ZN => n11327);
   U8491 : AOI22_X1 port map( A1 => n16467, A2 => net227186, B1 => n16464, B2 
                           => registers_68_16_port, ZN => n11283);
   U8492 : AOI221_X1 port map( B1 => n16686, B2 => net227184, C1 => n16683, C2 
                           => net227183, A => n11286, ZN => n11285);
   U8493 : AOI221_X1 port map( B1 => n16674, B2 => net227187, C1 => n16671, C2 
                           => net227185, A => n11287, ZN => n11284);
   U8494 : AOI22_X1 port map( A1 => n16467, A2 => net227204, B1 => n16464, B2 
                           => registers_68_17_port, ZN => n11240);
   U8495 : AOI221_X1 port map( B1 => n16686, B2 => net227202, C1 => n16683, C2 
                           => net227201, A => n11243, ZN => n11242);
   U8496 : AOI221_X1 port map( B1 => n16674, B2 => net227205, C1 => n16671, C2 
                           => net227203, A => n11244, ZN => n11241);
   U8497 : AOI22_X1 port map( A1 => n16467, A2 => net227222, B1 => n16464, B2 
                           => registers_68_18_port, ZN => n11197);
   U8498 : AOI221_X1 port map( B1 => n16685, B2 => net227220, C1 => n16683, C2 
                           => net227219, A => n11200, ZN => n11199);
   U8499 : AOI221_X1 port map( B1 => n16673, B2 => net227223, C1 => n16671, C2 
                           => net227221, A => n11201, ZN => n11198);
   U8500 : AOI22_X1 port map( A1 => n16467, A2 => net227240, B1 => n16464, B2 
                           => registers_68_19_port, ZN => n11154);
   U8501 : AOI221_X1 port map( B1 => n16685, B2 => net227238, C1 => n16683, C2 
                           => net227237, A => n11157, ZN => n11156);
   U8502 : AOI221_X1 port map( B1 => n16673, B2 => net227241, C1 => n16671, C2 
                           => net227239, A => n11158, ZN => n11155);
   U8503 : AOI22_X1 port map( A1 => n16467, A2 => net227258, B1 => n16464, B2 
                           => registers_68_20_port, ZN => n11111);
   U8504 : AOI221_X1 port map( B1 => n16685, B2 => net227256, C1 => n16683, C2 
                           => net227255, A => n11114, ZN => n11113);
   U8505 : AOI221_X1 port map( B1 => n16673, B2 => net227259, C1 => n16671, C2 
                           => net227257, A => n11115, ZN => n11112);
   U8506 : AOI22_X1 port map( A1 => n16467, A2 => net227276, B1 => n16464, B2 
                           => registers_68_21_port, ZN => n11068);
   U8507 : AOI221_X1 port map( B1 => n16685, B2 => net227274, C1 => n16683, C2 
                           => net227273, A => n11071, ZN => n11070);
   U8508 : AOI221_X1 port map( B1 => n16673, B2 => net227277, C1 => n16671, C2 
                           => net227275, A => n11072, ZN => n11069);
   U8509 : AOI22_X1 port map( A1 => n16467, A2 => net227294, B1 => n16464, B2 
                           => registers_68_22_port, ZN => n11025);
   U8510 : AOI221_X1 port map( B1 => n16685, B2 => net227292, C1 => n16683, C2 
                           => net227291, A => n11028, ZN => n11027);
   U8511 : AOI221_X1 port map( B1 => n16673, B2 => net227295, C1 => n16671, C2 
                           => net227293, A => n11029, ZN => n11026);
   U8512 : AOI22_X1 port map( A1 => n16467, A2 => net227312, B1 => n16464, B2 
                           => registers_68_23_port, ZN => n10982);
   U8513 : AOI221_X1 port map( B1 => n16686, B2 => net227310, C1 => n16683, C2 
                           => net227309, A => n10985, ZN => n10984);
   U8514 : AOI221_X1 port map( B1 => n16674, B2 => net227313, C1 => n16671, C2 
                           => net227311, A => n10986, ZN => n10983);
   U8515 : AOI22_X1 port map( A1 => n16466, A2 => net227330, B1 => n16463, B2 
                           => registers_68_24_port, ZN => n10939);
   U8516 : AOI221_X1 port map( B1 => n16685, B2 => net227328, C1 => n16682, C2 
                           => net227327, A => n10942, ZN => n10941);
   U8517 : AOI221_X1 port map( B1 => n16673, B2 => net227331, C1 => n16670, C2 
                           => net227329, A => n10943, ZN => n10940);
   U8518 : AOI22_X1 port map( A1 => n16466, A2 => net227348, B1 => n16463, B2 
                           => registers_68_25_port, ZN => n10896);
   U8519 : AOI221_X1 port map( B1 => n16685, B2 => net227346, C1 => n16682, C2 
                           => net227345, A => n10899, ZN => n10898);
   U8520 : AOI221_X1 port map( B1 => n16673, B2 => net227349, C1 => n16670, C2 
                           => net227347, A => n10900, ZN => n10897);
   U8521 : AOI22_X1 port map( A1 => n16466, A2 => net227366, B1 => n16463, B2 
                           => registers_68_26_port, ZN => n10853);
   U8522 : AOI221_X1 port map( B1 => n16685, B2 => net227364, C1 => n16682, C2 
                           => net227363, A => n10856, ZN => n10855);
   U8523 : AOI221_X1 port map( B1 => n16673, B2 => net227367, C1 => n16670, C2 
                           => net227365, A => n10857, ZN => n10854);
   U8524 : AOI22_X1 port map( A1 => n16466, A2 => net227384, B1 => n16463, B2 
                           => registers_68_27_port, ZN => n10810);
   U8525 : AOI221_X1 port map( B1 => n16685, B2 => net227382, C1 => n16682, C2 
                           => net227381, A => n10813, ZN => n10812);
   U8526 : AOI221_X1 port map( B1 => n16673, B2 => net227385, C1 => n16670, C2 
                           => net227383, A => n10814, ZN => n10811);
   U8527 : AOI22_X1 port map( A1 => n16466, A2 => net227402, B1 => n16463, B2 
                           => registers_68_28_port, ZN => n10767);
   U8528 : AOI221_X1 port map( B1 => n16685, B2 => net227400, C1 => n16682, C2 
                           => net227399, A => n10770, ZN => n10769);
   U8529 : AOI221_X1 port map( B1 => n16673, B2 => net227403, C1 => n16670, C2 
                           => net227401, A => n10771, ZN => n10768);
   U8530 : AOI22_X1 port map( A1 => n16466, A2 => net227420, B1 => n16463, B2 
                           => registers_68_29_port, ZN => n10724);
   U8531 : AOI221_X1 port map( B1 => n16685, B2 => net227418, C1 => n16682, C2 
                           => net227417, A => n10727, ZN => n10726);
   U8532 : AOI221_X1 port map( B1 => n16673, B2 => net227421, C1 => n16670, C2 
                           => net227419, A => n10728, ZN => n10725);
   U8533 : AOI22_X1 port map( A1 => n16466, A2 => net227438, B1 => n16463, B2 
                           => registers_68_30_port, ZN => n10665);
   U8534 : AOI221_X1 port map( B1 => n16685, B2 => net227436, C1 => n16682, C2 
                           => net227435, A => n10668, ZN => n10667);
   U8535 : AOI221_X1 port map( B1 => n16673, B2 => net227439, C1 => n16670, C2 
                           => net227437, A => n10669, ZN => n10666);
   U8536 : AND4_X1 port map( A1 => n14233, A2 => wr, A3 => add_wr(3), A4 => 
                           add_wr(4), ZN => n14223);
   U8537 : AND2_X1 port map( A1 => n14016, A2 => r590_carry_5_port, ZN => 
                           n14194);
   U8538 : NOR4_X1 port map( A1 => n13989, A2 => add_rd2(0), A3 => add_rd2(4), 
                           A4 => add_rd2(3), ZN => n13974);
   U8539 : INV_X1 port map( A => n13985, ZN => n13989);
   U8540 : AND4_X1 port map( A1 => n14026, A2 => n14027, A3 => n14028, A4 => 
                           n14029, ZN => n14024);
   U8541 : XNOR2_X1 port map( A => swp_2_port, B => N9909, ZN => n14027);
   U8542 : XNOR2_X1 port map( A => swp_0_port, B => N9641, ZN => n14026);
   U8543 : XNOR2_X1 port map( A => swp_3_port, B => N9910, ZN => n14028);
   U8544 : NOR4_X1 port map( A1 => n12508, A2 => add_rd1(0), A3 => add_rd1(4), 
                           A4 => add_rd1(3), ZN => n12493);
   U8545 : INV_X1 port map( A => n12504, ZN => n12508);
   U8546 : INV_X1 port map( A => n11859, ZN => n8037);
   U8547 : AOI221_X1 port map( B1 => n17989, B2 => registers_56_3_port, C1 => 
                           n17991, C2 => datain(3), A => n18049, ZN => n11859);
   U8548 : INV_X1 port map( A => n11853, ZN => n8043);
   U8549 : AOI221_X1 port map( B1 => n16989, B2 => registers_42_3_port, C1 => 
                           n16991, C2 => datain(3), A => n18049, ZN => n11853);
   U8550 : INV_X1 port map( A => n11848, ZN => n8048);
   U8551 : AOI221_X1 port map( B1 => n17150, B2 => registers_29_3_port, C1 => 
                           n17152, C2 => datain(3), A => n18048, ZN => n11848);
   U8552 : INV_X1 port map( A => n10448, ZN => n8134);
   U8553 : AOI221_X1 port map( B1 => n17216, B2 => registers_23_4_port, C1 => 
                           n17218, C2 => datain(4), A => n18048, ZN => n10448);
   U8554 : INV_X1 port map( A => n10444, ZN => n8138);
   U8555 : AOI221_X1 port map( B1 => n17268, B2 => registers_19_4_port, C1 => 
                           n17270, C2 => datain(4), A => n18048, ZN => n10444);
   U8556 : INV_X1 port map( A => n10416, ZN => n8165);
   U8557 : AOI221_X1 port map( B1 => n17989, B2 => registers_56_4_port, C1 => 
                           n17992, C2 => datain(4), A => n18048, ZN => n10416);
   U8558 : INV_X1 port map( A => n10413, ZN => n8168);
   U8559 : AOI221_X1 port map( B1 => n16866, B2 => net226980, C1 => n16868, C2 
                           => datain(4), A => n18047, ZN => n10413);
   U8560 : INV_X1 port map( A => n10410, ZN => n8171);
   U8561 : AOI221_X1 port map( B1 => n16900, B2 => registers_50_4_port, C1 => 
                           n16902, C2 => datain(4), A => n18047, ZN => n10410);
   U8562 : INV_X1 port map( A => n10405, ZN => n8176);
   U8563 : AOI221_X1 port map( B1 => n17150, B2 => registers_29_4_port, C1 => 
                           n17152, C2 => datain(4), A => n18047, ZN => n10405);
   U8564 : INV_X1 port map( A => n10306, ZN => n8237);
   U8565 : AOI221_X1 port map( B1 => n17989, B2 => registers_56_5_port, C1 => 
                           n17991, C2 => datain(5), A => n18047, ZN => n10306);
   U8566 : INV_X1 port map( A => n10303, ZN => n8240);
   U8567 : AOI221_X1 port map( B1 => n16866, B2 => net227000, C1 => n16868, C2 
                           => datain(5), A => n18046, ZN => n10303);
   U8568 : INV_X1 port map( A => n10300, ZN => n8243);
   U8569 : AOI221_X1 port map( B1 => n16900, B2 => registers_50_5_port, C1 => 
                           n16902, C2 => datain(5), A => n18046, ZN => n10300);
   U8570 : INV_X1 port map( A => n10292, ZN => n8251);
   U8571 : AOI221_X1 port map( B1 => n16989, B2 => registers_42_5_port, C1 => 
                           n16991, C2 => datain(5), A => n18046, ZN => n10292);
   U8572 : INV_X1 port map( A => n10288, ZN => n8254);
   U8573 : AOI221_X1 port map( B1 => n17534, B2 => net227003, C1 => n17536, C2 
                           => datain(6), A => n18046, ZN => n10288);
   U8574 : INV_X1 port map( A => n10287, ZN => n8255);
   U8575 : AOI221_X1 port map( B1 => n17548, B2 => net227004, C1 => n17550, C2 
                           => datain(6), A => n18045, ZN => n10287);
   U8576 : INV_X1 port map( A => n10286, ZN => n8256);
   U8577 : AOI221_X1 port map( B1 => n17562, B2 => registers_68_6_port, C1 => 
                           n17564, C2 => datain(6), A => n18045, ZN => n10286);
   U8578 : INV_X1 port map( A => n10283, ZN => n8258);
   U8579 : AOI221_X1 port map( B1 => n17589, B2 => net227005, C1 => n17591, C2 
                           => datain(6), A => n18045, ZN => n10283);
   U8580 : INV_X1 port map( A => n10282, ZN => n8259);
   U8581 : AOI221_X1 port map( B1 => n17603, B2 => net227006, C1 => n17605, C2 
                           => datain(6), A => n18045, ZN => n10282);
   U8582 : INV_X1 port map( A => n10280, ZN => n8260);
   U8583 : AOI221_X1 port map( B1 => n17617, B2 => net227007, C1 => n17619, C2 
                           => datain(6), A => n18049, ZN => n10280);
   U8584 : NOR2_X1 port map( A1 => n10187, A2 => n14017, ZN => n14021);
   U8585 : OAI22_X1 port map( A1 => n14820, A2 => n14000, B1 => 
                           r590_carry_5_port, B2 => n14001, ZN => n10182);
   U8586 : OAI22_X1 port map( A1 => n3043, A2 => n14000, B1 => n14002, B2 => 
                           n14001, ZN => n10181);
   U8587 : NOR2_X1 port map( A1 => call, A2 => n14003, ZN => n14002);
   U8588 : NOR2_X1 port map( A1 => r590_carry_5_port, A2 => n14021, ZN => 
                           n14011);
   U8589 : NAND2_X1 port map( A1 => add_wr(1), A2 => n14229, ZN => n14220);
   U8590 : NAND2_X1 port map( A1 => add_wr(1), A2 => add_wr(0), ZN => n12412);
   U8591 : NOR2_X1 port map( A1 => n13984, A2 => add_rd2(1), ZN => n13905);
   U8592 : NOR2_X1 port map( A1 => n12503, A2 => add_rd1(1), ZN => n12424);
   U8593 : AND2_X1 port map( A1 => add_rd2(1), A2 => n13984, ZN => n13902);
   U8594 : AND2_X1 port map( A1 => add_rd2(1), A2 => add_rd2(2), ZN => n13903);
   U8595 : AND2_X1 port map( A1 => add_rd1(1), A2 => n12503, ZN => n12421);
   U8596 : OR2_X1 port map( A1 => n14229, A2 => add_wr(1), ZN => n14217);
   U8597 : AND2_X1 port map( A1 => add_rd1(1), A2 => add_rd1(2), ZN => n12422);
   U8598 : NAND2_X1 port map( A1 => n7685, A2 => n17823, ZN => n10148);
   U8599 : NAND2_X1 port map( A1 => n7684, A2 => n17823, ZN => n10149);
   U8600 : NAND2_X1 port map( A1 => n7683, A2 => n17823, ZN => n10150);
   U8601 : NAND2_X1 port map( A1 => n7682, A2 => n17823, ZN => n10151);
   U8602 : NAND2_X1 port map( A1 => n7681, A2 => n17823, ZN => n10152);
   U8603 : NAND2_X1 port map( A1 => n7680, A2 => n17823, ZN => n10153);
   U8604 : NAND2_X1 port map( A1 => n7679, A2 => n17823, ZN => n10154);
   U8605 : NAND2_X1 port map( A1 => n7678, A2 => n17823, ZN => n10155);
   U8606 : NAND2_X1 port map( A1 => n7677, A2 => n17823, ZN => n10156);
   U8607 : NAND2_X1 port map( A1 => n7676, A2 => n17823, ZN => n10157);
   U8608 : NAND2_X1 port map( A1 => n7675, A2 => n17823, ZN => n10158);
   U8609 : NAND2_X1 port map( A1 => n7674, A2 => n17823, ZN => n10159);
   U8610 : NAND2_X1 port map( A1 => n7673, A2 => n17825, ZN => n10160);
   U8611 : NAND2_X1 port map( A1 => n7672, A2 => n17825, ZN => n10161);
   U8612 : NAND2_X1 port map( A1 => n7671, A2 => n17825, ZN => n10162);
   U8613 : NAND2_X1 port map( A1 => n7670, A2 => n17825, ZN => n10163);
   U8614 : NAND2_X1 port map( A1 => n7669, A2 => n17825, ZN => n10164);
   U8615 : NAND2_X1 port map( A1 => n7668, A2 => n17825, ZN => n10165);
   U8616 : NAND2_X1 port map( A1 => n7667, A2 => n17825, ZN => n10166);
   U8617 : NAND2_X1 port map( A1 => n7666, A2 => n17825, ZN => n10167);
   U8618 : NAND2_X1 port map( A1 => n7665, A2 => n17825, ZN => n10168);
   U8619 : NAND2_X1 port map( A1 => n7664, A2 => n17825, ZN => n10169);
   U8620 : NAND2_X1 port map( A1 => n7663, A2 => n17824, ZN => n10170);
   U8621 : NAND2_X1 port map( A1 => n7662, A2 => n17824, ZN => n10171);
   U8622 : NAND2_X1 port map( A1 => n7693, A2 => n17824, ZN => n10140);
   U8623 : NAND2_X1 port map( A1 => n7692, A2 => n17824, ZN => n10141);
   U8624 : NAND2_X1 port map( A1 => n7691, A2 => n17824, ZN => n10142);
   U8625 : NAND2_X1 port map( A1 => n7690, A2 => n17824, ZN => n10143);
   U8626 : NAND2_X1 port map( A1 => n7689, A2 => n17824, ZN => n10144);
   U8627 : NAND2_X1 port map( A1 => n7688, A2 => n17824, ZN => n10145);
   U8628 : NAND2_X1 port map( A1 => n7687, A2 => n17824, ZN => n10146);
   U8629 : NAND2_X1 port map( A1 => n7686, A2 => n17824, ZN => n10147);
   U8630 : OR2_X1 port map( A1 => n18050, A2 => swp_5_port, ZN => n10173);
   U8631 : AND2_X1 port map( A1 => n18044, A2 => swp_4_port, ZN => n10172);
   U8632 : AND2_X1 port map( A1 => n18044, A2 => swp_3_port, ZN => n10174);
   U8633 : AND2_X1 port map( A1 => n18044, A2 => swp_2_port, ZN => n10176);
   U8634 : AND2_X1 port map( A1 => n18044, A2 => swp_1_port, ZN => n10178);
   U8635 : AND2_X1 port map( A1 => n18044, A2 => swp_0_port, ZN => n10184);
   U8636 : INV_X1 port map( A => call, ZN => n14020);
   U8637 : INV_X1 port map( A => wr, ZN => n12514);
   U8638 : NOR2_X1 port map( A1 => ret, A2 => call, ZN => n14005);
   U8639 : NAND3_X2 port map( A1 => n14240, A2 => n14239, A3 => N276, ZN => 
                           n14241);
   U8640 : CLKBUF_X1 port map( A => n12527, Z => n16417);
   U8641 : CLKBUF_X1 port map( A => n10525, Z => n16669);
   U8642 : INV_X1 port map( A => n16696, ZN => n16692);
   U8643 : CLKBUF_X1 port map( A => n7652, Z => n16730);
   U8644 : INV_X1 port map( A => n17455, ZN => n17451);
   U8645 : INV_X1 port map( A => n17581, ZN => n17577);
   U8646 : INV_X1 port map( A => n17834, ZN => n17825);
   U8647 : INV_X1 port map( A => n17855, ZN => n17838);
   U8648 : CLKBUF_X1 port map( A => n17854, Z => n17839);
   U8649 : CLKBUF_X1 port map( A => n17856, Z => n17840);
   U8650 : CLKBUF_X1 port map( A => n17856, Z => n17841);
   U8651 : CLKBUF_X1 port map( A => n17856, Z => n17842);
   U8652 : CLKBUF_X1 port map( A => n17856, Z => n17843);
   U8653 : CLKBUF_X1 port map( A => n17856, Z => n17844);
   U8654 : CLKBUF_X1 port map( A => n17856, Z => n17845);
   U8655 : CLKBUF_X1 port map( A => n17856, Z => n17846);
   U8656 : CLKBUF_X1 port map( A => n17853, Z => n17847);
   U8657 : CLKBUF_X1 port map( A => n17840, Z => n17848);
   U8658 : CLKBUF_X1 port map( A => n17845, Z => n17849);
   U8659 : CLKBUF_X1 port map( A => n17856, Z => n17850);
   U8660 : CLKBUF_X1 port map( A => n17856, Z => n17851);
   U8661 : CLKBUF_X1 port map( A => n17856, Z => n17852);
   U8662 : CLKBUF_X1 port map( A => n17856, Z => n17853);
   U8663 : CLKBUF_X1 port map( A => n17856, Z => n17854);
   U8664 : CLKBUF_X1 port map( A => n17856, Z => n17855);
   U8665 : INV_X1 port map( A => n17835, ZN => n17856);
   U8666 : INV_X1 port map( A => n17877, ZN => n17860);
   U8667 : CLKBUF_X1 port map( A => n17878, Z => n17861);
   U8668 : CLKBUF_X1 port map( A => n17878, Z => n17862);
   U8669 : CLKBUF_X1 port map( A => n17878, Z => n17863);
   U8670 : CLKBUF_X1 port map( A => n17878, Z => n17864);
   U8671 : CLKBUF_X1 port map( A => n17878, Z => n17865);
   U8672 : CLKBUF_X1 port map( A => n17878, Z => n17866);
   U8673 : CLKBUF_X1 port map( A => n17865, Z => n17867);
   U8674 : CLKBUF_X1 port map( A => n17861, Z => n17868);
   U8675 : CLKBUF_X1 port map( A => n17866, Z => n17869);
   U8676 : CLKBUF_X1 port map( A => n17864, Z => n17870);
   U8677 : CLKBUF_X1 port map( A => n17876, Z => n17871);
   U8678 : CLKBUF_X1 port map( A => n17878, Z => n17872);
   U8679 : CLKBUF_X1 port map( A => n17878, Z => n17873);
   U8680 : CLKBUF_X1 port map( A => n17878, Z => n17874);
   U8681 : CLKBUF_X1 port map( A => n17863, Z => n17875);
   U8682 : CLKBUF_X1 port map( A => n17878, Z => n17876);
   U8683 : CLKBUF_X1 port map( A => n17878, Z => n17877);
   U8684 : INV_X1 port map( A => n17857, ZN => n17878);
   U8685 : INV_X1 port map( A => n17899, ZN => n17882);
   U8686 : CLKBUF_X1 port map( A => n17900, Z => n17883);
   U8687 : CLKBUF_X1 port map( A => n17887, Z => n17884);
   U8688 : CLKBUF_X1 port map( A => n17900, Z => n17885);
   U8689 : CLKBUF_X1 port map( A => n17900, Z => n17886);
   U8690 : CLKBUF_X1 port map( A => n17900, Z => n17887);
   U8691 : CLKBUF_X1 port map( A => n17900, Z => n17888);
   U8692 : CLKBUF_X1 port map( A => n17900, Z => n17889);
   U8693 : CLKBUF_X1 port map( A => n17900, Z => n17890);
   U8694 : CLKBUF_X1 port map( A => n17888, Z => n17891);
   U8695 : CLKBUF_X1 port map( A => n17890, Z => n17892);
   U8696 : CLKBUF_X1 port map( A => n17883, Z => n17893);
   U8697 : CLKBUF_X1 port map( A => n17900, Z => n17894);
   U8698 : CLKBUF_X1 port map( A => n17898, Z => n17895);
   U8699 : CLKBUF_X1 port map( A => n17900, Z => n17896);
   U8700 : CLKBUF_X1 port map( A => n17889, Z => n17897);
   U8701 : CLKBUF_X1 port map( A => n17900, Z => n17898);
   U8702 : CLKBUF_X1 port map( A => n17900, Z => n17899);
   U8703 : INV_X1 port map( A => n17879, ZN => n17900);
   U8704 : INV_X1 port map( A => n17921, ZN => n17904);
   U8705 : CLKBUF_X1 port map( A => n17922, Z => n17905);
   U8706 : CLKBUF_X1 port map( A => n17922, Z => n17906);
   U8707 : CLKBUF_X1 port map( A => n17922, Z => n17907);
   U8708 : CLKBUF_X1 port map( A => n17922, Z => n17908);
   U8709 : CLKBUF_X1 port map( A => n17922, Z => n17909);
   U8710 : CLKBUF_X1 port map( A => n17922, Z => n17910);
   U8711 : CLKBUF_X1 port map( A => n17909, Z => n17911);
   U8712 : CLKBUF_X1 port map( A => n17905, Z => n17912);
   U8713 : CLKBUF_X1 port map( A => n17910, Z => n17913);
   U8714 : CLKBUF_X1 port map( A => n17908, Z => n17914);
   U8715 : CLKBUF_X1 port map( A => n17920, Z => n17915);
   U8716 : CLKBUF_X1 port map( A => n17922, Z => n17916);
   U8717 : CLKBUF_X1 port map( A => n17922, Z => n17917);
   U8718 : CLKBUF_X1 port map( A => n17922, Z => n17918);
   U8719 : CLKBUF_X1 port map( A => n17907, Z => n17919);
   U8720 : CLKBUF_X1 port map( A => n17922, Z => n17920);
   U8721 : CLKBUF_X1 port map( A => n17922, Z => n17921);
   U8722 : INV_X1 port map( A => n17901, ZN => n17922);
   U8723 : INV_X1 port map( A => n17942, ZN => n17925);
   U8724 : CLKBUF_X1 port map( A => n17943, Z => n17926);
   U8725 : CLKBUF_X1 port map( A => n17930, Z => n17927);
   U8726 : CLKBUF_X1 port map( A => n17943, Z => n17928);
   U8727 : CLKBUF_X1 port map( A => n17943, Z => n17929);
   U8728 : CLKBUF_X1 port map( A => n17943, Z => n17930);
   U8729 : CLKBUF_X1 port map( A => n17943, Z => n17931);
   U8730 : CLKBUF_X1 port map( A => n17943, Z => n17932);
   U8731 : CLKBUF_X1 port map( A => n17943, Z => n17933);
   U8732 : CLKBUF_X1 port map( A => n17931, Z => n17934);
   U8733 : CLKBUF_X1 port map( A => n17933, Z => n17935);
   U8734 : CLKBUF_X1 port map( A => n17926, Z => n17936);
   U8735 : CLKBUF_X1 port map( A => n17943, Z => n17937);
   U8736 : CLKBUF_X1 port map( A => n17941, Z => n17938);
   U8737 : CLKBUF_X1 port map( A => n17943, Z => n17939);
   U8738 : CLKBUF_X1 port map( A => n17932, Z => n17940);
   U8739 : CLKBUF_X1 port map( A => n17943, Z => n17941);
   U8740 : CLKBUF_X1 port map( A => n17943, Z => n17942);
   U8741 : INV_X1 port map( A => n4076, ZN => n17943);
   U8742 : INV_X1 port map( A => n17963, ZN => n17946);
   U8743 : CLKBUF_X1 port map( A => n17964, Z => n17947);
   U8744 : CLKBUF_X1 port map( A => n17964, Z => n17948);
   U8745 : CLKBUF_X1 port map( A => n17964, Z => n17949);
   U8746 : CLKBUF_X1 port map( A => n17964, Z => n17950);
   U8747 : CLKBUF_X1 port map( A => n17964, Z => n17951);
   U8748 : CLKBUF_X1 port map( A => n17964, Z => n17952);
   U8749 : CLKBUF_X1 port map( A => n17951, Z => n17953);
   U8750 : CLKBUF_X1 port map( A => n17947, Z => n17954);
   U8751 : CLKBUF_X1 port map( A => n17952, Z => n17955);
   U8752 : CLKBUF_X1 port map( A => n17950, Z => n17956);
   U8753 : CLKBUF_X1 port map( A => n17962, Z => n17957);
   U8754 : CLKBUF_X1 port map( A => n17964, Z => n17958);
   U8755 : CLKBUF_X1 port map( A => n17964, Z => n17959);
   U8756 : CLKBUF_X1 port map( A => n17964, Z => n17960);
   U8757 : CLKBUF_X1 port map( A => n17949, Z => n17961);
   U8758 : CLKBUF_X1 port map( A => n17964, Z => n17962);
   U8759 : CLKBUF_X1 port map( A => n17964, Z => n17963);
   U8760 : INV_X1 port map( A => n4073, ZN => n17964);
   U8761 : INV_X1 port map( A => n17984, ZN => n17967);
   U8762 : CLKBUF_X1 port map( A => n17985, Z => n17968);
   U8763 : CLKBUF_X1 port map( A => n17972, Z => n17969);
   U8764 : CLKBUF_X1 port map( A => n17985, Z => n17970);
   U8765 : CLKBUF_X1 port map( A => n17985, Z => n17971);
   U8766 : CLKBUF_X1 port map( A => n17985, Z => n17972);
   U8767 : CLKBUF_X1 port map( A => n17985, Z => n17973);
   U8768 : CLKBUF_X1 port map( A => n17985, Z => n17974);
   U8769 : CLKBUF_X1 port map( A => n17985, Z => n17975);
   U8770 : CLKBUF_X1 port map( A => n17973, Z => n17976);
   U8771 : CLKBUF_X1 port map( A => n17975, Z => n17977);
   U8772 : CLKBUF_X1 port map( A => n17968, Z => n17978);
   U8773 : CLKBUF_X1 port map( A => n17983, Z => n17979);
   U8774 : CLKBUF_X1 port map( A => n17985, Z => n17980);
   U8775 : CLKBUF_X1 port map( A => n17985, Z => n17981);
   U8776 : CLKBUF_X1 port map( A => n17974, Z => n17982);
   U8777 : CLKBUF_X1 port map( A => n17985, Z => n17983);
   U8778 : CLKBUF_X1 port map( A => n17985, Z => n17984);
   U8779 : INV_X1 port map( A => n4070, ZN => n17985);
   U8780 : INV_X1 port map( A => n18051, ZN => n18033);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N5_1 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0);  
         d_out : out std_logic_vector (4 downto 0));

end reg_N5_1;

architecture SYN_behav of reg_N5_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, n1, n6_port, n7, n8, n9 : std_logic;

begin
   
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n1);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n6_port);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n7);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n8);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n9);
   U3 : AND2_X1 port map( A1 => d_in(2), A2 => rst, ZN => N4);
   U4 : AND2_X1 port map( A1 => d_in(3), A2 => rst, ZN => N5);
   U5 : AND2_X1 port map( A1 => d_in(1), A2 => rst, ZN => N3);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U7 : AND2_X1 port map( A1 => rst, A2 => d_in(4), ZN => N6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N5_2 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0);  
         d_out : out std_logic_vector (4 downto 0));

end reg_N5_2;

architecture SYN_behav of reg_N5_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, n1, n6_port, n7, n8, n9 : std_logic;

begin
   
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n1);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n6_port);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n7);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n8);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n9);
   U3 : AND2_X1 port map( A1 => d_in(2), A2 => rst, ZN => N4);
   U4 : AND2_X1 port map( A1 => d_in(3), A2 => rst, ZN => N5);
   U5 : AND2_X1 port map( A1 => d_in(1), A2 => rst, ZN => N3);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U7 : AND2_X1 port map( A1 => rst, A2 => d_in(4), ZN => N6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N5_0 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0);  
         d_out : out std_logic_vector (4 downto 0));

end reg_N5_0;

architecture SYN_behav of reg_N5_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, n2_port, n3_port, n4_port, n5_port, n6_port : 
      std_logic;

begin
   
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n6_port);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n5_port);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n4_port);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n3_port);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n2_port);
   U3 : AND2_X1 port map( A1 => d_in(1), A2 => rst, ZN => N3);
   U4 : AND2_X1 port map( A1 => d_in(2), A2 => rst, ZN => N4);
   U5 : AND2_X1 port map( A1 => rst, A2 => d_in(4), ZN => N6);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(3), A2 => rst, ZN => N5);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N6_1 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (5 downto 0);  
         d_out : out std_logic_vector (5 downto 0));

end reg_N6_1;

architecture SYN_behav of reg_N6_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, n1, n7_port, n8, n9, n10, n11 : std_logic;

begin
   
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n1);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n7_port);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n8);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n9);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n10);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n11);
   U3 : AND2_X1 port map( A1 => rst, A2 => d_in(5), ZN => N7);
   U4 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U5 : AND2_X1 port map( A1 => d_in(1), A2 => rst, ZN => N3);
   U6 : AND2_X1 port map( A1 => d_in(2), A2 => rst, ZN => N4);
   U7 : AND2_X1 port map( A1 => d_in(3), A2 => rst, ZN => N5);
   U8 : AND2_X1 port map( A1 => d_in(4), A2 => rst, ZN => N6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N6_0 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (5 downto 0);  
         d_out : out std_logic_vector (5 downto 0));

end reg_N6_0;

architecture SYN_behav of reg_N6_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, n2_port, n3_port, n4_port, n5_port, n6_port, 
      n7_port : std_logic;

begin
   
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n7_port);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n6_port);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n5_port);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n4_port);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n3_port);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n2_port);
   U3 : AND2_X1 port map( A1 => d_in(3), A2 => rst, ZN => N5);
   U4 : AND2_X1 port map( A1 => d_in(4), A2 => rst, ZN => N6);
   U5 : AND2_X1 port map( A1 => rst, A2 => d_in(5), ZN => N7);
   U6 : AND2_X1 port map( A1 => d_in(2), A2 => rst, ZN => N4);
   U7 : AND2_X1 port map( A1 => d_in(0), A2 => rst, ZN => N2);
   U8 : AND2_X1 port map( A1 => d_in(1), A2 => rst, ZN => N3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity reg_N32_0 is

   port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);  
         d_out : out std_logic_vector (31 downto 0));

end reg_N32_0;

architecture SYN_behav of reg_N32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   d_out_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => d_out(31), QN
                           => n36);
   d_out_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => d_out(30), QN
                           => n37);
   d_out_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => d_out(29), QN
                           => n38);
   d_out_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => d_out(28), QN
                           => n39);
   d_out_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => d_out(27), QN
                           => n40);
   d_out_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => d_out(26), QN
                           => n41);
   d_out_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => d_out(25), QN
                           => n42);
   d_out_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => d_out(24), QN
                           => n43);
   d_out_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => d_out(23), QN
                           => n44);
   d_out_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => d_out(22), QN
                           => n45);
   d_out_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => d_out(21), QN
                           => n46);
   d_out_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => d_out(20), QN
                           => n47);
   d_out_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => d_out(19), QN
                           => n48);
   d_out_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => d_out(18), QN
                           => n49);
   d_out_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => d_out(17), QN
                           => n50);
   d_out_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => d_out(16), QN
                           => n51);
   d_out_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => d_out(15), QN
                           => n52);
   d_out_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => d_out(14), QN
                           => n53);
   d_out_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => d_out(13), QN
                           => n54);
   d_out_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => d_out(12), QN
                           => n55);
   d_out_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => d_out(11), QN
                           => n56);
   d_out_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => d_out(10), QN
                           => n57);
   d_out_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => d_out(9), QN 
                           => n58);
   d_out_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => d_out(8), QN 
                           => n59);
   d_out_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => d_out(7), QN =>
                           n60);
   d_out_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => d_out(6), QN =>
                           n61);
   d_out_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => d_out(5), QN =>
                           n62);
   d_out_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => d_out(4), QN =>
                           n63);
   d_out_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => d_out(3), QN =>
                           n64);
   d_out_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => d_out(2), QN =>
                           n65);
   d_out_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => d_out(1), QN =>
                           n66);
   d_out_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => d_out(0), QN =>
                           n67);
   U3 : BUF_X1 port map( A => rst, Z => n68);
   U4 : BUF_X1 port map( A => rst, Z => n69);
   U5 : BUF_X1 port map( A => rst, Z => n70);
   U6 : AND2_X1 port map( A1 => d_in(0), A2 => n68, ZN => N2);
   U7 : AND2_X1 port map( A1 => d_in(1), A2 => n69, ZN => N3);
   U8 : AND2_X1 port map( A1 => d_in(8), A2 => n68, ZN => N10);
   U9 : AND2_X1 port map( A1 => d_in(9), A2 => n68, ZN => N11);
   U10 : AND2_X1 port map( A1 => d_in(10), A2 => n68, ZN => N12);
   U11 : AND2_X1 port map( A1 => d_in(11), A2 => n68, ZN => N13);
   U12 : AND2_X1 port map( A1 => d_in(12), A2 => n68, ZN => N14);
   U13 : AND2_X1 port map( A1 => d_in(13), A2 => n68, ZN => N15);
   U14 : AND2_X1 port map( A1 => d_in(14), A2 => n68, ZN => N16);
   U15 : AND2_X1 port map( A1 => d_in(15), A2 => n68, ZN => N17);
   U16 : AND2_X1 port map( A1 => d_in(16), A2 => n68, ZN => N18);
   U17 : AND2_X1 port map( A1 => d_in(17), A2 => n68, ZN => N19);
   U18 : AND2_X1 port map( A1 => d_in(18), A2 => n68, ZN => N20);
   U19 : AND2_X1 port map( A1 => d_in(19), A2 => n69, ZN => N21);
   U20 : AND2_X1 port map( A1 => d_in(20), A2 => n69, ZN => N22);
   U21 : AND2_X1 port map( A1 => d_in(21), A2 => n69, ZN => N23);
   U22 : AND2_X1 port map( A1 => d_in(22), A2 => n69, ZN => N24);
   U23 : AND2_X1 port map( A1 => d_in(23), A2 => n69, ZN => N25);
   U24 : AND2_X1 port map( A1 => d_in(24), A2 => n69, ZN => N26);
   U25 : AND2_X1 port map( A1 => d_in(25), A2 => n69, ZN => N27);
   U26 : AND2_X1 port map( A1 => d_in(26), A2 => n69, ZN => N28);
   U27 : AND2_X1 port map( A1 => d_in(27), A2 => n69, ZN => N29);
   U28 : AND2_X1 port map( A1 => d_in(28), A2 => n69, ZN => N30);
   U29 : AND2_X1 port map( A1 => d_in(29), A2 => n69, ZN => N31);
   U30 : AND2_X1 port map( A1 => n70, A2 => d_in(7), ZN => N9);
   U31 : AND2_X1 port map( A1 => d_in(2), A2 => n70, ZN => N4);
   U32 : AND2_X1 port map( A1 => d_in(3), A2 => n70, ZN => N5);
   U33 : AND2_X1 port map( A1 => d_in(4), A2 => n70, ZN => N6);
   U34 : AND2_X1 port map( A1 => d_in(5), A2 => n70, ZN => N7);
   U35 : AND2_X1 port map( A1 => d_in(6), A2 => n70, ZN => N8);
   U36 : AND2_X1 port map( A1 => d_in(30), A2 => n70, ZN => N32);
   U37 : AND2_X1 port map( A1 => d_in(31), A2 => n70, ZN => N33);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity cla_adder_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end cla_adder_N32;

architecture SYN_struct of cla_adder_N32 is

   component sum_generator_Nbits32_Nblocks8
      port( A, B : in std_logic_vector (31 downto 0);  Carry : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_Nblocks8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal Carry_8_port, Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port,
      Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port : std_logic;

begin
   
   CG : carry_generator_N32_Nblocks8 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci, Cout(8) => 
                           Carry_8_port, Cout(7) => Carry_7_port, Cout(6) => 
                           Carry_6_port, Cout(5) => Carry_5_port, Cout(4) => 
                           Carry_4_port, Cout(3) => Carry_3_port, Cout(2) => 
                           Carry_2_port, Cout(1) => Carry_1_port, Cout(0) => 
                           Carry_0_port);
   SG : sum_generator_Nbits32_Nblocks8 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Carry(8) => Carry_8_port, 
                           Carry(7) => Carry_7_port, Carry(6) => Carry_6_port, 
                           Carry(5) => Carry_5_port, Carry(4) => Carry_4_port, 
                           Carry(3) => Carry_3_port, Carry(2) => Carry_2_port, 
                           Carry(1) => Carry_1_port, Carry(0) => Carry_0_port, 
                           S(31) => Sum(31), S(30) => Sum(30), S(29) => Sum(29)
                           , S(28) => Sum(28), S(27) => Sum(27), S(26) => 
                           Sum(26), S(25) => Sum(25), S(24) => Sum(24), S(23) 
                           => Sum(23), S(22) => Sum(22), S(21) => Sum(21), 
                           S(20) => Sum(20), S(19) => Sum(19), S(18) => Sum(18)
                           , S(17) => Sum(17), S(16) => Sum(16), S(15) => 
                           Sum(15), S(14) => Sum(14), S(13) => Sum(13), S(12) 
                           => Sum(12), S(11) => Sum(11), S(10) => Sum(10), S(9)
                           => Sum(9), S(8) => Sum(8), S(7) => Sum(7), S(6) => 
                           Sum(6), S(5) => Sum(5), S(4) => Sum(4), S(3) => 
                           Sum(3), S(2) => Sum(2), S(1) => Sum(1), S(0) => 
                           Sum(0), Cout => Cout);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity alu is

   port( A, B : in std_logic_vector (31 downto 0);  OP : in std_logic_vector (0
         to 4);  Y1 : out std_logic_vector (31 downto 0);  cout : out std_logic
         );

end alu;

architecture SYN_behav of alu is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component mux_alu
      port( addsub, mul, log, shift, lhi : in std_logic_vector (31 downto 0);  
            gt, get, lt, let, eq, neq : in std_logic;  sel : in 
            std_logic_vector (0 to 4);  out_mux : out std_logic_vector (31 
            downto 0));
   end component;
   
   component comparator
      port( C : in std_logic;  Sum : in std_logic_vector (31 downto 0);  sign :
            in std_logic;  gt, get, lt, let, eq, neq : out std_logic);
   end component;
   
   component shifter
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  C : out std_logic_vector (31 downto
            0));
   end component;
   
   component logical
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (3 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component booth_mul_N16
      port( A, B : in std_logic_vector (15 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component adder_sub_N32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, cout_port, add_sub, A_add_31_port, A_add_30_port, 
      A_add_29_port, A_add_28_port, A_add_27_port, A_add_26_port, A_add_25_port
      , A_add_24_port, A_add_23_port, A_add_22_port, A_add_21_port, 
      A_add_20_port, A_add_19_port, A_add_18_port, A_add_17_port, A_add_16_port
      , A_add_15_port, A_add_14_port, A_add_13_port, A_add_12_port, 
      A_add_11_port, A_add_10_port, A_add_9_port, A_add_8_port, A_add_7_port, 
      A_add_6_port, A_add_5_port, A_add_4_port, A_add_3_port, A_add_2_port, 
      A_add_1_port, A_add_0_port, B_add_31_port, B_add_30_port, B_add_29_port, 
      B_add_28_port, B_add_27_port, B_add_26_port, B_add_25_port, B_add_24_port
      , B_add_23_port, B_add_22_port, B_add_21_port, B_add_20_port, 
      B_add_19_port, B_add_18_port, B_add_17_port, B_add_16_port, B_add_15_port
      , B_add_14_port, B_add_13_port, B_add_12_port, B_add_11_port, 
      B_add_10_port, B_add_9_port, B_add_8_port, B_add_7_port, B_add_6_port, 
      B_add_5_port, B_add_4_port, B_add_3_port, B_add_2_port, B_add_1_port, 
      B_add_0_port, A_mul_15_port, A_mul_14_port, A_mul_13_port, A_mul_12_port,
      A_mul_11_port, A_mul_10_port, A_mul_9_port, A_mul_8_port, A_mul_7_port, 
      A_mul_6_port, A_mul_5_port, A_mul_4_port, A_mul_3_port, A_mul_2_port, 
      A_mul_1_port, B_mul_15_port, B_mul_14_port, B_mul_13_port, B_mul_12_port,
      B_mul_11_port, B_mul_10_port, B_mul_9_port, B_mul_8_port, B_mul_7_port, 
      B_mul_6_port, B_mul_5_port, B_mul_4_port, B_mul_3_port, B_mul_2_port, 
      B_mul_1_port, B_mul_0_port, sel_log_3_port, sel_log_2_port, 
      sel_log_1_port, sel_log_0_port, A_log_31_port, A_log_30_port, 
      A_log_29_port, A_log_28_port, A_log_27_port, A_log_26_port, A_log_25_port
      , A_log_24_port, A_log_23_port, A_log_22_port, A_log_21_port, 
      A_log_20_port, A_log_19_port, A_log_18_port, A_log_17_port, A_log_16_port
      , A_log_15_port, A_log_14_port, A_log_13_port, A_log_12_port, 
      A_log_11_port, A_log_10_port, A_log_9_port, A_log_8_port, A_log_7_port, 
      A_log_6_port, A_log_5_port, A_log_4_port, A_log_3_port, A_log_2_port, 
      A_log_1_port, A_log_0_port, B_log_31_port, B_log_30_port, B_log_29_port, 
      B_log_28_port, B_log_27_port, B_log_26_port, B_log_25_port, B_log_24_port
      , B_log_23_port, B_log_22_port, B_log_21_port, B_log_20_port, 
      B_log_19_port, B_log_18_port, B_log_17_port, B_log_16_port, B_log_15_port
      , B_log_14_port, B_log_13_port, B_log_12_port, B_log_11_port, 
      B_log_10_port, B_log_9_port, B_log_8_port, B_log_7_port, B_log_6_port, 
      B_log_5_port, B_log_4_port, B_log_3_port, B_log_2_port, B_log_1_port, 
      B_log_0_port, sel_shift_1_port, sel_shift_0_port, A_sht_31_port, 
      A_sht_30_port, A_sht_29_port, A_sht_28_port, A_sht_27_port, A_sht_26_port
      , A_sht_25_port, A_sht_24_port, A_sht_23_port, A_sht_22_port, 
      A_sht_21_port, A_sht_20_port, A_sht_19_port, A_sht_18_port, A_sht_17_port
      , A_sht_16_port, A_sht_15_port, A_sht_14_port, A_sht_13_port, 
      A_sht_12_port, A_sht_11_port, A_sht_10_port, A_sht_9_port, A_sht_8_port, 
      A_sht_7_port, A_sht_6_port, A_sht_5_port, A_sht_4_port, A_sht_3_port, 
      A_sht_2_port, A_sht_1_port, A_sht_0_port, B_sht_31_port, B_sht_30_port, 
      B_sht_29_port, B_sht_28_port, B_sht_27_port, B_sht_26_port, B_sht_25_port
      , B_sht_24_port, B_sht_23_port, B_sht_22_port, B_sht_21_port, 
      B_sht_20_port, B_sht_19_port, B_sht_18_port, B_sht_17_port, B_sht_16_port
      , B_sht_15_port, B_sht_14_port, B_sht_13_port, B_sht_12_port, 
      B_sht_11_port, B_sht_10_port, B_sht_9_port, B_sht_8_port, B_sht_7_port, 
      B_sht_6_port, B_sht_5_port, B_sht_4_port, B_sht_3_port, B_sht_2_port, 
      B_sht_1_port, B_sht_0_port, sign, B_lhi_15_port, B_lhi_14_port, 
      B_lhi_13_port, B_lhi_12_port, B_lhi_11_port, B_lhi_10_port, B_lhi_9_port,
      B_lhi_8_port, B_lhi_7_port, B_lhi_6_port, B_lhi_5_port, B_lhi_4_port, 
      B_lhi_3_port, B_lhi_2_port, B_lhi_1_port, B_lhi_0_port, N25, N26, N27, 
      N28, N29, N31, N32, N33, N34, N35, N36, out_add_31_port, out_add_30_port,
      out_add_29_port, out_add_28_port, out_add_27_port, out_add_26_port, 
      out_add_25_port, out_add_24_port, out_add_23_port, out_add_22_port, 
      out_add_21_port, out_add_20_port, out_add_19_port, out_add_18_port, 
      out_add_17_port, out_add_16_port, out_add_15_port, out_add_14_port, 
      out_add_13_port, out_add_12_port, out_add_11_port, out_add_10_port, 
      out_add_9_port, out_add_8_port, out_add_7_port, out_add_6_port, 
      out_add_5_port, out_add_4_port, out_add_3_port, out_add_2_port, 
      out_add_1_port, out_add_0_port, out_mul_31_port, out_mul_30_port, 
      out_mul_29_port, out_mul_28_port, out_mul_27_port, out_mul_26_port, 
      out_mul_25_port, out_mul_24_port, out_mul_23_port, out_mul_22_port, 
      out_mul_21_port, out_mul_20_port, out_mul_19_port, out_mul_18_port, 
      out_mul_17_port, out_mul_16_port, out_mul_15_port, out_mul_14_port, 
      out_mul_13_port, out_mul_12_port, out_mul_11_port, out_mul_10_port, 
      out_mul_9_port, out_mul_8_port, out_mul_7_port, out_mul_6_port, 
      out_mul_5_port, out_mul_4_port, out_mul_3_port, out_mul_2_port, 
      out_mul_1_port, out_mul_0_port, out_log_31_port, out_log_30_port, 
      out_log_29_port, out_log_28_port, out_log_27_port, out_log_26_port, 
      out_log_25_port, out_log_24_port, out_log_23_port, out_log_22_port, 
      out_log_21_port, out_log_20_port, out_log_19_port, out_log_18_port, 
      out_log_17_port, out_log_16_port, out_log_15_port, out_log_14_port, 
      out_log_13_port, out_log_12_port, out_log_11_port, out_log_10_port, 
      out_log_9_port, out_log_8_port, out_log_7_port, out_log_6_port, 
      out_log_5_port, out_log_4_port, out_log_3_port, out_log_2_port, 
      out_log_1_port, out_log_0_port, out_shift_31_port, out_shift_30_port, 
      out_shift_29_port, out_shift_28_port, out_shift_27_port, 
      out_shift_26_port, out_shift_25_port, out_shift_24_port, 
      out_shift_23_port, out_shift_22_port, out_shift_21_port, 
      out_shift_20_port, out_shift_19_port, out_shift_18_port, 
      out_shift_17_port, out_shift_16_port, out_shift_15_port, 
      out_shift_14_port, out_shift_13_port, out_shift_12_port, 
      out_shift_11_port, out_shift_10_port, out_shift_9_port, out_shift_8_port,
      out_shift_7_port, out_shift_6_port, out_shift_5_port, out_shift_4_port, 
      out_shift_3_port, out_shift_2_port, out_shift_1_port, out_shift_0_port, 
      gt, get, lt, let, eq, neq, n23, n24, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98 : std_logic;

begin
   cout <= cout_port;
   
   adder_subtr : adder_sub_N32 port map( A(31) => A_add_31_port, A(30) => 
                           A_add_30_port, A(29) => A_add_29_port, A(28) => 
                           A_add_28_port, A(27) => A_add_27_port, A(26) => 
                           A_add_26_port, A(25) => A_add_25_port, A(24) => 
                           A_add_24_port, A(23) => A_add_23_port, A(22) => 
                           A_add_22_port, A(21) => A_add_21_port, A(20) => 
                           A_add_20_port, A(19) => A_add_19_port, A(18) => 
                           A_add_18_port, A(17) => A_add_17_port, A(16) => 
                           A_add_16_port, A(15) => A_add_15_port, A(14) => 
                           A_add_14_port, A(13) => A_add_13_port, A(12) => 
                           A_add_12_port, A(11) => A_add_11_port, A(10) => 
                           A_add_10_port, A(9) => A_add_9_port, A(8) => 
                           A_add_8_port, A(7) => A_add_7_port, A(6) => 
                           A_add_6_port, A(5) => A_add_5_port, A(4) => 
                           A_add_4_port, A(3) => A_add_3_port, A(2) => 
                           A_add_2_port, A(1) => A_add_1_port, A(0) => 
                           A_add_0_port, B(31) => B_add_31_port, B(30) => 
                           B_add_30_port, B(29) => B_add_29_port, B(28) => 
                           B_add_28_port, B(27) => B_add_27_port, B(26) => 
                           B_add_26_port, B(25) => B_add_25_port, B(24) => 
                           B_add_24_port, B(23) => B_add_23_port, B(22) => 
                           B_add_22_port, B(21) => B_add_21_port, B(20) => 
                           B_add_20_port, B(19) => B_add_19_port, B(18) => 
                           B_add_18_port, B(17) => B_add_17_port, B(16) => 
                           B_add_16_port, B(15) => B_add_15_port, B(14) => 
                           B_add_14_port, B(13) => B_add_13_port, B(12) => 
                           B_add_12_port, B(11) => B_add_11_port, B(10) => 
                           B_add_10_port, B(9) => B_add_9_port, B(8) => 
                           B_add_8_port, B(7) => B_add_7_port, B(6) => 
                           B_add_6_port, B(5) => B_add_5_port, B(4) => 
                           B_add_4_port, B(3) => B_add_3_port, B(2) => 
                           B_add_2_port, B(1) => B_add_1_port, B(0) => 
                           B_add_0_port, Ci => add_sub, Cout => cout_port, 
                           Sum(31) => out_add_31_port, Sum(30) => 
                           out_add_30_port, Sum(29) => out_add_29_port, Sum(28)
                           => out_add_28_port, Sum(27) => out_add_27_port, 
                           Sum(26) => out_add_26_port, Sum(25) => 
                           out_add_25_port, Sum(24) => out_add_24_port, Sum(23)
                           => out_add_23_port, Sum(22) => out_add_22_port, 
                           Sum(21) => out_add_21_port, Sum(20) => 
                           out_add_20_port, Sum(19) => out_add_19_port, Sum(18)
                           => out_add_18_port, Sum(17) => out_add_17_port, 
                           Sum(16) => out_add_16_port, Sum(15) => 
                           out_add_15_port, Sum(14) => out_add_14_port, Sum(13)
                           => out_add_13_port, Sum(12) => out_add_12_port, 
                           Sum(11) => out_add_11_port, Sum(10) => 
                           out_add_10_port, Sum(9) => out_add_9_port, Sum(8) =>
                           out_add_8_port, Sum(7) => out_add_7_port, Sum(6) => 
                           out_add_6_port, Sum(5) => out_add_5_port, Sum(4) => 
                           out_add_4_port, Sum(3) => out_add_3_port, Sum(2) => 
                           out_add_2_port, Sum(1) => out_add_1_port, Sum(0) => 
                           out_add_0_port);
   mul : booth_mul_N16 port map( A(15) => A_mul_15_port, A(14) => A_mul_14_port
                           , A(13) => A_mul_13_port, A(12) => A_mul_12_port, 
                           A(11) => A_mul_11_port, A(10) => A_mul_10_port, A(9)
                           => A_mul_9_port, A(8) => A_mul_8_port, A(7) => 
                           A_mul_7_port, A(6) => A_mul_6_port, A(5) => 
                           A_mul_5_port, A(4) => A_mul_4_port, A(3) => 
                           A_mul_3_port, A(2) => A_mul_2_port, A(1) => 
                           A_mul_1_port, A(0) => n23, B(15) => B_mul_15_port, 
                           B(14) => B_mul_14_port, B(13) => B_mul_13_port, 
                           B(12) => B_mul_12_port, B(11) => B_mul_11_port, 
                           B(10) => B_mul_10_port, B(9) => B_mul_9_port, B(8) 
                           => B_mul_8_port, B(7) => B_mul_7_port, B(6) => 
                           B_mul_6_port, B(5) => B_mul_5_port, B(4) => 
                           B_mul_4_port, B(3) => B_mul_3_port, B(2) => 
                           B_mul_2_port, B(1) => B_mul_1_port, B(0) => 
                           B_mul_0_port, Y(31) => out_mul_31_port, Y(30) => 
                           out_mul_30_port, Y(29) => out_mul_29_port, Y(28) => 
                           out_mul_28_port, Y(27) => out_mul_27_port, Y(26) => 
                           out_mul_26_port, Y(25) => out_mul_25_port, Y(24) => 
                           out_mul_24_port, Y(23) => out_mul_23_port, Y(22) => 
                           out_mul_22_port, Y(21) => out_mul_21_port, Y(20) => 
                           out_mul_20_port, Y(19) => out_mul_19_port, Y(18) => 
                           out_mul_18_port, Y(17) => out_mul_17_port, Y(16) => 
                           out_mul_16_port, Y(15) => out_mul_15_port, Y(14) => 
                           out_mul_14_port, Y(13) => out_mul_13_port, Y(12) => 
                           out_mul_12_port, Y(11) => out_mul_11_port, Y(10) => 
                           out_mul_10_port, Y(9) => out_mul_9_port, Y(8) => 
                           out_mul_8_port, Y(7) => out_mul_7_port, Y(6) => 
                           out_mul_6_port, Y(5) => out_mul_5_port, Y(4) => 
                           out_mul_4_port, Y(3) => out_mul_3_port, Y(2) => 
                           out_mul_2_port, Y(1) => out_mul_1_port, Y(0) => 
                           out_mul_0_port);
   logic : logical port map( A(31) => A_log_31_port, A(30) => A_log_30_port, 
                           A(29) => A_log_29_port, A(28) => A_log_28_port, 
                           A(27) => A_log_27_port, A(26) => A_log_26_port, 
                           A(25) => A_log_25_port, A(24) => A_log_24_port, 
                           A(23) => A_log_23_port, A(22) => A_log_22_port, 
                           A(21) => A_log_21_port, A(20) => A_log_20_port, 
                           A(19) => A_log_19_port, A(18) => A_log_18_port, 
                           A(17) => A_log_17_port, A(16) => A_log_16_port, 
                           A(15) => A_log_15_port, A(14) => A_log_14_port, 
                           A(13) => A_log_13_port, A(12) => A_log_12_port, 
                           A(11) => A_log_11_port, A(10) => A_log_10_port, A(9)
                           => A_log_9_port, A(8) => A_log_8_port, A(7) => 
                           A_log_7_port, A(6) => A_log_6_port, A(5) => 
                           A_log_5_port, A(4) => A_log_4_port, A(3) => 
                           A_log_3_port, A(2) => A_log_2_port, A(1) => 
                           A_log_1_port, A(0) => A_log_0_port, B(31) => 
                           B_log_31_port, B(30) => B_log_30_port, B(29) => 
                           B_log_29_port, B(28) => B_log_28_port, B(27) => 
                           B_log_27_port, B(26) => B_log_26_port, B(25) => 
                           B_log_25_port, B(24) => B_log_24_port, B(23) => 
                           B_log_23_port, B(22) => B_log_22_port, B(21) => 
                           B_log_21_port, B(20) => B_log_20_port, B(19) => 
                           B_log_19_port, B(18) => B_log_18_port, B(17) => 
                           B_log_17_port, B(16) => B_log_16_port, B(15) => 
                           B_log_15_port, B(14) => B_log_14_port, B(13) => 
                           B_log_13_port, B(12) => B_log_12_port, B(11) => 
                           B_log_11_port, B(10) => B_log_10_port, B(9) => 
                           B_log_9_port, B(8) => B_log_8_port, B(7) => 
                           B_log_7_port, B(6) => B_log_6_port, B(5) => 
                           B_log_5_port, B(4) => B_log_4_port, B(3) => 
                           B_log_3_port, B(2) => B_log_2_port, B(1) => 
                           B_log_1_port, B(0) => B_log_0_port, sel(3) => 
                           sel_log_3_port, sel(2) => sel_log_2_port, sel(1) => 
                           sel_log_1_port, sel(0) => sel_log_0_port, Y(31) => 
                           out_log_31_port, Y(30) => out_log_30_port, Y(29) => 
                           out_log_29_port, Y(28) => out_log_28_port, Y(27) => 
                           out_log_27_port, Y(26) => out_log_26_port, Y(25) => 
                           out_log_25_port, Y(24) => out_log_24_port, Y(23) => 
                           out_log_23_port, Y(22) => out_log_22_port, Y(21) => 
                           out_log_21_port, Y(20) => out_log_20_port, Y(19) => 
                           out_log_19_port, Y(18) => out_log_18_port, Y(17) => 
                           out_log_17_port, Y(16) => out_log_16_port, Y(15) => 
                           out_log_15_port, Y(14) => out_log_14_port, Y(13) => 
                           out_log_13_port, Y(12) => out_log_12_port, Y(11) => 
                           out_log_11_port, Y(10) => out_log_10_port, Y(9) => 
                           out_log_9_port, Y(8) => out_log_8_port, Y(7) => 
                           out_log_7_port, Y(6) => out_log_6_port, Y(5) => 
                           out_log_5_port, Y(4) => out_log_4_port, Y(3) => 
                           out_log_3_port, Y(2) => out_log_2_port, Y(1) => 
                           out_log_1_port, Y(0) => out_log_0_port);
   shift : shifter port map( A(31) => A_sht_31_port, A(30) => A_sht_30_port, 
                           A(29) => A_sht_29_port, A(28) => A_sht_28_port, 
                           A(27) => A_sht_27_port, A(26) => A_sht_26_port, 
                           A(25) => A_sht_25_port, A(24) => A_sht_24_port, 
                           A(23) => A_sht_23_port, A(22) => A_sht_22_port, 
                           A(21) => A_sht_21_port, A(20) => A_sht_20_port, 
                           A(19) => A_sht_19_port, A(18) => A_sht_18_port, 
                           A(17) => A_sht_17_port, A(16) => A_sht_16_port, 
                           A(15) => A_sht_15_port, A(14) => A_sht_14_port, 
                           A(13) => A_sht_13_port, A(12) => A_sht_12_port, 
                           A(11) => A_sht_11_port, A(10) => A_sht_10_port, A(9)
                           => A_sht_9_port, A(8) => A_sht_8_port, A(7) => 
                           A_sht_7_port, A(6) => A_sht_6_port, A(5) => 
                           A_sht_5_port, A(4) => A_sht_4_port, A(3) => 
                           A_sht_3_port, A(2) => A_sht_2_port, A(1) => 
                           A_sht_1_port, A(0) => A_sht_0_port, B(31) => 
                           B_sht_31_port, B(30) => B_sht_30_port, B(29) => 
                           B_sht_29_port, B(28) => B_sht_28_port, B(27) => 
                           B_sht_27_port, B(26) => B_sht_26_port, B(25) => 
                           B_sht_25_port, B(24) => B_sht_24_port, B(23) => 
                           B_sht_23_port, B(22) => B_sht_22_port, B(21) => 
                           B_sht_21_port, B(20) => B_sht_20_port, B(19) => 
                           B_sht_19_port, B(18) => B_sht_18_port, B(17) => 
                           B_sht_17_port, B(16) => B_sht_16_port, B(15) => 
                           B_sht_15_port, B(14) => B_sht_14_port, B(13) => 
                           B_sht_13_port, B(12) => B_sht_12_port, B(11) => 
                           B_sht_11_port, B(10) => B_sht_10_port, B(9) => 
                           B_sht_9_port, B(8) => B_sht_8_port, B(7) => 
                           B_sht_7_port, B(6) => B_sht_6_port, B(5) => 
                           B_sht_5_port, B(4) => B_sht_4_port, B(3) => 
                           B_sht_3_port, B(2) => B_sht_2_port, B(1) => 
                           B_sht_1_port, B(0) => B_sht_0_port, sel(1) => 
                           sel_shift_1_port, sel(0) => sel_shift_0_port, C(31) 
                           => out_shift_31_port, C(30) => out_shift_30_port, 
                           C(29) => out_shift_29_port, C(28) => 
                           out_shift_28_port, C(27) => out_shift_27_port, C(26)
                           => out_shift_26_port, C(25) => out_shift_25_port, 
                           C(24) => out_shift_24_port, C(23) => 
                           out_shift_23_port, C(22) => out_shift_22_port, C(21)
                           => out_shift_21_port, C(20) => out_shift_20_port, 
                           C(19) => out_shift_19_port, C(18) => 
                           out_shift_18_port, C(17) => out_shift_17_port, C(16)
                           => out_shift_16_port, C(15) => out_shift_15_port, 
                           C(14) => out_shift_14_port, C(13) => 
                           out_shift_13_port, C(12) => out_shift_12_port, C(11)
                           => out_shift_11_port, C(10) => out_shift_10_port, 
                           C(9) => out_shift_9_port, C(8) => out_shift_8_port, 
                           C(7) => out_shift_7_port, C(6) => out_shift_6_port, 
                           C(5) => out_shift_5_port, C(4) => out_shift_4_port, 
                           C(3) => out_shift_3_port, C(2) => out_shift_2_port, 
                           C(1) => out_shift_1_port, C(0) => out_shift_0_port);
   compar : comparator port map( C => cout_port, Sum(31) => out_add_31_port, 
                           Sum(30) => out_add_30_port, Sum(29) => 
                           out_add_29_port, Sum(28) => out_add_28_port, Sum(27)
                           => out_add_27_port, Sum(26) => out_add_26_port, 
                           Sum(25) => out_add_25_port, Sum(24) => 
                           out_add_24_port, Sum(23) => out_add_23_port, Sum(22)
                           => out_add_22_port, Sum(21) => out_add_21_port, 
                           Sum(20) => out_add_20_port, Sum(19) => 
                           out_add_19_port, Sum(18) => out_add_18_port, Sum(17)
                           => out_add_17_port, Sum(16) => out_add_16_port, 
                           Sum(15) => out_add_15_port, Sum(14) => 
                           out_add_14_port, Sum(13) => out_add_13_port, Sum(12)
                           => out_add_12_port, Sum(11) => out_add_11_port, 
                           Sum(10) => out_add_10_port, Sum(9) => out_add_9_port
                           , Sum(8) => out_add_8_port, Sum(7) => out_add_7_port
                           , Sum(6) => out_add_6_port, Sum(5) => out_add_5_port
                           , Sum(4) => out_add_4_port, Sum(3) => out_add_3_port
                           , Sum(2) => out_add_2_port, Sum(1) => out_add_1_port
                           , Sum(0) => out_add_0_port, sign => sign, gt => gt, 
                           get => get, lt => lt, let => let, eq => eq, neq => 
                           neq);
   muxy1 : mux_alu port map( addsub(31) => out_add_31_port, addsub(30) => 
                           out_add_30_port, addsub(29) => out_add_29_port, 
                           addsub(28) => out_add_28_port, addsub(27) => 
                           out_add_27_port, addsub(26) => out_add_26_port, 
                           addsub(25) => out_add_25_port, addsub(24) => 
                           out_add_24_port, addsub(23) => out_add_23_port, 
                           addsub(22) => out_add_22_port, addsub(21) => 
                           out_add_21_port, addsub(20) => out_add_20_port, 
                           addsub(19) => out_add_19_port, addsub(18) => 
                           out_add_18_port, addsub(17) => out_add_17_port, 
                           addsub(16) => out_add_16_port, addsub(15) => 
                           out_add_15_port, addsub(14) => out_add_14_port, 
                           addsub(13) => out_add_13_port, addsub(12) => 
                           out_add_12_port, addsub(11) => out_add_11_port, 
                           addsub(10) => out_add_10_port, addsub(9) => 
                           out_add_9_port, addsub(8) => out_add_8_port, 
                           addsub(7) => out_add_7_port, addsub(6) => 
                           out_add_6_port, addsub(5) => out_add_5_port, 
                           addsub(4) => out_add_4_port, addsub(3) => 
                           out_add_3_port, addsub(2) => out_add_2_port, 
                           addsub(1) => out_add_1_port, addsub(0) => 
                           out_add_0_port, mul(31) => out_mul_31_port, mul(30) 
                           => out_mul_30_port, mul(29) => out_mul_29_port, 
                           mul(28) => out_mul_28_port, mul(27) => 
                           out_mul_27_port, mul(26) => out_mul_26_port, mul(25)
                           => out_mul_25_port, mul(24) => out_mul_24_port, 
                           mul(23) => out_mul_23_port, mul(22) => 
                           out_mul_22_port, mul(21) => out_mul_21_port, mul(20)
                           => out_mul_20_port, mul(19) => out_mul_19_port, 
                           mul(18) => out_mul_18_port, mul(17) => 
                           out_mul_17_port, mul(16) => out_mul_16_port, mul(15)
                           => out_mul_15_port, mul(14) => out_mul_14_port, 
                           mul(13) => out_mul_13_port, mul(12) => 
                           out_mul_12_port, mul(11) => out_mul_11_port, mul(10)
                           => out_mul_10_port, mul(9) => out_mul_9_port, mul(8)
                           => out_mul_8_port, mul(7) => out_mul_7_port, mul(6) 
                           => out_mul_6_port, mul(5) => out_mul_5_port, mul(4) 
                           => out_mul_4_port, mul(3) => out_mul_3_port, mul(2) 
                           => out_mul_2_port, mul(1) => out_mul_1_port, mul(0) 
                           => out_mul_0_port, log(31) => out_log_31_port, 
                           log(30) => out_log_30_port, log(29) => 
                           out_log_29_port, log(28) => out_log_28_port, log(27)
                           => out_log_27_port, log(26) => out_log_26_port, 
                           log(25) => out_log_25_port, log(24) => 
                           out_log_24_port, log(23) => out_log_23_port, log(22)
                           => out_log_22_port, log(21) => out_log_21_port, 
                           log(20) => out_log_20_port, log(19) => 
                           out_log_19_port, log(18) => out_log_18_port, log(17)
                           => out_log_17_port, log(16) => out_log_16_port, 
                           log(15) => out_log_15_port, log(14) => 
                           out_log_14_port, log(13) => out_log_13_port, log(12)
                           => out_log_12_port, log(11) => out_log_11_port, 
                           log(10) => out_log_10_port, log(9) => out_log_9_port
                           , log(8) => out_log_8_port, log(7) => out_log_7_port
                           , log(6) => out_log_6_port, log(5) => out_log_5_port
                           , log(4) => out_log_4_port, log(3) => out_log_3_port
                           , log(2) => out_log_2_port, log(1) => out_log_1_port
                           , log(0) => out_log_0_port, shift(31) => 
                           out_shift_31_port, shift(30) => out_shift_30_port, 
                           shift(29) => out_shift_29_port, shift(28) => 
                           out_shift_28_port, shift(27) => out_shift_27_port, 
                           shift(26) => out_shift_26_port, shift(25) => 
                           out_shift_25_port, shift(24) => out_shift_24_port, 
                           shift(23) => out_shift_23_port, shift(22) => 
                           out_shift_22_port, shift(21) => out_shift_21_port, 
                           shift(20) => out_shift_20_port, shift(19) => 
                           out_shift_19_port, shift(18) => out_shift_18_port, 
                           shift(17) => out_shift_17_port, shift(16) => 
                           out_shift_16_port, shift(15) => out_shift_15_port, 
                           shift(14) => out_shift_14_port, shift(13) => 
                           out_shift_13_port, shift(12) => out_shift_12_port, 
                           shift(11) => out_shift_11_port, shift(10) => 
                           out_shift_10_port, shift(9) => out_shift_9_port, 
                           shift(8) => out_shift_8_port, shift(7) => 
                           out_shift_7_port, shift(6) => out_shift_6_port, 
                           shift(5) => out_shift_5_port, shift(4) => 
                           out_shift_4_port, shift(3) => out_shift_3_port, 
                           shift(2) => out_shift_2_port, shift(1) => 
                           out_shift_1_port, shift(0) => out_shift_0_port, 
                           lhi(31) => B_lhi_15_port, lhi(30) => B_lhi_14_port, 
                           lhi(29) => B_lhi_13_port, lhi(28) => B_lhi_12_port, 
                           lhi(27) => B_lhi_11_port, lhi(26) => B_lhi_10_port, 
                           lhi(25) => B_lhi_9_port, lhi(24) => B_lhi_8_port, 
                           lhi(23) => B_lhi_7_port, lhi(22) => B_lhi_6_port, 
                           lhi(21) => B_lhi_5_port, lhi(20) => B_lhi_4_port, 
                           lhi(19) => B_lhi_3_port, lhi(18) => B_lhi_2_port, 
                           lhi(17) => B_lhi_1_port, lhi(16) => B_lhi_0_port, 
                           lhi(15) => X_Logic0_port, lhi(14) => X_Logic0_port, 
                           lhi(13) => X_Logic0_port, lhi(12) => X_Logic0_port, 
                           lhi(11) => X_Logic0_port, lhi(10) => X_Logic0_port, 
                           lhi(9) => X_Logic0_port, lhi(8) => X_Logic0_port, 
                           lhi(7) => X_Logic0_port, lhi(6) => X_Logic0_port, 
                           lhi(5) => X_Logic0_port, lhi(4) => X_Logic0_port, 
                           lhi(3) => X_Logic0_port, lhi(2) => X_Logic0_port, 
                           lhi(1) => X_Logic0_port, lhi(0) => X_Logic0_port, gt
                           => gt, get => get, lt => lt, let => let, eq => eq, 
                           neq => neq, sel(0) => OP(0), sel(1) => OP(1), sel(2)
                           => OP(2), sel(3) => OP(3), sel(4) => OP(4), 
                           out_mux(31) => Y1(31), out_mux(30) => Y1(30), 
                           out_mux(29) => Y1(29), out_mux(28) => Y1(28), 
                           out_mux(27) => Y1(27), out_mux(26) => Y1(26), 
                           out_mux(25) => Y1(25), out_mux(24) => Y1(24), 
                           out_mux(23) => Y1(23), out_mux(22) => Y1(22), 
                           out_mux(21) => Y1(21), out_mux(20) => Y1(20), 
                           out_mux(19) => Y1(19), out_mux(18) => Y1(18), 
                           out_mux(17) => Y1(17), out_mux(16) => Y1(16), 
                           out_mux(15) => Y1(15), out_mux(14) => Y1(14), 
                           out_mux(13) => Y1(13), out_mux(12) => Y1(12), 
                           out_mux(11) => Y1(11), out_mux(10) => Y1(10), 
                           out_mux(9) => Y1(9), out_mux(8) => Y1(8), out_mux(7)
                           => Y1(7), out_mux(6) => Y1(6), out_mux(5) => Y1(5), 
                           out_mux(4) => Y1(4), out_mux(3) => Y1(3), out_mux(2)
                           => Y1(2), out_mux(1) => Y1(1), out_mux(0) => Y1(0));
   X_Logic0_port <= '0';
   B_lhi_reg_15_inst : DLH_X1 port map( G => N36, D => B(15), Q => 
                           B_lhi_15_port);
   B_lhi_reg_14_inst : DLH_X1 port map( G => N36, D => B(14), Q => 
                           B_lhi_14_port);
   B_lhi_reg_13_inst : DLH_X1 port map( G => N36, D => B(13), Q => 
                           B_lhi_13_port);
   B_lhi_reg_12_inst : DLH_X1 port map( G => N36, D => B(12), Q => 
                           B_lhi_12_port);
   B_lhi_reg_11_inst : DLH_X1 port map( G => N36, D => B(11), Q => 
                           B_lhi_11_port);
   B_lhi_reg_10_inst : DLH_X1 port map( G => N36, D => B(10), Q => 
                           B_lhi_10_port);
   B_lhi_reg_9_inst : DLH_X1 port map( G => N36, D => B(9), Q => B_lhi_9_port);
   B_lhi_reg_8_inst : DLH_X1 port map( G => N36, D => B(8), Q => B_lhi_8_port);
   B_lhi_reg_7_inst : DLH_X1 port map( G => N36, D => B(7), Q => B_lhi_7_port);
   B_lhi_reg_6_inst : DLH_X1 port map( G => N36, D => B(6), Q => B_lhi_6_port);
   B_lhi_reg_5_inst : DLH_X1 port map( G => N36, D => B(5), Q => B_lhi_5_port);
   B_lhi_reg_4_inst : DLH_X1 port map( G => N36, D => B(4), Q => B_lhi_4_port);
   B_lhi_reg_3_inst : DLH_X1 port map( G => N36, D => B(3), Q => B_lhi_3_port);
   B_lhi_reg_2_inst : DLH_X1 port map( G => N36, D => B(2), Q => B_lhi_2_port);
   B_lhi_reg_1_inst : DLH_X1 port map( G => N36, D => B(1), Q => B_lhi_1_port);
   B_lhi_reg_0_inst : DLH_X1 port map( G => N36, D => B(0), Q => B_lhi_0_port);
   A_add_reg_31_inst : DLH_X1 port map( G => n98, D => A(31), Q => 
                           A_add_31_port);
   A_add_reg_30_inst : DLH_X1 port map( G => n98, D => A(30), Q => 
                           A_add_30_port);
   A_add_reg_29_inst : DLH_X1 port map( G => n98, D => A(29), Q => 
                           A_add_29_port);
   A_add_reg_28_inst : DLH_X1 port map( G => n98, D => A(28), Q => 
                           A_add_28_port);
   A_add_reg_27_inst : DLH_X1 port map( G => n98, D => A(27), Q => 
                           A_add_27_port);
   A_add_reg_26_inst : DLH_X1 port map( G => n98, D => A(26), Q => 
                           A_add_26_port);
   A_add_reg_25_inst : DLH_X1 port map( G => n98, D => A(25), Q => 
                           A_add_25_port);
   A_add_reg_24_inst : DLH_X1 port map( G => n98, D => A(24), Q => 
                           A_add_24_port);
   A_add_reg_23_inst : DLH_X1 port map( G => n98, D => A(23), Q => 
                           A_add_23_port);
   A_add_reg_22_inst : DLH_X1 port map( G => n98, D => A(22), Q => 
                           A_add_22_port);
   A_add_reg_21_inst : DLH_X1 port map( G => n97, D => A(21), Q => 
                           A_add_21_port);
   A_add_reg_20_inst : DLH_X1 port map( G => n97, D => A(20), Q => 
                           A_add_20_port);
   A_add_reg_19_inst : DLH_X1 port map( G => n97, D => A(19), Q => 
                           A_add_19_port);
   A_add_reg_18_inst : DLH_X1 port map( G => n97, D => A(18), Q => 
                           A_add_18_port);
   A_add_reg_17_inst : DLH_X1 port map( G => n97, D => A(17), Q => 
                           A_add_17_port);
   A_add_reg_16_inst : DLH_X1 port map( G => n97, D => A(16), Q => 
                           A_add_16_port);
   A_add_reg_15_inst : DLH_X1 port map( G => n97, D => A(15), Q => 
                           A_add_15_port);
   A_add_reg_14_inst : DLH_X1 port map( G => n97, D => A(14), Q => 
                           A_add_14_port);
   A_add_reg_13_inst : DLH_X1 port map( G => n97, D => A(13), Q => 
                           A_add_13_port);
   A_add_reg_12_inst : DLH_X1 port map( G => n97, D => A(12), Q => 
                           A_add_12_port);
   A_add_reg_11_inst : DLH_X1 port map( G => n97, D => A(11), Q => 
                           A_add_11_port);
   A_add_reg_10_inst : DLH_X1 port map( G => n96, D => A(10), Q => 
                           A_add_10_port);
   A_add_reg_9_inst : DLH_X1 port map( G => n96, D => A(9), Q => A_add_9_port);
   A_add_reg_8_inst : DLH_X1 port map( G => n96, D => A(8), Q => A_add_8_port);
   A_add_reg_7_inst : DLH_X1 port map( G => n96, D => A(7), Q => A_add_7_port);
   A_add_reg_6_inst : DLH_X1 port map( G => n96, D => A(6), Q => A_add_6_port);
   A_add_reg_5_inst : DLH_X1 port map( G => n96, D => A(5), Q => A_add_5_port);
   A_add_reg_4_inst : DLH_X1 port map( G => n96, D => A(4), Q => A_add_4_port);
   A_add_reg_3_inst : DLH_X1 port map( G => n96, D => A(3), Q => A_add_3_port);
   A_add_reg_2_inst : DLH_X1 port map( G => n96, D => A(2), Q => A_add_2_port);
   A_add_reg_1_inst : DLH_X1 port map( G => n96, D => A(1), Q => A_add_1_port);
   A_add_reg_0_inst : DLH_X1 port map( G => n96, D => A(0), Q => A_add_0_port);
   B_add_reg_31_inst : DLH_X1 port map( G => n95, D => B(31), Q => 
                           B_add_31_port);
   B_add_reg_30_inst : DLH_X1 port map( G => n95, D => B(30), Q => 
                           B_add_30_port);
   B_add_reg_29_inst : DLH_X1 port map( G => n95, D => B(29), Q => 
                           B_add_29_port);
   B_add_reg_28_inst : DLH_X1 port map( G => n95, D => B(28), Q => 
                           B_add_28_port);
   B_add_reg_27_inst : DLH_X1 port map( G => n95, D => B(27), Q => 
                           B_add_27_port);
   B_add_reg_26_inst : DLH_X1 port map( G => n95, D => B(26), Q => 
                           B_add_26_port);
   B_add_reg_25_inst : DLH_X1 port map( G => n95, D => B(25), Q => 
                           B_add_25_port);
   B_add_reg_24_inst : DLH_X1 port map( G => n95, D => B(24), Q => 
                           B_add_24_port);
   B_add_reg_23_inst : DLH_X1 port map( G => n95, D => B(23), Q => 
                           B_add_23_port);
   B_add_reg_22_inst : DLH_X1 port map( G => n95, D => B(22), Q => 
                           B_add_22_port);
   B_add_reg_21_inst : DLH_X1 port map( G => n95, D => B(21), Q => 
                           B_add_21_port);
   B_add_reg_20_inst : DLH_X1 port map( G => n94, D => B(20), Q => 
                           B_add_20_port);
   B_add_reg_19_inst : DLH_X1 port map( G => n94, D => B(19), Q => 
                           B_add_19_port);
   B_add_reg_18_inst : DLH_X1 port map( G => n94, D => B(18), Q => 
                           B_add_18_port);
   B_add_reg_17_inst : DLH_X1 port map( G => n94, D => B(17), Q => 
                           B_add_17_port);
   B_add_reg_16_inst : DLH_X1 port map( G => n94, D => B(16), Q => 
                           B_add_16_port);
   B_add_reg_15_inst : DLH_X1 port map( G => n94, D => B(15), Q => 
                           B_add_15_port);
   B_add_reg_14_inst : DLH_X1 port map( G => n94, D => B(14), Q => 
                           B_add_14_port);
   B_add_reg_13_inst : DLH_X1 port map( G => n94, D => B(13), Q => 
                           B_add_13_port);
   B_add_reg_12_inst : DLH_X1 port map( G => n94, D => B(12), Q => 
                           B_add_12_port);
   B_add_reg_11_inst : DLH_X1 port map( G => n94, D => B(11), Q => 
                           B_add_11_port);
   B_add_reg_10_inst : DLH_X1 port map( G => n94, D => B(10), Q => 
                           B_add_10_port);
   B_add_reg_9_inst : DLH_X1 port map( G => n93, D => B(9), Q => B_add_9_port);
   B_add_reg_8_inst : DLH_X1 port map( G => n93, D => B(8), Q => B_add_8_port);
   B_add_reg_7_inst : DLH_X1 port map( G => n93, D => B(7), Q => B_add_7_port);
   B_add_reg_6_inst : DLH_X1 port map( G => n93, D => B(6), Q => B_add_6_port);
   B_add_reg_5_inst : DLH_X1 port map( G => n93, D => B(5), Q => B_add_5_port);
   B_add_reg_4_inst : DLH_X1 port map( G => n93, D => B(4), Q => B_add_4_port);
   B_add_reg_3_inst : DLH_X1 port map( G => n93, D => B(3), Q => B_add_3_port);
   B_add_reg_2_inst : DLH_X1 port map( G => n93, D => B(2), Q => B_add_2_port);
   B_add_reg_1_inst : DLH_X1 port map( G => n93, D => B(1), Q => B_add_1_port);
   B_add_reg_0_inst : DLH_X1 port map( G => n93, D => B(0), Q => B_add_0_port);
   A_mul_reg_15_inst : DLH_X1 port map( G => n92, D => A(15), Q => 
                           A_mul_15_port);
   A_mul_reg_0_inst : DLH_X1 port map( G => n92, D => A(0), Q => n23);
   B_mul_reg_15_inst : DLH_X1 port map( G => n92, D => B(15), Q => 
                           B_mul_15_port);
   B_mul_reg_14_inst : DLH_X1 port map( G => n92, D => B(14), Q => 
                           B_mul_14_port);
   B_mul_reg_13_inst : DLH_X1 port map( G => n92, D => B(13), Q => 
                           B_mul_13_port);
   B_mul_reg_12_inst : DLH_X1 port map( G => n92, D => B(12), Q => 
                           B_mul_12_port);
   B_mul_reg_11_inst : DLH_X1 port map( G => n92, D => B(11), Q => 
                           B_mul_11_port);
   B_mul_reg_10_inst : DLH_X1 port map( G => n92, D => B(10), Q => 
                           B_mul_10_port);
   B_mul_reg_9_inst : DLH_X1 port map( G => n92, D => B(9), Q => B_mul_9_port);
   B_mul_reg_8_inst : DLH_X1 port map( G => n92, D => B(8), Q => B_mul_8_port);
   B_mul_reg_7_inst : DLH_X1 port map( G => n91, D => B(7), Q => B_mul_7_port);
   B_mul_reg_6_inst : DLH_X1 port map( G => n91, D => B(6), Q => B_mul_6_port);
   B_mul_reg_5_inst : DLH_X1 port map( G => n91, D => B(5), Q => B_mul_5_port);
   B_mul_reg_4_inst : DLH_X1 port map( G => n91, D => B(4), Q => B_mul_4_port);
   B_mul_reg_3_inst : DLH_X1 port map( G => n91, D => B(3), Q => B_mul_3_port);
   B_mul_reg_2_inst : DLH_X1 port map( G => n91, D => B(2), Q => B_mul_2_port);
   B_mul_reg_1_inst : DLH_X1 port map( G => n91, D => B(1), Q => B_mul_1_port);
   B_mul_reg_0_inst : DLH_X1 port map( G => n91, D => B(0), Q => B_mul_0_port);
   sel_log_reg_2_inst : DLH_X1 port map( G => n78, D => N29, Q => 
                           sel_log_2_port);
   sel_log_reg_1_inst : DLH_X1 port map( G => n78, D => N29, Q => 
                           sel_log_1_port);
   sel_log_reg_0_inst : DLH_X1 port map( G => n78, D => N28, Q => 
                           sel_log_0_port);
   A_log_reg_31_inst : DLH_X1 port map( G => n78, D => A(31), Q => 
                           A_log_31_port);
   A_log_reg_30_inst : DLH_X1 port map( G => n78, D => A(30), Q => 
                           A_log_30_port);
   A_log_reg_29_inst : DLH_X1 port map( G => n78, D => A(29), Q => 
                           A_log_29_port);
   A_log_reg_28_inst : DLH_X1 port map( G => n78, D => A(28), Q => 
                           A_log_28_port);
   A_log_reg_27_inst : DLH_X1 port map( G => n78, D => A(27), Q => 
                           A_log_27_port);
   A_log_reg_26_inst : DLH_X1 port map( G => n78, D => A(26), Q => 
                           A_log_26_port);
   A_log_reg_25_inst : DLH_X1 port map( G => n78, D => A(25), Q => 
                           A_log_25_port);
   A_log_reg_24_inst : DLH_X1 port map( G => n78, D => A(24), Q => 
                           A_log_24_port);
   A_log_reg_23_inst : DLH_X1 port map( G => n79, D => A(23), Q => 
                           A_log_23_port);
   A_log_reg_22_inst : DLH_X1 port map( G => n79, D => A(22), Q => 
                           A_log_22_port);
   A_log_reg_21_inst : DLH_X1 port map( G => n79, D => A(21), Q => 
                           A_log_21_port);
   A_log_reg_20_inst : DLH_X1 port map( G => n79, D => A(20), Q => 
                           A_log_20_port);
   A_log_reg_19_inst : DLH_X1 port map( G => n79, D => A(19), Q => 
                           A_log_19_port);
   A_log_reg_18_inst : DLH_X1 port map( G => n79, D => A(18), Q => 
                           A_log_18_port);
   A_log_reg_17_inst : DLH_X1 port map( G => n79, D => A(17), Q => 
                           A_log_17_port);
   A_log_reg_16_inst : DLH_X1 port map( G => n79, D => A(16), Q => 
                           A_log_16_port);
   A_log_reg_15_inst : DLH_X1 port map( G => n79, D => A(15), Q => 
                           A_log_15_port);
   A_log_reg_14_inst : DLH_X1 port map( G => n79, D => A(14), Q => 
                           A_log_14_port);
   A_log_reg_13_inst : DLH_X1 port map( G => n79, D => A(13), Q => 
                           A_log_13_port);
   A_log_reg_12_inst : DLH_X1 port map( G => n80, D => A(12), Q => 
                           A_log_12_port);
   A_log_reg_11_inst : DLH_X1 port map( G => n80, D => A(11), Q => 
                           A_log_11_port);
   A_log_reg_10_inst : DLH_X1 port map( G => n80, D => A(10), Q => 
                           A_log_10_port);
   A_log_reg_9_inst : DLH_X1 port map( G => n80, D => A(9), Q => A_log_9_port);
   A_log_reg_8_inst : DLH_X1 port map( G => n80, D => A(8), Q => A_log_8_port);
   A_log_reg_7_inst : DLH_X1 port map( G => n80, D => A(7), Q => A_log_7_port);
   A_log_reg_6_inst : DLH_X1 port map( G => n80, D => A(6), Q => A_log_6_port);
   A_log_reg_5_inst : DLH_X1 port map( G => n80, D => A(5), Q => A_log_5_port);
   A_log_reg_4_inst : DLH_X1 port map( G => n80, D => A(4), Q => A_log_4_port);
   A_log_reg_3_inst : DLH_X1 port map( G => n80, D => A(3), Q => A_log_3_port);
   A_log_reg_2_inst : DLH_X1 port map( G => n80, D => A(2), Q => A_log_2_port);
   A_log_reg_1_inst : DLH_X1 port map( G => n81, D => A(1), Q => A_log_1_port);
   A_log_reg_0_inst : DLH_X1 port map( G => n81, D => A(0), Q => A_log_0_port);
   B_log_reg_31_inst : DLH_X1 port map( G => n81, D => B(31), Q => 
                           B_log_31_port);
   B_log_reg_30_inst : DLH_X1 port map( G => n81, D => B(30), Q => 
                           B_log_30_port);
   B_log_reg_29_inst : DLH_X1 port map( G => n81, D => B(29), Q => 
                           B_log_29_port);
   B_log_reg_28_inst : DLH_X1 port map( G => n81, D => B(28), Q => 
                           B_log_28_port);
   B_log_reg_27_inst : DLH_X1 port map( G => n81, D => B(27), Q => 
                           B_log_27_port);
   B_log_reg_26_inst : DLH_X1 port map( G => n81, D => B(26), Q => 
                           B_log_26_port);
   B_log_reg_25_inst : DLH_X1 port map( G => n81, D => B(25), Q => 
                           B_log_25_port);
   B_log_reg_24_inst : DLH_X1 port map( G => n81, D => B(24), Q => 
                           B_log_24_port);
   B_log_reg_23_inst : DLH_X1 port map( G => n81, D => B(23), Q => 
                           B_log_23_port);
   B_log_reg_22_inst : DLH_X1 port map( G => n82, D => B(22), Q => 
                           B_log_22_port);
   B_log_reg_21_inst : DLH_X1 port map( G => n82, D => B(21), Q => 
                           B_log_21_port);
   B_log_reg_20_inst : DLH_X1 port map( G => n82, D => B(20), Q => 
                           B_log_20_port);
   B_log_reg_19_inst : DLH_X1 port map( G => n82, D => B(19), Q => 
                           B_log_19_port);
   B_log_reg_18_inst : DLH_X1 port map( G => n82, D => B(18), Q => 
                           B_log_18_port);
   B_log_reg_17_inst : DLH_X1 port map( G => n82, D => B(17), Q => 
                           B_log_17_port);
   B_log_reg_16_inst : DLH_X1 port map( G => n82, D => B(16), Q => 
                           B_log_16_port);
   B_log_reg_15_inst : DLH_X1 port map( G => n82, D => B(15), Q => 
                           B_log_15_port);
   B_log_reg_14_inst : DLH_X1 port map( G => n82, D => B(14), Q => 
                           B_log_14_port);
   B_log_reg_13_inst : DLH_X1 port map( G => n82, D => B(13), Q => 
                           B_log_13_port);
   B_log_reg_12_inst : DLH_X1 port map( G => n82, D => B(12), Q => 
                           B_log_12_port);
   B_log_reg_11_inst : DLH_X1 port map( G => n83, D => B(11), Q => 
                           B_log_11_port);
   B_log_reg_10_inst : DLH_X1 port map( G => n83, D => B(10), Q => 
                           B_log_10_port);
   B_log_reg_9_inst : DLH_X1 port map( G => n83, D => B(9), Q => B_log_9_port);
   B_log_reg_8_inst : DLH_X1 port map( G => n83, D => B(8), Q => B_log_8_port);
   B_log_reg_7_inst : DLH_X1 port map( G => n83, D => B(7), Q => B_log_7_port);
   B_log_reg_6_inst : DLH_X1 port map( G => n83, D => B(6), Q => B_log_6_port);
   B_log_reg_5_inst : DLH_X1 port map( G => n83, D => B(5), Q => B_log_5_port);
   B_log_reg_4_inst : DLH_X1 port map( G => n83, D => B(4), Q => B_log_4_port);
   B_log_reg_3_inst : DLH_X1 port map( G => n83, D => B(3), Q => B_log_3_port);
   B_log_reg_2_inst : DLH_X1 port map( G => n83, D => B(2), Q => B_log_2_port);
   B_log_reg_1_inst : DLH_X1 port map( G => n83, D => B(1), Q => B_log_1_port);
   B_log_reg_0_inst : DLH_X1 port map( G => n24, D => B(0), Q => B_log_0_port);
   sel_shift_reg_1_inst : DLH_X1 port map( G => n89, D => N32, Q => 
                           sel_shift_1_port);
   sel_shift_reg_0_inst : DLH_X1 port map( G => n89, D => N31, Q => 
                           sel_shift_0_port);
   A_sht_reg_31_inst : DLH_X1 port map( G => n89, D => A(31), Q => 
                           A_sht_31_port);
   A_sht_reg_30_inst : DLH_X1 port map( G => n89, D => A(30), Q => 
                           A_sht_30_port);
   A_sht_reg_29_inst : DLH_X1 port map( G => n89, D => A(29), Q => 
                           A_sht_29_port);
   A_sht_reg_28_inst : DLH_X1 port map( G => n89, D => A(28), Q => 
                           A_sht_28_port);
   A_sht_reg_27_inst : DLH_X1 port map( G => n89, D => A(27), Q => 
                           A_sht_27_port);
   A_sht_reg_26_inst : DLH_X1 port map( G => n89, D => A(26), Q => 
                           A_sht_26_port);
   A_sht_reg_25_inst : DLH_X1 port map( G => n89, D => A(25), Q => 
                           A_sht_25_port);
   A_sht_reg_24_inst : DLH_X1 port map( G => n89, D => A(24), Q => 
                           A_sht_24_port);
   A_sht_reg_23_inst : DLH_X1 port map( G => n89, D => A(23), Q => 
                           A_sht_23_port);
   A_sht_reg_22_inst : DLH_X1 port map( G => n88, D => A(22), Q => 
                           A_sht_22_port);
   A_sht_reg_21_inst : DLH_X1 port map( G => n88, D => A(21), Q => 
                           A_sht_21_port);
   A_sht_reg_20_inst : DLH_X1 port map( G => n88, D => A(20), Q => 
                           A_sht_20_port);
   A_sht_reg_19_inst : DLH_X1 port map( G => n88, D => A(19), Q => 
                           A_sht_19_port);
   A_sht_reg_18_inst : DLH_X1 port map( G => n88, D => A(18), Q => 
                           A_sht_18_port);
   A_sht_reg_17_inst : DLH_X1 port map( G => n88, D => A(17), Q => 
                           A_sht_17_port);
   A_sht_reg_16_inst : DLH_X1 port map( G => n88, D => A(16), Q => 
                           A_sht_16_port);
   A_sht_reg_15_inst : DLH_X1 port map( G => n88, D => A(15), Q => 
                           A_sht_15_port);
   A_sht_reg_14_inst : DLH_X1 port map( G => n88, D => A(14), Q => 
                           A_sht_14_port);
   A_sht_reg_13_inst : DLH_X1 port map( G => n88, D => A(13), Q => 
                           A_sht_13_port);
   A_sht_reg_12_inst : DLH_X1 port map( G => n88, D => A(12), Q => 
                           A_sht_12_port);
   A_sht_reg_11_inst : DLH_X1 port map( G => n87, D => A(11), Q => 
                           A_sht_11_port);
   A_sht_reg_10_inst : DLH_X1 port map( G => n87, D => A(10), Q => 
                           A_sht_10_port);
   A_sht_reg_9_inst : DLH_X1 port map( G => n87, D => A(9), Q => A_sht_9_port);
   A_sht_reg_8_inst : DLH_X1 port map( G => n87, D => A(8), Q => A_sht_8_port);
   A_sht_reg_7_inst : DLH_X1 port map( G => n87, D => A(7), Q => A_sht_7_port);
   A_sht_reg_6_inst : DLH_X1 port map( G => n87, D => A(6), Q => A_sht_6_port);
   A_sht_reg_5_inst : DLH_X1 port map( G => n87, D => A(5), Q => A_sht_5_port);
   A_sht_reg_4_inst : DLH_X1 port map( G => n87, D => A(4), Q => A_sht_4_port);
   A_sht_reg_3_inst : DLH_X1 port map( G => n87, D => A(3), Q => A_sht_3_port);
   A_sht_reg_2_inst : DLH_X1 port map( G => n87, D => A(2), Q => A_sht_2_port);
   A_sht_reg_1_inst : DLH_X1 port map( G => n87, D => A(1), Q => A_sht_1_port);
   A_sht_reg_0_inst : DLH_X1 port map( G => n86, D => A(0), Q => A_sht_0_port);
   B_sht_reg_31_inst : DLH_X1 port map( G => n86, D => B(31), Q => 
                           B_sht_31_port);
   B_sht_reg_30_inst : DLH_X1 port map( G => n86, D => B(30), Q => 
                           B_sht_30_port);
   B_sht_reg_29_inst : DLH_X1 port map( G => n86, D => B(29), Q => 
                           B_sht_29_port);
   B_sht_reg_28_inst : DLH_X1 port map( G => n86, D => B(28), Q => 
                           B_sht_28_port);
   B_sht_reg_27_inst : DLH_X1 port map( G => n86, D => B(27), Q => 
                           B_sht_27_port);
   B_sht_reg_26_inst : DLH_X1 port map( G => n86, D => B(26), Q => 
                           B_sht_26_port);
   B_sht_reg_25_inst : DLH_X1 port map( G => n86, D => B(25), Q => 
                           B_sht_25_port);
   B_sht_reg_24_inst : DLH_X1 port map( G => n86, D => B(24), Q => 
                           B_sht_24_port);
   B_sht_reg_23_inst : DLH_X1 port map( G => n86, D => B(23), Q => 
                           B_sht_23_port);
   B_sht_reg_22_inst : DLH_X1 port map( G => n86, D => B(22), Q => 
                           B_sht_22_port);
   B_sht_reg_21_inst : DLH_X1 port map( G => n85, D => B(21), Q => 
                           B_sht_21_port);
   B_sht_reg_20_inst : DLH_X1 port map( G => n85, D => B(20), Q => 
                           B_sht_20_port);
   B_sht_reg_19_inst : DLH_X1 port map( G => n85, D => B(19), Q => 
                           B_sht_19_port);
   B_sht_reg_18_inst : DLH_X1 port map( G => n85, D => B(18), Q => 
                           B_sht_18_port);
   B_sht_reg_17_inst : DLH_X1 port map( G => n85, D => B(17), Q => 
                           B_sht_17_port);
   B_sht_reg_16_inst : DLH_X1 port map( G => n85, D => B(16), Q => 
                           B_sht_16_port);
   B_sht_reg_15_inst : DLH_X1 port map( G => n85, D => B(15), Q => 
                           B_sht_15_port);
   B_sht_reg_14_inst : DLH_X1 port map( G => n85, D => B(14), Q => 
                           B_sht_14_port);
   B_sht_reg_13_inst : DLH_X1 port map( G => n85, D => B(13), Q => 
                           B_sht_13_port);
   B_sht_reg_12_inst : DLH_X1 port map( G => n85, D => B(12), Q => 
                           B_sht_12_port);
   B_sht_reg_11_inst : DLH_X1 port map( G => n85, D => B(11), Q => 
                           B_sht_11_port);
   B_sht_reg_10_inst : DLH_X1 port map( G => n84, D => B(10), Q => 
                           B_sht_10_port);
   B_sht_reg_9_inst : DLH_X1 port map( G => n84, D => B(9), Q => B_sht_9_port);
   B_sht_reg_8_inst : DLH_X1 port map( G => n84, D => B(8), Q => B_sht_8_port);
   B_sht_reg_7_inst : DLH_X1 port map( G => n84, D => B(7), Q => B_sht_7_port);
   B_sht_reg_6_inst : DLH_X1 port map( G => n84, D => B(6), Q => B_sht_6_port);
   B_sht_reg_5_inst : DLH_X1 port map( G => n84, D => B(5), Q => B_sht_5_port);
   B_sht_reg_4_inst : DLH_X1 port map( G => n84, D => B(4), Q => B_sht_4_port);
   B_sht_reg_3_inst : DLH_X1 port map( G => n84, D => B(3), Q => B_sht_3_port);
   B_sht_reg_2_inst : DLH_X1 port map( G => n84, D => B(2), Q => B_sht_2_port);
   B_sht_reg_1_inst : DLH_X1 port map( G => n84, D => B(1), Q => B_sht_1_port);
   B_sht_reg_0_inst : DLH_X1 port map( G => n84, D => B(0), Q => B_sht_0_port);
   sign_reg : DLH_X1 port map( G => N34, D => N35, Q => sign);
   sel_log_3_port <= '0';
   U63 : NAND3_X1 port map( A1 => n59, A2 => n60, A3 => n61, ZN => n58);
   U64 : XOR2_X1 port map( A => n66, B => OP(2), Z => n63);
   U65 : NAND3_X1 port map( A1 => n70, A2 => OP(2), A3 => OP(4), ZN => n69);
   U66 : NAND3_X1 port map( A1 => OP(2), A2 => n59, A3 => n70, ZN => n72);
   U67 : NAND3_X1 port map( A1 => n66, A2 => n60, A3 => n61, ZN => n57);
   U68 : NAND3_X1 port map( A1 => n65, A2 => n60, A3 => OP(3), ZN => n73);
   A_mul_reg_13_inst : DLH_X1 port map( G => n91, D => A(13), Q => 
                           A_mul_13_port);
   A_mul_reg_3_inst : DLH_X1 port map( G => n91, D => A(3), Q => A_mul_3_port);
   A_mul_reg_5_inst : DLH_X1 port map( G => n91, D => A(5), Q => A_mul_5_port);
   A_mul_reg_9_inst : DLH_X1 port map( G => n90, D => A(9), Q => A_mul_9_port);
   A_mul_reg_7_inst : DLH_X1 port map( G => n90, D => A(7), Q => A_mul_7_port);
   A_mul_reg_14_inst : DLH_X1 port map( G => n90, D => A(14), Q => 
                           A_mul_14_port);
   A_mul_reg_11_inst : DLH_X1 port map( G => n90, D => A(11), Q => 
                           A_mul_11_port);
   A_mul_reg_1_inst : DLH_X1 port map( G => n90, D => A(1), Q => A_mul_1_port);
   A_mul_reg_12_inst : DLH_X1 port map( G => n90, D => A(12), Q => 
                           A_mul_12_port);
   A_mul_reg_8_inst : DLH_X1 port map( G => n90, D => A(8), Q => A_mul_8_port);
   A_mul_reg_10_inst : DLH_X1 port map( G => n90, D => A(10), Q => 
                           A_mul_10_port);
   A_mul_reg_6_inst : DLH_X1 port map( G => n90, D => A(6), Q => A_mul_6_port);
   A_mul_reg_4_inst : DLH_X1 port map( G => n90, D => A(4), Q => A_mul_4_port);
   add_sub_reg : DLH_X1 port map( G => n93, D => N25, Q => add_sub);
   A_mul_reg_2_inst : DLH_X1 port map( G => n90, D => A(2), Q => A_mul_2_port);
   U69 : NOR4_X4 port map( A1 => OP(3), A2 => OP(4), A3 => n62, A4 => n60, ZN 
                           => N36);
   U70 : INV_X1 port map( A => n57, ZN => N28);
   U71 : OAI21_X1 port map( B1 => n73, B2 => n76, A => n67, ZN => N25);
   U72 : NAND2_X1 port map( A1 => n59, A2 => n71, ZN => n76);
   U73 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n24);
   U74 : BUF_X1 port map( A => N27, Z => n90);
   U75 : BUF_X1 port map( A => N27, Z => n91);
   U76 : BUF_X1 port map( A => N27, Z => n92);
   U77 : INV_X1 port map( A => n73, ZN => n70);
   U78 : NOR2_X1 port map( A1 => n59, A2 => n68, ZN => N32);
   U79 : INV_X1 port map( A => n67, ZN => N34);
   U80 : INV_X1 port map( A => n62, ZN => n61);
   U81 : OAI221_X1 port map( B1 => n77, B2 => n65, C1 => OP(0), C2 => OP(1), A 
                           => n62, ZN => n67);
   U82 : AOI21_X1 port map( B1 => n66, B2 => n71, A => OP(0), ZN => n77);
   U83 : NOR3_X1 port map( A1 => n59, A2 => OP(2), A3 => n73, ZN => N27);
   U84 : NOR4_X1 port map( A1 => OP(0), A2 => n63, A3 => n64, A4 => n65, ZN => 
                           N35);
   U85 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n64);
   U86 : NAND4_X1 port map( A1 => OP(1), A2 => n66, A3 => n71, A4 => n60, ZN =>
                           n68);
   U87 : INV_X1 port map( A => OP(4), ZN => n59);
   U88 : INV_X1 port map( A => OP(1), ZN => n65);
   U89 : INV_X1 port map( A => OP(3), ZN => n66);
   U90 : INV_X1 port map( A => OP(2), ZN => n71);
   U91 : INV_X1 port map( A => OP(0), ZN => n60);
   U92 : NAND2_X1 port map( A1 => OP(2), A2 => n65, ZN => n62);
   U93 : OAI21_X1 port map( B1 => n59, B2 => n57, A => n72, ZN => N29);
   U94 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N33);
   U95 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => N26);
   U96 : INV_X1 port map( A => N25, ZN => n75);
   U97 : NAND4_X1 port map( A1 => OP(4), A2 => n66, A3 => n71, A4 => n65, ZN =>
                           n74);
   U98 : NOR2_X1 port map( A1 => OP(4), A2 => n68, ZN => N31);
   U99 : CLKBUF_X1 port map( A => n24, Z => n78);
   U100 : CLKBUF_X1 port map( A => n24, Z => n79);
   U101 : CLKBUF_X1 port map( A => n24, Z => n80);
   U102 : CLKBUF_X1 port map( A => n24, Z => n81);
   U103 : CLKBUF_X1 port map( A => n24, Z => n82);
   U104 : CLKBUF_X1 port map( A => n24, Z => n83);
   U105 : CLKBUF_X1 port map( A => N33, Z => n84);
   U106 : CLKBUF_X1 port map( A => N33, Z => n85);
   U107 : CLKBUF_X1 port map( A => N33, Z => n86);
   U108 : CLKBUF_X1 port map( A => N33, Z => n87);
   U109 : CLKBUF_X1 port map( A => N33, Z => n88);
   U110 : CLKBUF_X1 port map( A => N33, Z => n89);
   U111 : CLKBUF_X1 port map( A => N26, Z => n93);
   U112 : CLKBUF_X1 port map( A => N26, Z => n94);
   U113 : CLKBUF_X1 port map( A => N26, Z => n95);
   U114 : CLKBUF_X1 port map( A => N26, Z => n96);
   U115 : CLKBUF_X1 port map( A => N26, Z => n97);
   U116 : CLKBUF_X1 port map( A => N26, Z => n98);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity CU_HW is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         flush : in std_logic_vector (1 downto 0);  JUMP_EN, RF_RD1_EN, 
         RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, MUXA_SEL, MUXB_SEL, EQ_COND : 
         out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 4);  
         SEL_STORE1, SEL_STORE0, SEL_LOAD2, SEL_LOAD1, SEL_LOAD0, DRAM_WR, 
         WB_MUX_SEL, RF_WR : out std_logic);

end CU_HW;

architecture SYN_rtl of CU_HW is

begin
   
   JUMP_EN <= '0';
   ALU_OPCODE(4) <= '0';
   ALU_OPCODE(3) <= '0';
   ALU_OPCODE(2) <= '0';
   ALU_OPCODE(1) <= '0';
   ALU_OPCODE(0) <= '0';
   RF_WR <= '0';
   WB_MUX_SEL <= '0';
   DRAM_WR <= '0';
   SEL_LOAD0 <= '0';
   SEL_LOAD1 <= '0';
   SEL_LOAD2 <= '0';
   SEL_STORE0 <= '0';
   SEL_STORE1 <= '0';
   EQ_COND <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   IMM_SEL <= '0';
   RET <= '0';
   CALL <= '0';
   RF_EN <= '0';
   RF_RD2_EN <= '0';
   RF_RD1_EN <= '0';

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity datapath is

   port( Clk, Rst : in std_logic;  Instr : in std_logic_vector (31 downto 0);  
         JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, MUXA_SEL, 
         MUXB_SEL, EQ_COND : in std_logic;  ALU_OPCODE : in std_logic_vector (0
         to 4);  SEL_STORE1, SEL_STORE0, SEL_LOAD2, SEL_LOAD1, SEL_LOAD0, 
         DRAM_WR, WB_MUX_SEL, RF_WR : in std_logic;  flush : out 
         std_logic_vector (1 downto 0);  PC_out : out std_logic_vector (31 
         downto 0));

end datapath;

architecture SYN_rtl of datapath is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff_1
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_2
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_3
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_4
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_5
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_6
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_7
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_8
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_9
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_10
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component mux_fwd_1
      port( OP, alu_out, alu_wb_in, lmd_out : in std_logic_vector (31 downto 0)
            ;  OPF : out std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (2 downto 0));
   end component;
   
   component ff_11
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_12
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_13
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component mux_fwd_0
      port( OP, alu_out, alu_wb_in, lmd_out : in std_logic_vector (31 downto 0)
            ;  OPF : out std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (2 downto 0));
   end component;
   
   component ff_14
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_15
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_16
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_17
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_18
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_19
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_20
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_21
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_22
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_23
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_24
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_25
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_26
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_27
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component counter
      port( clk, rst : in std_logic;  tc : out std_logic);
   end component;
   
   component ff_28
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component reg_N2_1
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (1 downto 0); 
            d_out : out std_logic_vector (1 downto 0));
   end component;
   
   component reg_N2_0
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (1 downto 0); 
            d_out : out std_logic_vector (1 downto 0));
   end component;
   
   component mux_pc
      port( A, B, C, D, E, F : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component ff_29
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_30
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_31
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component ff_0
      port( clk, rst, d_in : in std_logic;  d_out : out std_logic);
   end component;
   
   component reg_N32_1
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_2
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_3
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_4
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component PC_incr
      port( PC : in std_logic_vector (31 downto 0);  NPC : out std_logic_vector
            (31 downto 0));
   end component;
   
   component reg_en_N32
      port( clk, rst, en : in std_logic;  d_in : in std_logic_vector (31 downto
            0);  d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_5
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_6
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_7
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_8
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component DRAM
      port( clk, rst, WR : in std_logic;  sel_store : in std_logic_vector (1 
            downto 0);  sel_load : in std_logic_vector (2 downto 0);  addr : in
            std_logic_vector (11 downto 0);  d_in : in std_logic_vector (31 
            downto 0);  d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_9
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_10
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_11
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component sign_ext_Nstart26_Nend32
      port( Ain : in std_logic_vector (25 downto 0);  Aout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component sign_ext_Nstart16_Nend32
      port( Ain : in std_logic_vector (15 downto 0);  Aout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_12
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_13
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component stack
      port( clk, reset, enable, RD, wr : in std_logic;  datain : in 
            std_logic_vector (31 downto 0);  dataout : out std_logic_vector (31
            downto 0));
   end component;
   
   component w_reg_file_M8_N8_F4_Nbit32
      port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
            add_rd2 : in std_logic_vector (4 downto 0);  datain : in 
            std_logic_vector (31 downto 0);  out1, out2 : out std_logic_vector 
            (31 downto 0);  call, ret : in std_logic;  spill, fill : out 
            std_logic;  to_mem : out std_logic_vector (31 downto 0);  from_mem 
            : in std_logic_vector (31 downto 0));
   end component;
   
   component reg_N5_1
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0); 
            d_out : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_N5_2
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0); 
            d_out : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_N5_0
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (4 downto 0); 
            d_out : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_N6_1
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (5 downto 0); 
            d_out : out std_logic_vector (5 downto 0));
   end component;
   
   component reg_N6_0
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (5 downto 0); 
            d_out : out std_logic_vector (5 downto 0));
   end component;
   
   component reg_N32_0
      port( clk, rst : in std_logic;  d_in : in std_logic_vector (31 downto 0);
            d_out : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component cla_adder_N32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component alu
      port( A, B : in std_logic_vector (31 downto 0);  OP : in std_logic_vector
            (0 to 4);  Y1 : out std_logic_vector (31 downto 0);  cout : out 
            std_logic);
   end component;
   
   signal X_Logic0_port, flush_1_port, flush_0_port, PC_out_31, PC_out_28_port,
      PC_out_27_port, PC_out_26_port, PC_out_25_port, PC_out_24_port, 
      PC_out_23_port, PC_out_22_port, PC_out_21_port, PC_out_20_port, 
      PC_out_19_port, PC_out_18_port, PC_out_17_port, PC_out_16_port, 
      PC_out_15_port, PC_out_14_port, PC_out_13_port, PC_out_12_port, 
      PC_out_11_port, PC_out_10_port, PC_out_9_port, PC_out_8_port, 
      PC_out_7_port, PC_out_6_port, PC_out_5_port, PC_out_4_port, PC_out_3_port
      , PC_out_2_port, PC_out_1_port, PC_out_0_port, PC_enable1, 
      Instr_reg_out_31_port, Instr_reg_out_30_port, Instr_reg_out_29_port, 
      Instr_reg_out_28_port, Instr_reg_out_27_port, Instr_reg_out_26_port, 
      Instr_reg_out_25_port, Instr_reg_out_24_port, Instr_reg_out_23_port, 
      Instr_reg_out_22_port, Instr_reg_out_21_port, Instr_reg_out_20_port, 
      Instr_reg_out_19_port, Instr_reg_out_18_port, Instr_reg_out_17_port, 
      Instr_reg_out_16_port, Instr_reg_out_15_port, Instr_reg_out_14_port, 
      Instr_reg_out_13_port, Instr_reg_out_12_port, Instr_reg_out_11_port, 
      Instr_reg_out_10_port, Instr_reg_out_9_port, Instr_reg_out_8_port, 
      Instr_reg_out_7_port, Instr_reg_out_6_port, Instr_reg_out_5_port, 
      Instr_reg_out_4_port, Instr_reg_out_3_port, Instr_reg_out_2_port, 
      Instr_reg_out_1_port, Instr_reg_out_0_port, OPCODE1_5_port, 
      OPCODE1_4_port, OPCODE1_3_port, OPCODE1_2_port, OPCODE1_1_port, 
      OPCODE1_0_port, OPCODE2_5_port, OPCODE2_4_port, OPCODE2_3_port, 
      OPCODE2_2_port, OPCODE2_1_port, OPCODE2_0_port, RD_4_port, RD_3_port, 
      RD_2_port, RD_1_port, RD_0_port, RD1_4_port, RD1_3_port, RD1_2_port, 
      RD1_1_port, RD1_0_port, RD2_4_port, RD2_3_port, RD2_2_port, RD2_1_port, 
      RD2_0_port, RD3_4_port, RD3_3_port, RD3_2_port, RD3_1_port, RD3_0_port, 
      RF_write_data_31_port, RF_write_data_30_port, RF_write_data_29_port, 
      RF_write_data_28_port, RF_write_data_27_port, RF_write_data_26_port, 
      RF_write_data_25_port, RF_write_data_24_port, RF_write_data_23_port, 
      RF_write_data_22_port, RF_write_data_21_port, RF_write_data_20_port, 
      RF_write_data_19_port, RF_write_data_18_port, RF_write_data_17_port, 
      RF_write_data_16_port, RF_write_data_15_port, RF_write_data_14_port, 
      RF_write_data_13_port, RF_write_data_12_port, RF_write_data_11_port, 
      RF_write_data_10_port, RF_write_data_9_port, RF_write_data_8_port, 
      RF_write_data_7_port, RF_write_data_6_port, RF_write_data_5_port, 
      RF_write_data_4_port, RF_write_data_3_port, RF_write_data_2_port, 
      RF_write_data_1_port, RF_write_data_0_port, RF_out_A_31_port, 
      RF_out_A_30_port, RF_out_A_29_port, RF_out_A_28_port, RF_out_A_27_port, 
      RF_out_A_26_port, RF_out_A_25_port, RF_out_A_24_port, RF_out_A_23_port, 
      RF_out_A_22_port, RF_out_A_21_port, RF_out_A_20_port, RF_out_A_19_port, 
      RF_out_A_18_port, RF_out_A_17_port, RF_out_A_16_port, RF_out_A_15_port, 
      RF_out_A_14_port, RF_out_A_13_port, RF_out_A_12_port, RF_out_A_11_port, 
      RF_out_A_10_port, RF_out_A_9_port, RF_out_A_8_port, RF_out_A_7_port, 
      RF_out_A_6_port, RF_out_A_5_port, RF_out_A_4_port, RF_out_A_3_port, 
      RF_out_A_2_port, RF_out_A_1_port, RF_out_A_0_port, RF_out_B_31_port, 
      RF_out_B_30_port, RF_out_B_29_port, RF_out_B_28_port, RF_out_B_27_port, 
      RF_out_B_26_port, RF_out_B_25_port, RF_out_B_24_port, RF_out_B_23_port, 
      RF_out_B_22_port, RF_out_B_21_port, RF_out_B_20_port, RF_out_B_19_port, 
      RF_out_B_18_port, RF_out_B_17_port, RF_out_B_16_port, RF_out_B_15_port, 
      RF_out_B_14_port, RF_out_B_13_port, RF_out_B_12_port, RF_out_B_11_port, 
      RF_out_B_10_port, RF_out_B_9_port, RF_out_B_8_port, RF_out_B_7_port, 
      RF_out_B_6_port, RF_out_B_5_port, RF_out_B_4_port, RF_out_B_3_port, 
      RF_out_B_2_port, RF_out_B_1_port, RF_out_B_0_port, SPILL, FILL, 
      spill_to_stack_31_port, spill_to_stack_30_port, spill_to_stack_29_port, 
      spill_to_stack_28_port, spill_to_stack_27_port, spill_to_stack_26_port, 
      spill_to_stack_25_port, spill_to_stack_24_port, spill_to_stack_23_port, 
      spill_to_stack_22_port, spill_to_stack_21_port, spill_to_stack_20_port, 
      spill_to_stack_19_port, spill_to_stack_18_port, spill_to_stack_17_port, 
      spill_to_stack_16_port, spill_to_stack_15_port, spill_to_stack_14_port, 
      spill_to_stack_13_port, spill_to_stack_12_port, spill_to_stack_11_port, 
      spill_to_stack_10_port, spill_to_stack_9_port, spill_to_stack_8_port, 
      spill_to_stack_7_port, spill_to_stack_6_port, spill_to_stack_5_port, 
      spill_to_stack_4_port, spill_to_stack_3_port, spill_to_stack_2_port, 
      spill_to_stack_1_port, spill_to_stack_0_port, fill_from_stack_31_port, 
      fill_from_stack_30_port, fill_from_stack_29_port, fill_from_stack_28_port
      , fill_from_stack_27_port, fill_from_stack_26_port, 
      fill_from_stack_25_port, fill_from_stack_24_port, fill_from_stack_23_port
      , fill_from_stack_22_port, fill_from_stack_21_port, 
      fill_from_stack_20_port, fill_from_stack_19_port, fill_from_stack_18_port
      , fill_from_stack_17_port, fill_from_stack_16_port, 
      fill_from_stack_15_port, fill_from_stack_14_port, fill_from_stack_13_port
      , fill_from_stack_12_port, fill_from_stack_11_port, 
      fill_from_stack_10_port, fill_from_stack_9_port, fill_from_stack_8_port, 
      fill_from_stack_7_port, fill_from_stack_6_port, fill_from_stack_5_port, 
      fill_from_stack_4_port, fill_from_stack_3_port, fill_from_stack_2_port, 
      fill_from_stack_1_port, fill_from_stack_0_port, A_reg_out_31_port, 
      A_reg_out_30_port, A_reg_out_29_port, A_reg_out_28_port, 
      A_reg_out_27_port, A_reg_out_26_port, A_reg_out_25_port, 
      A_reg_out_24_port, A_reg_out_23_port, A_reg_out_22_port, 
      A_reg_out_21_port, A_reg_out_20_port, A_reg_out_19_port, 
      A_reg_out_18_port, A_reg_out_17_port, A_reg_out_16_port, 
      A_reg_out_15_port, A_reg_out_14_port, A_reg_out_13_port, 
      A_reg_out_12_port, A_reg_out_11_port, A_reg_out_10_port, A_reg_out_9_port
      , A_reg_out_8_port, A_reg_out_7_port, A_reg_out_6_port, A_reg_out_5_port,
      A_reg_out_4_port, A_reg_out_3_port, A_reg_out_2_port, A_reg_out_1_port, 
      A_reg_out_0_port, B_reg_out_31_port, B_reg_out_30_port, B_reg_out_29_port
      , B_reg_out_28_port, B_reg_out_27_port, B_reg_out_26_port, 
      B_reg_out_25_port, B_reg_out_24_port, B_reg_out_23_port, 
      B_reg_out_22_port, B_reg_out_21_port, B_reg_out_20_port, 
      B_reg_out_19_port, B_reg_out_18_port, B_reg_out_17_port, 
      B_reg_out_16_port, B_reg_out_15_port, B_reg_out_14_port, 
      B_reg_out_13_port, B_reg_out_12_port, B_reg_out_11_port, 
      B_reg_out_10_port, B_reg_out_9_port, B_reg_out_8_port, B_reg_out_7_port, 
      B_reg_out_6_port, B_reg_out_5_port, B_reg_out_4_port, B_reg_out_3_port, 
      B_reg_out_2_port, B_reg_out_1_port, B_reg_out_0_port, 
      Immediate_16_extended_31_port, Immediate_16_extended_30_port, 
      Immediate_16_extended_29_port, Immediate_16_extended_28_port, 
      Immediate_16_extended_27_port, Immediate_16_extended_26_port, 
      Immediate_16_extended_25_port, Immediate_16_extended_24_port, 
      Immediate_16_extended_23_port, Immediate_16_extended_22_port, 
      Immediate_16_extended_21_port, Immediate_16_extended_20_port, 
      Immediate_16_extended_19_port, Immediate_16_extended_18_port, 
      Immediate_16_extended_17_port, Immediate_16_extended_16_port, 
      Immediate_16_extended_15_port, Immediate_16_extended_14_port, 
      Immediate_16_extended_13_port, Immediate_16_extended_12_port, 
      Immediate_16_extended_11_port, Immediate_16_extended_10_port, 
      Immediate_16_extended_9_port, Immediate_16_extended_8_port, 
      Immediate_16_extended_7_port, Immediate_16_extended_6_port, 
      Immediate_16_extended_5_port, Immediate_16_extended_4_port, 
      Immediate_16_extended_3_port, Immediate_16_extended_2_port, 
      Immediate_16_extended_1_port, Immediate_16_extended_0_port, 
      Immediate_26_extended_31_port, Immediate_26_extended_30_port, 
      Immediate_26_extended_29_port, Immediate_26_extended_28_port, 
      Immediate_26_extended_27_port, Immediate_26_extended_26_port, 
      Immediate_26_extended_25_port, Immediate_26_extended_24_port, 
      Immediate_26_extended_23_port, Immediate_26_extended_22_port, 
      Immediate_26_extended_21_port, Immediate_26_extended_20_port, 
      Immediate_26_extended_19_port, Immediate_26_extended_18_port, 
      Immediate_26_extended_17_port, Immediate_26_extended_16_port, 
      Immediate_26_extended_15_port, Immediate_26_extended_14_port, 
      Immediate_26_extended_13_port, Immediate_26_extended_12_port, 
      Immediate_26_extended_11_port, Immediate_26_extended_10_port, 
      Immediate_26_extended_9_port, Immediate_26_extended_8_port, 
      Immediate_26_extended_7_port, Immediate_26_extended_6_port, 
      Immediate_26_extended_5_port, Immediate_26_extended_4_port, 
      Immediate_26_extended_3_port, Immediate_26_extended_2_port, 
      Immediate_26_extended_1_port, Immediate_26_extended_0_port, 
      Immediate_selected_31_port, Immediate_selected_30_port, 
      Immediate_selected_29_port, Immediate_selected_28_port, 
      Immediate_selected_27_port, Immediate_selected_26_port, 
      Immediate_selected_25_port, Immediate_selected_24_port, 
      Immediate_selected_23_port, Immediate_selected_22_port, 
      Immediate_selected_21_port, Immediate_selected_20_port, 
      Immediate_selected_19_port, Immediate_selected_18_port, 
      Immediate_selected_17_port, Immediate_selected_16_port, 
      Immediate_selected_15_port, Immediate_selected_14_port, 
      Immediate_selected_13_port, Immediate_selected_12_port, 
      Immediate_selected_11_port, Immediate_selected_10_port, 
      Immediate_selected_9_port, Immediate_selected_8_port, 
      Immediate_selected_7_port, Immediate_selected_6_port, 
      Immediate_selected_5_port, Immediate_selected_4_port, 
      Immediate_selected_3_port, Immediate_selected_2_port, 
      Immediate_selected_1_port, Immediate_selected_0_port, 
      Immediate_clocked_31_port, Immediate_clocked_30_port, 
      Immediate_clocked_29_port, Immediate_clocked_28_port, 
      Immediate_clocked_27_port, Immediate_clocked_26_port, 
      Immediate_clocked_25_port, Immediate_clocked_24_port, 
      Immediate_clocked_23_port, Immediate_clocked_22_port, 
      Immediate_clocked_21_port, Immediate_clocked_20_port, 
      Immediate_clocked_19_port, Immediate_clocked_18_port, 
      Immediate_clocked_17_port, Immediate_clocked_16_port, 
      Immediate_clocked_15_port, Immediate_clocked_14_port, 
      Immediate_clocked_13_port, Immediate_clocked_12_port, 
      Immediate_clocked_11_port, Immediate_clocked_10_port, 
      Immediate_clocked_9_port, Immediate_clocked_8_port, 
      Immediate_clocked_7_port, Immediate_clocked_6_port, 
      Immediate_clocked_5_port, Immediate_clocked_4_port, 
      Immediate_clocked_3_port, Immediate_clocked_2_port, 
      Immediate_clocked_1_port, Immediate_clocked_0_port, NPC2_31_port, 
      NPC2_30_port, NPC2_29_port, NPC2_28_port, NPC2_27_port, NPC2_26_port, 
      NPC2_25_port, NPC2_24_port, NPC2_23_port, NPC2_22_port, NPC2_21_port, 
      NPC2_20_port, NPC2_19_port, NPC2_18_port, NPC2_17_port, NPC2_16_port, 
      NPC2_15_port, NPC2_14_port, NPC2_13_port, NPC2_12_port, NPC2_11_port, 
      NPC2_10_port, NPC2_9_port, NPC2_8_port, NPC2_7_port, NPC2_6_port, 
      NPC2_5_port, NPC2_4_port, NPC2_3_port, NPC2_2_port, NPC2_1_port, 
      NPC2_0_port, ALU_operand_1_31_port, ALU_operand_1_30_port, 
      ALU_operand_1_29_port, ALU_operand_1_28_port, ALU_operand_1_27_port, 
      ALU_operand_1_26_port, ALU_operand_1_25_port, ALU_operand_1_24_port, 
      ALU_operand_1_23_port, ALU_operand_1_22_port, ALU_operand_1_21_port, 
      ALU_operand_1_20_port, ALU_operand_1_19_port, ALU_operand_1_18_port, 
      ALU_operand_1_17_port, ALU_operand_1_16_port, ALU_operand_1_15_port, 
      ALU_operand_1_14_port, ALU_operand_1_13_port, ALU_operand_1_12_port, 
      ALU_operand_1_11_port, ALU_operand_1_10_port, ALU_operand_1_9_port, 
      ALU_operand_1_8_port, ALU_operand_1_7_port, ALU_operand_1_6_port, 
      ALU_operand_1_5_port, ALU_operand_1_4_port, ALU_operand_1_3_port, 
      ALU_operand_1_2_port, ALU_operand_1_1_port, ALU_operand_1_0_port, 
      ALU_operand_2_31_port, ALU_operand_2_30_port, ALU_operand_2_29_port, 
      ALU_operand_2_28_port, ALU_operand_2_27_port, ALU_operand_2_26_port, 
      ALU_operand_2_25_port, ALU_operand_2_24_port, ALU_operand_2_23_port, 
      ALU_operand_2_22_port, ALU_operand_2_21_port, ALU_operand_2_20_port, 
      ALU_operand_2_19_port, ALU_operand_2_18_port, ALU_operand_2_17_port, 
      ALU_operand_2_16_port, ALU_operand_2_15_port, ALU_operand_2_14_port, 
      ALU_operand_2_13_port, ALU_operand_2_12_port, ALU_operand_2_11_port, 
      ALU_operand_2_10_port, ALU_operand_2_9_port, ALU_operand_2_8_port, 
      ALU_operand_2_7_port, ALU_operand_2_6_port, ALU_operand_2_5_port, 
      ALU_operand_2_4_port, ALU_operand_2_3_port, ALU_operand_2_2_port, 
      ALU_operand_2_1_port, ALU_operand_2_0_port, ALU_OPCODE_in_4_port, 
      ALU_OPCODE_in_3_port, ALU_OPCODE_in_2_port, ALU_OPCODE_in_1_port, 
      ALU_OPCODE_in_0_port, ALU_operand_1_FWD_31_port, 
      ALU_operand_1_FWD_30_port, ALU_operand_1_FWD_29_port, 
      ALU_operand_1_FWD_28_port, ALU_operand_1_FWD_27_port, 
      ALU_operand_1_FWD_26_port, ALU_operand_1_FWD_25_port, 
      ALU_operand_1_FWD_24_port, ALU_operand_1_FWD_23_port, 
      ALU_operand_1_FWD_22_port, ALU_operand_1_FWD_21_port, 
      ALU_operand_1_FWD_20_port, ALU_operand_1_FWD_19_port, 
      ALU_operand_1_FWD_18_port, ALU_operand_1_FWD_17_port, 
      ALU_operand_1_FWD_16_port, ALU_operand_1_FWD_15_port, 
      ALU_operand_1_FWD_14_port, ALU_operand_1_FWD_13_port, 
      ALU_operand_1_FWD_12_port, ALU_operand_1_FWD_11_port, 
      ALU_operand_1_FWD_10_port, ALU_operand_1_FWD_9_port, 
      ALU_operand_1_FWD_8_port, ALU_operand_1_FWD_7_port, 
      ALU_operand_1_FWD_6_port, ALU_operand_1_FWD_5_port, 
      ALU_operand_1_FWD_4_port, ALU_operand_1_FWD_3_port, 
      ALU_operand_1_FWD_2_port, ALU_operand_1_FWD_1_port, 
      ALU_operand_1_FWD_0_port, ALU_operand_2_FWD_31_port, 
      ALU_operand_2_FWD_30_port, ALU_operand_2_FWD_29_port, 
      ALU_operand_2_FWD_28_port, ALU_operand_2_FWD_27_port, 
      ALU_operand_2_FWD_26_port, ALU_operand_2_FWD_25_port, 
      ALU_operand_2_FWD_24_port, ALU_operand_2_FWD_23_port, 
      ALU_operand_2_FWD_22_port, ALU_operand_2_FWD_21_port, 
      ALU_operand_2_FWD_20_port, ALU_operand_2_FWD_19_port, 
      ALU_operand_2_FWD_18_port, ALU_operand_2_FWD_17_port, 
      ALU_operand_2_FWD_16_port, ALU_operand_2_FWD_15_port, 
      ALU_operand_2_FWD_14_port, ALU_operand_2_FWD_13_port, 
      ALU_operand_2_FWD_12_port, ALU_operand_2_FWD_11_port, 
      ALU_operand_2_FWD_10_port, ALU_operand_2_FWD_9_port, 
      ALU_operand_2_FWD_8_port, ALU_operand_2_FWD_7_port, 
      ALU_operand_2_FWD_6_port, ALU_operand_2_FWD_5_port, 
      ALU_operand_2_FWD_4_port, ALU_operand_2_FWD_3_port, 
      ALU_operand_2_FWD_2_port, ALU_operand_2_FWD_1_port, 
      ALU_operand_2_FWD_0_port, ALU_output_31_port, ALU_output_30_port, 
      ALU_output_29_port, ALU_output_28_port, ALU_output_27_port, 
      ALU_output_26_port, ALU_output_25_port, ALU_output_24_port, 
      ALU_output_23_port, ALU_output_22_port, ALU_output_21_port, 
      ALU_output_20_port, ALU_output_19_port, ALU_output_18_port, 
      ALU_output_17_port, ALU_output_16_port, ALU_output_15_port, 
      ALU_output_14_port, ALU_output_13_port, ALU_output_12_port, 
      ALU_output_11_port, ALU_output_10_port, ALU_output_9_port, 
      ALU_output_8_port, ALU_output_7_port, ALU_output_6_port, 
      ALU_output_5_port, ALU_output_4_port, ALU_output_3_port, 
      ALU_output_2_port, ALU_output_1_port, ALU_output_0_port, JAL_op2, 
      ALU_output_FWD_31_port, ALU_output_FWD_30_port, ALU_output_FWD_29_port, 
      ALU_output_FWD_28_port, ALU_output_FWD_27_port, ALU_output_FWD_26_port, 
      ALU_output_FWD_25_port, ALU_output_FWD_24_port, ALU_output_FWD_23_port, 
      ALU_output_FWD_22_port, ALU_output_FWD_21_port, ALU_output_FWD_20_port, 
      ALU_output_FWD_19_port, ALU_output_FWD_18_port, ALU_output_FWD_17_port, 
      ALU_output_FWD_16_port, ALU_output_FWD_15_port, ALU_output_FWD_14_port, 
      ALU_output_FWD_13_port, ALU_output_FWD_12_port, ALU_output_FWD_11_port, 
      ALU_output_FWD_10_port, ALU_output_FWD_9_port, ALU_output_FWD_8_port, 
      ALU_output_FWD_7_port, ALU_output_FWD_6_port, ALU_output_FWD_5_port, 
      ALU_output_FWD_4_port, ALU_output_FWD_3_port, ALU_output_FWD_2_port, 
      ALU_output_FWD_1_port, ALU_output_FWD_0_port, ALU_reg_out_31_port, 
      ALU_reg_out_30_port, ALU_reg_out_29_port, ALU_reg_out_28_port, 
      ALU_reg_out_27_port, ALU_reg_out_26_port, ALU_reg_out_25_port, 
      ALU_reg_out_24_port, ALU_reg_out_23_port, ALU_reg_out_22_port, 
      ALU_reg_out_21_port, ALU_reg_out_20_port, ALU_reg_out_19_port, 
      ALU_reg_out_18_port, ALU_reg_out_17_port, ALU_reg_out_16_port, 
      ALU_reg_out_15_port, ALU_reg_out_14_port, ALU_reg_out_13_port, 
      ALU_reg_out_12_port, ALU_reg_out_11_port, ALU_reg_out_10_port, 
      ALU_reg_out_9_port, ALU_reg_out_8_port, ALU_reg_out_7_port, 
      ALU_reg_out_6_port, ALU_reg_out_5_port, ALU_reg_out_4_port, 
      ALU_reg_out_3_port, ALU_reg_out_2_port, ALU_reg_out_1_port, 
      ALU_reg_out_0_port, DRAM_write_data_31_port, DRAM_write_data_30_port, 
      DRAM_write_data_29_port, DRAM_write_data_28_port, DRAM_write_data_27_port
      , DRAM_write_data_26_port, DRAM_write_data_25_port, 
      DRAM_write_data_24_port, DRAM_write_data_23_port, DRAM_write_data_22_port
      , DRAM_write_data_21_port, DRAM_write_data_20_port, 
      DRAM_write_data_19_port, DRAM_write_data_18_port, DRAM_write_data_17_port
      , DRAM_write_data_16_port, DRAM_write_data_15_port, 
      DRAM_write_data_14_port, DRAM_write_data_13_port, DRAM_write_data_12_port
      , DRAM_write_data_11_port, DRAM_write_data_10_port, 
      DRAM_write_data_9_port, DRAM_write_data_8_port, DRAM_write_data_7_port, 
      DRAM_write_data_6_port, DRAM_write_data_5_port, DRAM_write_data_4_port, 
      DRAM_write_data_3_port, DRAM_write_data_2_port, DRAM_write_data_1_port, 
      DRAM_write_data_0_port, DRAM_write_data_FWD_31_port, 
      DRAM_write_data_FWD_30_port, DRAM_write_data_FWD_29_port, 
      DRAM_write_data_FWD_28_port, DRAM_write_data_FWD_27_port, 
      DRAM_write_data_FWD_26_port, DRAM_write_data_FWD_25_port, 
      DRAM_write_data_FWD_24_port, DRAM_write_data_FWD_23_port, 
      DRAM_write_data_FWD_22_port, DRAM_write_data_FWD_21_port, 
      DRAM_write_data_FWD_20_port, DRAM_write_data_FWD_19_port, 
      DRAM_write_data_FWD_18_port, DRAM_write_data_FWD_17_port, 
      DRAM_write_data_FWD_16_port, DRAM_write_data_FWD_15_port, 
      DRAM_write_data_FWD_14_port, DRAM_write_data_FWD_13_port, 
      DRAM_write_data_FWD_12_port, DRAM_write_data_FWD_11_port, 
      DRAM_write_data_FWD_10_port, DRAM_write_data_FWD_9_port, 
      DRAM_write_data_FWD_8_port, DRAM_write_data_FWD_7_port, 
      DRAM_write_data_FWD_6_port, DRAM_write_data_FWD_5_port, 
      DRAM_write_data_FWD_4_port, DRAM_write_data_FWD_3_port, 
      DRAM_write_data_FWD_2_port, DRAM_write_data_FWD_1_port, 
      DRAM_write_data_FWD_0_port, DRAM_read_data_31_port, 
      DRAM_read_data_30_port, DRAM_read_data_29_port, DRAM_read_data_28_port, 
      DRAM_read_data_27_port, DRAM_read_data_26_port, DRAM_read_data_25_port, 
      DRAM_read_data_24_port, DRAM_read_data_23_port, DRAM_read_data_22_port, 
      DRAM_read_data_21_port, DRAM_read_data_20_port, DRAM_read_data_19_port, 
      DRAM_read_data_18_port, DRAM_read_data_17_port, DRAM_read_data_16_port, 
      DRAM_read_data_15_port, DRAM_read_data_14_port, DRAM_read_data_13_port, 
      DRAM_read_data_12_port, DRAM_read_data_11_port, DRAM_read_data_10_port, 
      DRAM_read_data_9_port, DRAM_read_data_8_port, DRAM_read_data_7_port, 
      DRAM_read_data_6_port, DRAM_read_data_5_port, DRAM_read_data_4_port, 
      DRAM_read_data_3_port, DRAM_read_data_2_port, DRAM_read_data_1_port, 
      DRAM_read_data_0_port, LMD_reg_out_31_port, LMD_reg_out_30_port, 
      LMD_reg_out_29_port, LMD_reg_out_28_port, LMD_reg_out_27_port, 
      LMD_reg_out_26_port, LMD_reg_out_25_port, LMD_reg_out_24_port, 
      LMD_reg_out_23_port, LMD_reg_out_22_port, LMD_reg_out_21_port, 
      LMD_reg_out_20_port, LMD_reg_out_19_port, LMD_reg_out_18_port, 
      LMD_reg_out_17_port, LMD_reg_out_16_port, LMD_reg_out_15_port, 
      LMD_reg_out_14_port, LMD_reg_out_13_port, LMD_reg_out_12_port, 
      LMD_reg_out_11_port, LMD_reg_out_10_port, LMD_reg_out_9_port, 
      LMD_reg_out_8_port, LMD_reg_out_7_port, LMD_reg_out_6_port, 
      LMD_reg_out_5_port, LMD_reg_out_4_port, LMD_reg_out_3_port, 
      LMD_reg_out_2_port, LMD_reg_out_1_port, LMD_reg_out_0_port, 
      LMD_reg_out1_31_port, LMD_reg_out1_30_port, LMD_reg_out1_29_port, 
      LMD_reg_out1_28_port, LMD_reg_out1_27_port, LMD_reg_out1_26_port, 
      LMD_reg_out1_25_port, LMD_reg_out1_24_port, LMD_reg_out1_23_port, 
      LMD_reg_out1_22_port, LMD_reg_out1_21_port, LMD_reg_out1_20_port, 
      LMD_reg_out1_19_port, LMD_reg_out1_18_port, LMD_reg_out1_17_port, 
      LMD_reg_out1_16_port, LMD_reg_out1_15_port, LMD_reg_out1_14_port, 
      LMD_reg_out1_13_port, LMD_reg_out1_12_port, LMD_reg_out1_11_port, 
      LMD_reg_out1_10_port, LMD_reg_out1_9_port, LMD_reg_out1_8_port, 
      LMD_reg_out1_7_port, LMD_reg_out1_6_port, LMD_reg_out1_5_port, 
      LMD_reg_out1_4_port, LMD_reg_out1_3_port, LMD_reg_out1_2_port, 
      LMD_reg_out1_1_port, LMD_reg_out1_0_port, ALU_WB_out_31_port, 
      ALU_WB_out_30_port, ALU_WB_out_29_port, ALU_WB_out_28_port, 
      ALU_WB_out_27_port, ALU_WB_out_26_port, ALU_WB_out_25_port, 
      ALU_WB_out_24_port, ALU_WB_out_23_port, ALU_WB_out_22_port, 
      ALU_WB_out_21_port, ALU_WB_out_20_port, ALU_WB_out_19_port, 
      ALU_WB_out_18_port, ALU_WB_out_17_port, ALU_WB_out_16_port, 
      ALU_WB_out_15_port, ALU_WB_out_14_port, ALU_WB_out_13_port, 
      ALU_WB_out_12_port, ALU_WB_out_11_port, ALU_WB_out_10_port, 
      ALU_WB_out_9_port, ALU_WB_out_8_port, ALU_WB_out_7_port, 
      ALU_WB_out_6_port, ALU_WB_out_5_port, ALU_WB_out_4_port, 
      ALU_WB_out_3_port, ALU_WB_out_2_port, ALU_WB_out_1_port, 
      ALU_WB_out_0_port, ALU_WB_out1_31_port, ALU_WB_out1_30_port, 
      ALU_WB_out1_29_port, ALU_WB_out1_28_port, ALU_WB_out1_27_port, 
      ALU_WB_out1_26_port, ALU_WB_out1_25_port, ALU_WB_out1_24_port, 
      ALU_WB_out1_23_port, ALU_WB_out1_22_port, ALU_WB_out1_21_port, 
      ALU_WB_out1_20_port, ALU_WB_out1_19_port, ALU_WB_out1_18_port, 
      ALU_WB_out1_17_port, ALU_WB_out1_16_port, ALU_WB_out1_15_port, 
      ALU_WB_out1_14_port, ALU_WB_out1_13_port, ALU_WB_out1_12_port, 
      ALU_WB_out1_11_port, ALU_WB_out1_10_port, ALU_WB_out1_9_port, 
      ALU_WB_out1_8_port, ALU_WB_out1_7_port, ALU_WB_out1_6_port, 
      ALU_WB_out1_5_port, ALU_WB_out1_4_port, ALU_WB_out1_3_port, 
      ALU_WB_out1_2_port, ALU_WB_out1_1_port, ALU_WB_out1_0_port, 
      WB_mux_out_31_port, WB_mux_out_30_port, WB_mux_out_29_port, 
      WB_mux_out_28_port, WB_mux_out_27_port, WB_mux_out_26_port, 
      WB_mux_out_25_port, WB_mux_out_24_port, WB_mux_out_23_port, 
      WB_mux_out_22_port, WB_mux_out_21_port, WB_mux_out_20_port, 
      WB_mux_out_19_port, WB_mux_out_18_port, WB_mux_out_17_port, 
      WB_mux_out_16_port, WB_mux_out_15_port, WB_mux_out_14_port, 
      WB_mux_out_13_port, WB_mux_out_12_port, WB_mux_out_11_port, 
      WB_mux_out_10_port, WB_mux_out_9_port, WB_mux_out_8_port, 
      WB_mux_out_7_port, WB_mux_out_6_port, WB_mux_out_5_port, 
      WB_mux_out_4_port, WB_mux_out_3_port, WB_mux_out_2_port, 
      WB_mux_out_1_port, WB_mux_out_0_port, NPC4_31_port, NPC4_30_port, 
      NPC4_29_port, NPC4_28_port, NPC4_27_port, NPC4_26_port, NPC4_25_port, 
      NPC4_24_port, NPC4_23_port, NPC4_22_port, NPC4_21_port, NPC4_20_port, 
      NPC4_19_port, NPC4_18_port, NPC4_17_port, NPC4_16_port, NPC4_15_port, 
      NPC4_14_port, NPC4_13_port, NPC4_12_port, NPC4_11_port, NPC4_10_port, 
      NPC4_9_port, NPC4_8_port, NPC4_7_port, NPC4_6_port, NPC4_5_port, 
      NPC4_4_port, NPC4_3_port, NPC4_2_port, NPC4_1_port, NPC4_0_port, JAL_op4,
      PC_enable_fixed, PC_reg_in_31_port, PC_reg_in_30_port, PC_reg_in_29_port,
      PC_reg_in_28_port, PC_reg_in_27_port, PC_reg_in_26_port, 
      PC_reg_in_25_port, PC_reg_in_24_port, PC_reg_in_23_port, 
      PC_reg_in_22_port, PC_reg_in_21_port, PC_reg_in_20_port, 
      PC_reg_in_19_port, PC_reg_in_18_port, PC_reg_in_17_port, 
      PC_reg_in_16_port, PC_reg_in_15_port, PC_reg_in_14_port, 
      PC_reg_in_13_port, PC_reg_in_12_port, PC_reg_in_11_port, 
      PC_reg_in_10_port, PC_reg_in_9_port, PC_reg_in_8_port, PC_reg_in_7_port, 
      PC_reg_in_6_port, PC_reg_in_5_port, PC_reg_in_4_port, PC_reg_in_3_port, 
      PC_reg_in_2_port, PC_reg_in_1_port, PC_reg_in_0_port, PC_reg_out_1_port, 
      PC_reg_out_0_port, NPC_31_port, NPC_30_port, NPC_29_port, NPC_28_port, 
      NPC_27_port, NPC_26_port, NPC_25_port, NPC_24_port, NPC_23_port, 
      NPC_22_port, NPC_21_port, NPC_20_port, NPC_19_port, NPC_18_port, 
      NPC_17_port, NPC_16_port, NPC_15_port, NPC_14_port, NPC_13_port, 
      NPC_12_port, NPC_11_port, NPC_10_port, NPC_9_port, NPC_8_port, NPC_7_port
      , NPC_6_port, NPC_5_port, NPC_4_port, NPC_3_port, NPC_2_port, NPC_1_port,
      NPC_0_port, NPC1_31_port, NPC1_30_port, NPC1_29_port, NPC1_28_port, 
      NPC1_27_port, NPC1_26_port, NPC1_25_port, NPC1_24_port, NPC1_23_port, 
      NPC1_22_port, NPC1_21_port, NPC1_20_port, NPC1_19_port, NPC1_18_port, 
      NPC1_17_port, NPC1_16_port, NPC1_15_port, NPC1_14_port, NPC1_13_port, 
      NPC1_12_port, NPC1_11_port, NPC1_10_port, NPC1_9_port, NPC1_8_port, 
      NPC1_7_port, NPC1_6_port, NPC1_5_port, NPC1_4_port, NPC1_3_port, 
      NPC1_2_port, NPC1_1_port, NPC1_0_port, NPC3_31_port, NPC3_30_port, 
      NPC3_29_port, NPC3_28_port, NPC3_27_port, NPC3_26_port, NPC3_25_port, 
      NPC3_24_port, NPC3_23_port, NPC3_22_port, NPC3_21_port, NPC3_20_port, 
      NPC3_19_port, NPC3_18_port, NPC3_17_port, NPC3_16_port, NPC3_15_port, 
      NPC3_14_port, NPC3_13_port, NPC3_12_port, NPC3_11_port, NPC3_10_port, 
      NPC3_9_port, NPC3_8_port, NPC3_7_port, NPC3_6_port, NPC3_5_port, 
      NPC3_4_port, NPC3_3_port, NPC3_2_port, NPC3_1_port, NPC3_0_port, JUMP_EN1
      , JUMP_EN2, BRANCH_op2, forward_branch, forward_branch1, forward_branch2,
      JR_op, BRANCH_op, PC_mux_sel_2_port, PC_mux_sel_0_port, JR_op1, PC_enable
      , PC_displaced_31_port, PC_displaced_30_port, PC_displaced_29_port, 
      PC_displaced_28_port, PC_displaced_27_port, PC_displaced_26_port, 
      PC_displaced_25_port, PC_displaced_24_port, PC_displaced_23_port, 
      PC_displaced_22_port, PC_displaced_21_port, PC_displaced_20_port, 
      PC_displaced_19_port, PC_displaced_18_port, PC_displaced_17_port, 
      PC_displaced_16_port, PC_displaced_15_port, PC_displaced_14_port, 
      PC_displaced_13_port, PC_displaced_12_port, PC_displaced_11_port, 
      PC_displaced_10_port, PC_displaced_9_port, PC_displaced_8_port, 
      PC_displaced_7_port, PC_displaced_6_port, PC_displaced_5_port, 
      PC_displaced_4_port, PC_displaced_3_port, PC_displaced_2_port, 
      PC_displaced_1_port, PC_displaced_0_port, RF_out_A_FWD_31_port, 
      RF_out_A_FWD_30_port, RF_out_A_FWD_29_port, RF_out_A_FWD_28_port, 
      RF_out_A_FWD_27_port, RF_out_A_FWD_26_port, RF_out_A_FWD_25_port, 
      RF_out_A_FWD_24_port, RF_out_A_FWD_23_port, RF_out_A_FWD_22_port, 
      RF_out_A_FWD_21_port, RF_out_A_FWD_20_port, RF_out_A_FWD_19_port, 
      RF_out_A_FWD_18_port, RF_out_A_FWD_17_port, RF_out_A_FWD_16_port, 
      RF_out_A_FWD_15_port, RF_out_A_FWD_14_port, RF_out_A_FWD_13_port, 
      RF_out_A_FWD_12_port, RF_out_A_FWD_11_port, RF_out_A_FWD_10_port, 
      RF_out_A_FWD_9_port, RF_out_A_FWD_8_port, RF_out_A_FWD_7_port, 
      RF_out_A_FWD_6_port, RF_out_A_FWD_5_port, RF_out_A_FWD_4_port, 
      RF_out_A_FWD_3_port, RF_out_A_FWD_2_port, RF_out_A_FWD_1_port, 
      RF_out_A_FWD_0_port, PC_Immediate_displacement_31_port, 
      PC_Immediate_displacement_24_port, PC_Immediate_displacement_23_port, 
      PC_Immediate_displacement_22_port, PC_Immediate_displacement_21_port, 
      PC_Immediate_displacement_20_port, PC_Immediate_displacement_19_port, 
      PC_Immediate_displacement_18_port, PC_Immediate_displacement_17_port, 
      PC_Immediate_displacement_16_port, LOAD_op1, STORE_op, flush0_1_port, 
      flush0_0_port, flush2_1_port, flush2_0_port, bootstrap, JAL_op, JAL_op1, 
      JAL_op3, BRANCH_op1, LOAD_op, LOAD_op2, STORE_op1, STORE_op2, 
      FWD_A_mem_dec, FWD_A_exe_dec, FWD_A_wb_dec, FWD_A_sel_2_port, 
      FWD_A_sel_1_port, FWD_A_sel_0_port, FWD_B_mem_exe, FWD_B_exe_dec, 
      FWD_B_wb_dec, FWD_B_sel_2_port, FWD_B_sel_1_port, FWD_B_sel_0_port, 
      FWD_B_exe_mem, FWD_B_exe_mem1, FWD_B_exe_mem2, FWD_B_wb_mem, 
      FWD_B_wb_mem1, FWD_B_wb_mem2, FWD_B_mem_mem, FWD_B_mem_mem1, 
      FWD_B_mem_mem2, FWD_B_lmd1_mem, FWD_B_lmd1_mem1, FWD_B_lmd1_mem2, 
      FWD_exe_branch, FWD_exe_branch1, FWD_wb_branch, FWD_wb_branch1, net2664, 
      net2665, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n114
      , n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n97, n98, n99, n100, n101, n102, n113, n210, n312, n313, n314
      , n330, n331, n332, n424, n425, n426, n427, n428, n429, n430, n431, n432,
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454 : std_logic;

begin
   flush <= ( flush_1_port, flush_0_port );
   PC_out <= ( PC_out_31, PC_out_31, PC_out_31, PC_out_28_port, PC_out_27_port,
      PC_out_26_port, PC_out_25_port, PC_out_24_port, PC_out_23_port, 
      PC_out_22_port, PC_out_21_port, PC_out_20_port, PC_out_19_port, 
      PC_out_18_port, PC_out_17_port, PC_out_16_port, PC_out_15_port, 
      PC_out_14_port, PC_out_13_port, PC_out_12_port, PC_out_11_port, 
      PC_out_10_port, PC_out_9_port, PC_out_8_port, PC_out_7_port, 
      PC_out_6_port, PC_out_5_port, PC_out_4_port, PC_out_3_port, PC_out_2_port
      , PC_out_1_port, PC_out_0_port );
   
   ALU_block : alu port map( A(31) => ALU_operand_1_FWD_31_port, A(30) => 
                           ALU_operand_1_FWD_30_port, A(29) => 
                           ALU_operand_1_FWD_29_port, A(28) => 
                           ALU_operand_1_FWD_28_port, A(27) => 
                           ALU_operand_1_FWD_27_port, A(26) => 
                           ALU_operand_1_FWD_26_port, A(25) => 
                           ALU_operand_1_FWD_25_port, A(24) => 
                           ALU_operand_1_FWD_24_port, A(23) => 
                           ALU_operand_1_FWD_23_port, A(22) => 
                           ALU_operand_1_FWD_22_port, A(21) => 
                           ALU_operand_1_FWD_21_port, A(20) => 
                           ALU_operand_1_FWD_20_port, A(19) => 
                           ALU_operand_1_FWD_19_port, A(18) => 
                           ALU_operand_1_FWD_18_port, A(17) => 
                           ALU_operand_1_FWD_17_port, A(16) => 
                           ALU_operand_1_FWD_16_port, A(15) => 
                           ALU_operand_1_FWD_15_port, A(14) => 
                           ALU_operand_1_FWD_14_port, A(13) => 
                           ALU_operand_1_FWD_13_port, A(12) => 
                           ALU_operand_1_FWD_12_port, A(11) => 
                           ALU_operand_1_FWD_11_port, A(10) => 
                           ALU_operand_1_FWD_10_port, A(9) => 
                           ALU_operand_1_FWD_9_port, A(8) => 
                           ALU_operand_1_FWD_8_port, A(7) => 
                           ALU_operand_1_FWD_7_port, A(6) => 
                           ALU_operand_1_FWD_6_port, A(5) => 
                           ALU_operand_1_FWD_5_port, A(4) => 
                           ALU_operand_1_FWD_4_port, A(3) => 
                           ALU_operand_1_FWD_3_port, A(2) => 
                           ALU_operand_1_FWD_2_port, A(1) => 
                           ALU_operand_1_FWD_1_port, A(0) => 
                           ALU_operand_1_FWD_0_port, B(31) => 
                           ALU_operand_2_FWD_31_port, B(30) => 
                           ALU_operand_2_FWD_30_port, B(29) => 
                           ALU_operand_2_FWD_29_port, B(28) => 
                           ALU_operand_2_FWD_28_port, B(27) => 
                           ALU_operand_2_FWD_27_port, B(26) => 
                           ALU_operand_2_FWD_26_port, B(25) => 
                           ALU_operand_2_FWD_25_port, B(24) => 
                           ALU_operand_2_FWD_24_port, B(23) => 
                           ALU_operand_2_FWD_23_port, B(22) => 
                           ALU_operand_2_FWD_22_port, B(21) => 
                           ALU_operand_2_FWD_21_port, B(20) => 
                           ALU_operand_2_FWD_20_port, B(19) => 
                           ALU_operand_2_FWD_19_port, B(18) => 
                           ALU_operand_2_FWD_18_port, B(17) => 
                           ALU_operand_2_FWD_17_port, B(16) => 
                           ALU_operand_2_FWD_16_port, B(15) => 
                           ALU_operand_2_FWD_15_port, B(14) => 
                           ALU_operand_2_FWD_14_port, B(13) => 
                           ALU_operand_2_FWD_13_port, B(12) => 
                           ALU_operand_2_FWD_12_port, B(11) => 
                           ALU_operand_2_FWD_11_port, B(10) => 
                           ALU_operand_2_FWD_10_port, B(9) => 
                           ALU_operand_2_FWD_9_port, B(8) => 
                           ALU_operand_2_FWD_8_port, B(7) => 
                           ALU_operand_2_FWD_7_port, B(6) => 
                           ALU_operand_2_FWD_6_port, B(5) => 
                           ALU_operand_2_FWD_5_port, B(4) => 
                           ALU_operand_2_FWD_4_port, B(3) => 
                           ALU_operand_2_FWD_3_port, B(2) => 
                           ALU_operand_2_FWD_2_port, B(1) => 
                           ALU_operand_2_FWD_1_port, B(0) => 
                           ALU_operand_2_FWD_0_port, OP(0) => 
                           ALU_OPCODE_in_4_port, OP(1) => ALU_OPCODE_in_3_port,
                           OP(2) => ALU_OPCODE_in_2_port, OP(3) => 
                           ALU_OPCODE_in_1_port, OP(4) => ALU_OPCODE_in_0_port,
                           Y1(31) => ALU_output_31_port, Y1(30) => 
                           ALU_output_30_port, Y1(29) => ALU_output_29_port, 
                           Y1(28) => ALU_output_28_port, Y1(27) => 
                           ALU_output_27_port, Y1(26) => ALU_output_26_port, 
                           Y1(25) => ALU_output_25_port, Y1(24) => 
                           ALU_output_24_port, Y1(23) => ALU_output_23_port, 
                           Y1(22) => ALU_output_22_port, Y1(21) => 
                           ALU_output_21_port, Y1(20) => ALU_output_20_port, 
                           Y1(19) => ALU_output_19_port, Y1(18) => 
                           ALU_output_18_port, Y1(17) => ALU_output_17_port, 
                           Y1(16) => ALU_output_16_port, Y1(15) => 
                           ALU_output_15_port, Y1(14) => ALU_output_14_port, 
                           Y1(13) => ALU_output_13_port, Y1(12) => 
                           ALU_output_12_port, Y1(11) => ALU_output_11_port, 
                           Y1(10) => ALU_output_10_port, Y1(9) => 
                           ALU_output_9_port, Y1(8) => ALU_output_8_port, Y1(7)
                           => ALU_output_7_port, Y1(6) => ALU_output_6_port, 
                           Y1(5) => ALU_output_5_port, Y1(4) => 
                           ALU_output_4_port, Y1(3) => ALU_output_3_port, Y1(2)
                           => ALU_output_2_port, Y1(1) => ALU_output_1_port, 
                           Y1(0) => ALU_output_0_port, cout => net2665);
   jump_adder : cla_adder_N32 port map( A(31) => NPC_31_port, A(30) => 
                           NPC_30_port, A(29) => NPC_29_port, A(28) => 
                           NPC_28_port, A(27) => NPC_27_port, A(26) => 
                           NPC_26_port, A(25) => NPC_25_port, A(24) => 
                           NPC_24_port, A(23) => NPC_23_port, A(22) => 
                           NPC_22_port, A(21) => NPC_21_port, A(20) => 
                           NPC_20_port, A(19) => NPC_19_port, A(18) => 
                           NPC_18_port, A(17) => NPC_17_port, A(16) => 
                           NPC_16_port, A(15) => NPC_15_port, A(14) => 
                           NPC_14_port, A(13) => NPC_13_port, A(12) => 
                           NPC_12_port, A(11) => NPC_11_port, A(10) => 
                           NPC_10_port, A(9) => NPC_9_port, A(8) => NPC_8_port,
                           A(7) => NPC_7_port, A(6) => NPC_6_port, A(5) => 
                           NPC_5_port, A(4) => NPC_4_port, A(3) => NPC_3_port, 
                           A(2) => NPC_2_port, A(1) => NPC_1_port, A(0) => 
                           NPC_0_port, B(31) => 
                           PC_Immediate_displacement_31_port, B(30) => 
                           PC_Immediate_displacement_31_port, B(29) => 
                           PC_Immediate_displacement_31_port, B(28) => 
                           PC_Immediate_displacement_31_port, B(27) => 
                           PC_Immediate_displacement_31_port, B(26) => 
                           PC_Immediate_displacement_31_port, B(25) => 
                           PC_Immediate_displacement_31_port, B(24) => 
                           PC_Immediate_displacement_24_port, B(23) => 
                           PC_Immediate_displacement_23_port, B(22) => 
                           PC_Immediate_displacement_22_port, B(21) => 
                           PC_Immediate_displacement_21_port, B(20) => 
                           PC_Immediate_displacement_20_port, B(19) => 
                           PC_Immediate_displacement_19_port, B(18) => 
                           PC_Immediate_displacement_18_port, B(17) => 
                           PC_Immediate_displacement_17_port, B(16) => 
                           PC_Immediate_displacement_16_port, B(15) => 
                           Instr(15), B(14) => Instr(14), B(13) => Instr(13), 
                           B(12) => Instr(12), B(11) => Instr(11), B(10) => 
                           Instr(10), B(9) => Instr(9), B(8) => Instr(8), B(7) 
                           => Instr(7), B(6) => Instr(6), B(5) => Instr(5), 
                           B(4) => Instr(4), B(3) => Instr(3), B(2) => Instr(2)
                           , B(1) => Instr(1), B(0) => Instr(0), Ci => 
                           X_Logic0_port, Cout => net2664, Sum(31) => 
                           PC_displaced_31_port, Sum(30) => 
                           PC_displaced_30_port, Sum(29) => 
                           PC_displaced_29_port, Sum(28) => 
                           PC_displaced_28_port, Sum(27) => 
                           PC_displaced_27_port, Sum(26) => 
                           PC_displaced_26_port, Sum(25) => 
                           PC_displaced_25_port, Sum(24) => 
                           PC_displaced_24_port, Sum(23) => 
                           PC_displaced_23_port, Sum(22) => 
                           PC_displaced_22_port, Sum(21) => 
                           PC_displaced_21_port, Sum(20) => 
                           PC_displaced_20_port, Sum(19) => 
                           PC_displaced_19_port, Sum(18) => 
                           PC_displaced_18_port, Sum(17) => 
                           PC_displaced_17_port, Sum(16) => 
                           PC_displaced_16_port, Sum(15) => 
                           PC_displaced_15_port, Sum(14) => 
                           PC_displaced_14_port, Sum(13) => 
                           PC_displaced_13_port, Sum(12) => 
                           PC_displaced_12_port, Sum(11) => 
                           PC_displaced_11_port, Sum(10) => 
                           PC_displaced_10_port, Sum(9) => PC_displaced_9_port,
                           Sum(8) => PC_displaced_8_port, Sum(7) => 
                           PC_displaced_7_port, Sum(6) => PC_displaced_6_port, 
                           Sum(5) => PC_displaced_5_port, Sum(4) => 
                           PC_displaced_4_port, Sum(3) => PC_displaced_3_port, 
                           Sum(2) => PC_displaced_2_port, Sum(1) => 
                           PC_displaced_1_port, Sum(0) => PC_displaced_0_port);
   X_Logic0_port <= '0';
   U456 : NAND3_X1 port map( A1 => Instr_reg_out_31_port, A2 => 
                           Instr_reg_out_29_port, A3 => n228, ZN => n109);
   U457 : OAI33_X1 port map( A1 => n232, A2 => FWD_exe_branch1, A3 => n233, B1 
                           => n234, B2 => n235, B3 => n236, ZN => n231);
   U458 : NAND3_X1 port map( A1 => n297, A2 => n298, A3 => n299, ZN => n296);
   U459 : NAND3_X1 port map( A1 => Instr_reg_out_27_port, A2 => n278, A3 => 
                           Instr_reg_out_26_port, ZN => n311);
   U460 : NAND3_X1 port map( A1 => n306, A2 => n307, A3 => n305, ZN => n327);
   U461 : XOR2_X1 port map( A => RD2_0_port, B => Instr_reg_out_21_port, Z => 
                           n341);
   U462 : XOR2_X1 port map( A => RD2_1_port, B => Instr_reg_out_22_port, Z => 
                           n340);
   U463 : XOR2_X1 port map( A => RD1_0_port, B => Instr_reg_out_21_port, Z => 
                           n349);
   U464 : XOR2_X1 port map( A => RD1_1_port, B => Instr_reg_out_22_port, Z => 
                           n348);
   IR : reg_N32_0 port map( clk => Clk, rst => n451, d_in(31) => Instr(31), 
                           d_in(30) => Instr(30), d_in(29) => Instr(29), 
                           d_in(28) => Instr(28), d_in(27) => Instr(27), 
                           d_in(26) => Instr(26), d_in(25) => Instr(25), 
                           d_in(24) => Instr(24), d_in(23) => Instr(23), 
                           d_in(22) => Instr(22), d_in(21) => Instr(21), 
                           d_in(20) => Instr(20), d_in(19) => Instr(19), 
                           d_in(18) => Instr(18), d_in(17) => Instr(17), 
                           d_in(16) => Instr(16), d_in(15) => Instr(15), 
                           d_in(14) => Instr(14), d_in(13) => Instr(13), 
                           d_in(12) => Instr(12), d_in(11) => Instr(11), 
                           d_in(10) => Instr(10), d_in(9) => Instr(9), d_in(8) 
                           => Instr(8), d_in(7) => Instr(7), d_in(6) => 
                           Instr(6), d_in(5) => Instr(5), d_in(4) => Instr(4), 
                           d_in(3) => Instr(3), d_in(2) => Instr(2), d_in(1) =>
                           Instr(1), d_in(0) => Instr(0), d_out(31) => 
                           Instr_reg_out_31_port, d_out(30) => 
                           Instr_reg_out_30_port, d_out(29) => 
                           Instr_reg_out_29_port, d_out(28) => 
                           Instr_reg_out_28_port, d_out(27) => 
                           Instr_reg_out_27_port, d_out(26) => 
                           Instr_reg_out_26_port, d_out(25) => 
                           Instr_reg_out_25_port, d_out(24) => 
                           Instr_reg_out_24_port, d_out(23) => 
                           Instr_reg_out_23_port, d_out(22) => 
                           Instr_reg_out_22_port, d_out(21) => 
                           Instr_reg_out_21_port, d_out(20) => 
                           Instr_reg_out_20_port, d_out(19) => 
                           Instr_reg_out_19_port, d_out(18) => 
                           Instr_reg_out_18_port, d_out(17) => 
                           Instr_reg_out_17_port, d_out(16) => 
                           Instr_reg_out_16_port, d_out(15) => 
                           Instr_reg_out_15_port, d_out(14) => 
                           Instr_reg_out_14_port, d_out(13) => 
                           Instr_reg_out_13_port, d_out(12) => 
                           Instr_reg_out_12_port, d_out(11) => 
                           Instr_reg_out_11_port, d_out(10) => 
                           Instr_reg_out_10_port, d_out(9) => 
                           Instr_reg_out_9_port, d_out(8) => 
                           Instr_reg_out_8_port, d_out(7) => 
                           Instr_reg_out_7_port, d_out(6) => 
                           Instr_reg_out_6_port, d_out(5) => 
                           Instr_reg_out_5_port, d_out(4) => 
                           Instr_reg_out_4_port, d_out(3) => 
                           Instr_reg_out_3_port, d_out(2) => 
                           Instr_reg_out_2_port, d_out(1) => 
                           Instr_reg_out_1_port, d_out(0) => 
                           Instr_reg_out_0_port);
   OPC1 : reg_N6_0 port map( clk => Clk, rst => n451, d_in(5) => 
                           Instr_reg_out_31_port, d_in(4) => 
                           Instr_reg_out_30_port, d_in(3) => 
                           Instr_reg_out_29_port, d_in(2) => 
                           Instr_reg_out_28_port, d_in(1) => 
                           Instr_reg_out_27_port, d_in(0) => 
                           Instr_reg_out_26_port, d_out(5) => OPCODE1_5_port, 
                           d_out(4) => OPCODE1_4_port, d_out(3) => 
                           OPCODE1_3_port, d_out(2) => OPCODE1_2_port, d_out(1)
                           => OPCODE1_1_port, d_out(0) => OPCODE1_0_port);
   OPC2 : reg_N6_1 port map( clk => Clk, rst => n451, d_in(5) => OPCODE1_5_port
                           , d_in(4) => OPCODE1_4_port, d_in(3) => 
                           OPCODE1_3_port, d_in(2) => OPCODE1_2_port, d_in(1) 
                           => OPCODE1_1_port, d_in(0) => OPCODE1_0_port, 
                           d_out(5) => OPCODE2_5_port, d_out(4) => 
                           OPCODE2_4_port, d_out(3) => OPCODE2_3_port, d_out(2)
                           => OPCODE2_2_port, d_out(1) => OPCODE2_1_port, 
                           d_out(0) => OPCODE2_0_port);
   RDreg1 : reg_N5_0 port map( clk => Clk, rst => n451, d_in(4) => RD_4_port, 
                           d_in(3) => RD_3_port, d_in(2) => RD_2_port, d_in(1) 
                           => RD_1_port, d_in(0) => RD_0_port, d_out(4) => 
                           RD1_4_port, d_out(3) => RD1_3_port, d_out(2) => 
                           RD1_2_port, d_out(1) => RD1_1_port, d_out(0) => 
                           RD1_0_port);
   RDreg2 : reg_N5_2 port map( clk => Clk, rst => n451, d_in(4) => RD1_4_port, 
                           d_in(3) => RD1_3_port, d_in(2) => RD1_2_port, 
                           d_in(1) => RD1_1_port, d_in(0) => RD1_0_port, 
                           d_out(4) => RD2_4_port, d_out(3) => RD2_3_port, 
                           d_out(2) => RD2_2_port, d_out(1) => RD2_1_port, 
                           d_out(0) => RD2_0_port);
   RDreg3 : reg_N5_1 port map( clk => Clk, rst => n451, d_in(4) => RD2_4_port, 
                           d_in(3) => RD2_3_port, d_in(2) => RD2_2_port, 
                           d_in(1) => RD2_1_port, d_in(0) => RD2_0_port, 
                           d_out(4) => RD3_4_port, d_out(3) => RD3_3_port, 
                           d_out(2) => RD3_2_port, d_out(1) => RD3_1_port, 
                           d_out(0) => RD3_0_port);
   RF : w_reg_file_M8_N8_F4_Nbit32 port map( clk => Clk, reset => n451, enable 
                           => RF_EN, rd1 => RF_RD1_EN, rd2 => RF_RD2_EN, wr => 
                           RF_WR, add_wr(4) => RD3_4_port, add_wr(3) => 
                           RD3_3_port, add_wr(2) => RD3_2_port, add_wr(1) => 
                           RD3_1_port, add_wr(0) => RD3_0_port, add_rd1(4) => 
                           Instr_reg_out_25_port, add_rd1(3) => 
                           Instr_reg_out_24_port, add_rd1(2) => 
                           Instr_reg_out_23_port, add_rd1(1) => 
                           Instr_reg_out_22_port, add_rd1(0) => 
                           Instr_reg_out_21_port, add_rd2(4) => 
                           Instr_reg_out_20_port, add_rd2(3) => 
                           Instr_reg_out_19_port, add_rd2(2) => 
                           Instr_reg_out_18_port, add_rd2(1) => 
                           Instr_reg_out_17_port, add_rd2(0) => 
                           Instr_reg_out_16_port, datain(31) => 
                           RF_write_data_31_port, datain(30) => 
                           RF_write_data_30_port, datain(29) => 
                           RF_write_data_29_port, datain(28) => 
                           RF_write_data_28_port, datain(27) => 
                           RF_write_data_27_port, datain(26) => 
                           RF_write_data_26_port, datain(25) => 
                           RF_write_data_25_port, datain(24) => 
                           RF_write_data_24_port, datain(23) => 
                           RF_write_data_23_port, datain(22) => 
                           RF_write_data_22_port, datain(21) => 
                           RF_write_data_21_port, datain(20) => 
                           RF_write_data_20_port, datain(19) => 
                           RF_write_data_19_port, datain(18) => 
                           RF_write_data_18_port, datain(17) => 
                           RF_write_data_17_port, datain(16) => 
                           RF_write_data_16_port, datain(15) => 
                           RF_write_data_15_port, datain(14) => 
                           RF_write_data_14_port, datain(13) => 
                           RF_write_data_13_port, datain(12) => 
                           RF_write_data_12_port, datain(11) => 
                           RF_write_data_11_port, datain(10) => 
                           RF_write_data_10_port, datain(9) => 
                           RF_write_data_9_port, datain(8) => 
                           RF_write_data_8_port, datain(7) => 
                           RF_write_data_7_port, datain(6) => 
                           RF_write_data_6_port, datain(5) => 
                           RF_write_data_5_port, datain(4) => 
                           RF_write_data_4_port, datain(3) => 
                           RF_write_data_3_port, datain(2) => 
                           RF_write_data_2_port, datain(1) => 
                           RF_write_data_1_port, datain(0) => 
                           RF_write_data_0_port, out1(31) => RF_out_A_31_port, 
                           out1(30) => RF_out_A_30_port, out1(29) => 
                           RF_out_A_29_port, out1(28) => RF_out_A_28_port, 
                           out1(27) => RF_out_A_27_port, out1(26) => 
                           RF_out_A_26_port, out1(25) => RF_out_A_25_port, 
                           out1(24) => RF_out_A_24_port, out1(23) => 
                           RF_out_A_23_port, out1(22) => RF_out_A_22_port, 
                           out1(21) => RF_out_A_21_port, out1(20) => 
                           RF_out_A_20_port, out1(19) => RF_out_A_19_port, 
                           out1(18) => RF_out_A_18_port, out1(17) => 
                           RF_out_A_17_port, out1(16) => RF_out_A_16_port, 
                           out1(15) => RF_out_A_15_port, out1(14) => 
                           RF_out_A_14_port, out1(13) => RF_out_A_13_port, 
                           out1(12) => RF_out_A_12_port, out1(11) => 
                           RF_out_A_11_port, out1(10) => RF_out_A_10_port, 
                           out1(9) => RF_out_A_9_port, out1(8) => 
                           RF_out_A_8_port, out1(7) => RF_out_A_7_port, out1(6)
                           => RF_out_A_6_port, out1(5) => RF_out_A_5_port, 
                           out1(4) => RF_out_A_4_port, out1(3) => 
                           RF_out_A_3_port, out1(2) => RF_out_A_2_port, out1(1)
                           => RF_out_A_1_port, out1(0) => RF_out_A_0_port, 
                           out2(31) => RF_out_B_31_port, out2(30) => 
                           RF_out_B_30_port, out2(29) => RF_out_B_29_port, 
                           out2(28) => RF_out_B_28_port, out2(27) => 
                           RF_out_B_27_port, out2(26) => RF_out_B_26_port, 
                           out2(25) => RF_out_B_25_port, out2(24) => 
                           RF_out_B_24_port, out2(23) => RF_out_B_23_port, 
                           out2(22) => RF_out_B_22_port, out2(21) => 
                           RF_out_B_21_port, out2(20) => RF_out_B_20_port, 
                           out2(19) => RF_out_B_19_port, out2(18) => 
                           RF_out_B_18_port, out2(17) => RF_out_B_17_port, 
                           out2(16) => RF_out_B_16_port, out2(15) => 
                           RF_out_B_15_port, out2(14) => RF_out_B_14_port, 
                           out2(13) => RF_out_B_13_port, out2(12) => 
                           RF_out_B_12_port, out2(11) => RF_out_B_11_port, 
                           out2(10) => RF_out_B_10_port, out2(9) => 
                           RF_out_B_9_port, out2(8) => RF_out_B_8_port, out2(7)
                           => RF_out_B_7_port, out2(6) => RF_out_B_6_port, 
                           out2(5) => RF_out_B_5_port, out2(4) => 
                           RF_out_B_4_port, out2(3) => RF_out_B_3_port, out2(2)
                           => RF_out_B_2_port, out2(1) => RF_out_B_1_port, 
                           out2(0) => RF_out_B_0_port, call => CALL, ret => RET
                           , spill => SPILL, fill => FILL, to_mem(31) => 
                           spill_to_stack_31_port, to_mem(30) => 
                           spill_to_stack_30_port, to_mem(29) => 
                           spill_to_stack_29_port, to_mem(28) => 
                           spill_to_stack_28_port, to_mem(27) => 
                           spill_to_stack_27_port, to_mem(26) => 
                           spill_to_stack_26_port, to_mem(25) => 
                           spill_to_stack_25_port, to_mem(24) => 
                           spill_to_stack_24_port, to_mem(23) => 
                           spill_to_stack_23_port, to_mem(22) => 
                           spill_to_stack_22_port, to_mem(21) => 
                           spill_to_stack_21_port, to_mem(20) => 
                           spill_to_stack_20_port, to_mem(19) => 
                           spill_to_stack_19_port, to_mem(18) => 
                           spill_to_stack_18_port, to_mem(17) => 
                           spill_to_stack_17_port, to_mem(16) => 
                           spill_to_stack_16_port, to_mem(15) => 
                           spill_to_stack_15_port, to_mem(14) => 
                           spill_to_stack_14_port, to_mem(13) => 
                           spill_to_stack_13_port, to_mem(12) => 
                           spill_to_stack_12_port, to_mem(11) => 
                           spill_to_stack_11_port, to_mem(10) => 
                           spill_to_stack_10_port, to_mem(9) => 
                           spill_to_stack_9_port, to_mem(8) => 
                           spill_to_stack_8_port, to_mem(7) => 
                           spill_to_stack_7_port, to_mem(6) => 
                           spill_to_stack_6_port, to_mem(5) => 
                           spill_to_stack_5_port, to_mem(4) => 
                           spill_to_stack_4_port, to_mem(3) => 
                           spill_to_stack_3_port, to_mem(2) => 
                           spill_to_stack_2_port, to_mem(1) => 
                           spill_to_stack_1_port, to_mem(0) => 
                           spill_to_stack_0_port, from_mem(31) => 
                           fill_from_stack_31_port, from_mem(30) => 
                           fill_from_stack_30_port, from_mem(29) => 
                           fill_from_stack_29_port, from_mem(28) => 
                           fill_from_stack_28_port, from_mem(27) => 
                           fill_from_stack_27_port, from_mem(26) => 
                           fill_from_stack_26_port, from_mem(25) => 
                           fill_from_stack_25_port, from_mem(24) => 
                           fill_from_stack_24_port, from_mem(23) => 
                           fill_from_stack_23_port, from_mem(22) => 
                           fill_from_stack_22_port, from_mem(21) => 
                           fill_from_stack_21_port, from_mem(20) => 
                           fill_from_stack_20_port, from_mem(19) => 
                           fill_from_stack_19_port, from_mem(18) => 
                           fill_from_stack_18_port, from_mem(17) => 
                           fill_from_stack_17_port, from_mem(16) => 
                           fill_from_stack_16_port, from_mem(15) => 
                           fill_from_stack_15_port, from_mem(14) => 
                           fill_from_stack_14_port, from_mem(13) => 
                           fill_from_stack_13_port, from_mem(12) => 
                           fill_from_stack_12_port, from_mem(11) => 
                           fill_from_stack_11_port, from_mem(10) => 
                           fill_from_stack_10_port, from_mem(9) => 
                           fill_from_stack_9_port, from_mem(8) => 
                           fill_from_stack_8_port, from_mem(7) => 
                           fill_from_stack_7_port, from_mem(6) => 
                           fill_from_stack_6_port, from_mem(5) => 
                           fill_from_stack_5_port, from_mem(4) => 
                           fill_from_stack_4_port, from_mem(3) => 
                           fill_from_stack_3_port, from_mem(2) => 
                           fill_from_stack_2_port, from_mem(1) => 
                           fill_from_stack_1_port, from_mem(0) => 
                           fill_from_stack_0_port);
   WRF_stack : stack port map( clk => Clk, reset => n453, enable => n454, RD =>
                           FILL, wr => SPILL, datain(31) => 
                           spill_to_stack_31_port, datain(30) => 
                           spill_to_stack_30_port, datain(29) => 
                           spill_to_stack_29_port, datain(28) => 
                           spill_to_stack_28_port, datain(27) => 
                           spill_to_stack_27_port, datain(26) => 
                           spill_to_stack_26_port, datain(25) => 
                           spill_to_stack_25_port, datain(24) => 
                           spill_to_stack_24_port, datain(23) => 
                           spill_to_stack_23_port, datain(22) => 
                           spill_to_stack_22_port, datain(21) => 
                           spill_to_stack_21_port, datain(20) => 
                           spill_to_stack_20_port, datain(19) => 
                           spill_to_stack_19_port, datain(18) => 
                           spill_to_stack_18_port, datain(17) => 
                           spill_to_stack_17_port, datain(16) => 
                           spill_to_stack_16_port, datain(15) => 
                           spill_to_stack_15_port, datain(14) => 
                           spill_to_stack_14_port, datain(13) => 
                           spill_to_stack_13_port, datain(12) => 
                           spill_to_stack_12_port, datain(11) => 
                           spill_to_stack_11_port, datain(10) => 
                           spill_to_stack_10_port, datain(9) => 
                           spill_to_stack_9_port, datain(8) => 
                           spill_to_stack_8_port, datain(7) => 
                           spill_to_stack_7_port, datain(6) => 
                           spill_to_stack_6_port, datain(5) => 
                           spill_to_stack_5_port, datain(4) => 
                           spill_to_stack_4_port, datain(3) => 
                           spill_to_stack_3_port, datain(2) => 
                           spill_to_stack_2_port, datain(1) => 
                           spill_to_stack_1_port, datain(0) => 
                           spill_to_stack_0_port, dataout(31) => 
                           fill_from_stack_31_port, dataout(30) => 
                           fill_from_stack_30_port, dataout(29) => 
                           fill_from_stack_29_port, dataout(28) => 
                           fill_from_stack_28_port, dataout(27) => 
                           fill_from_stack_27_port, dataout(26) => 
                           fill_from_stack_26_port, dataout(25) => 
                           fill_from_stack_25_port, dataout(24) => 
                           fill_from_stack_24_port, dataout(23) => 
                           fill_from_stack_23_port, dataout(22) => 
                           fill_from_stack_22_port, dataout(21) => 
                           fill_from_stack_21_port, dataout(20) => 
                           fill_from_stack_20_port, dataout(19) => 
                           fill_from_stack_19_port, dataout(18) => 
                           fill_from_stack_18_port, dataout(17) => 
                           fill_from_stack_17_port, dataout(16) => 
                           fill_from_stack_16_port, dataout(15) => 
                           fill_from_stack_15_port, dataout(14) => 
                           fill_from_stack_14_port, dataout(13) => 
                           fill_from_stack_13_port, dataout(12) => 
                           fill_from_stack_12_port, dataout(11) => 
                           fill_from_stack_11_port, dataout(10) => 
                           fill_from_stack_10_port, dataout(9) => 
                           fill_from_stack_9_port, dataout(8) => 
                           fill_from_stack_8_port, dataout(7) => 
                           fill_from_stack_7_port, dataout(6) => 
                           fill_from_stack_6_port, dataout(5) => 
                           fill_from_stack_5_port, dataout(4) => 
                           fill_from_stack_4_port, dataout(3) => 
                           fill_from_stack_3_port, dataout(2) => 
                           fill_from_stack_2_port, dataout(1) => 
                           fill_from_stack_1_port, dataout(0) => 
                           fill_from_stack_0_port);
   A : reg_N32_13 port map( clk => Clk, rst => n451, d_in(31) => 
                           RF_out_A_31_port, d_in(30) => RF_out_A_30_port, 
                           d_in(29) => RF_out_A_29_port, d_in(28) => 
                           RF_out_A_28_port, d_in(27) => RF_out_A_27_port, 
                           d_in(26) => RF_out_A_26_port, d_in(25) => 
                           RF_out_A_25_port, d_in(24) => RF_out_A_24_port, 
                           d_in(23) => RF_out_A_23_port, d_in(22) => 
                           RF_out_A_22_port, d_in(21) => RF_out_A_21_port, 
                           d_in(20) => RF_out_A_20_port, d_in(19) => 
                           RF_out_A_19_port, d_in(18) => RF_out_A_18_port, 
                           d_in(17) => RF_out_A_17_port, d_in(16) => 
                           RF_out_A_16_port, d_in(15) => RF_out_A_15_port, 
                           d_in(14) => RF_out_A_14_port, d_in(13) => 
                           RF_out_A_13_port, d_in(12) => RF_out_A_12_port, 
                           d_in(11) => RF_out_A_11_port, d_in(10) => 
                           RF_out_A_10_port, d_in(9) => RF_out_A_9_port, 
                           d_in(8) => RF_out_A_8_port, d_in(7) => 
                           RF_out_A_7_port, d_in(6) => RF_out_A_6_port, d_in(5)
                           => RF_out_A_5_port, d_in(4) => RF_out_A_4_port, 
                           d_in(3) => RF_out_A_3_port, d_in(2) => 
                           RF_out_A_2_port, d_in(1) => RF_out_A_1_port, d_in(0)
                           => RF_out_A_0_port, d_out(31) => A_reg_out_31_port, 
                           d_out(30) => A_reg_out_30_port, d_out(29) => 
                           A_reg_out_29_port, d_out(28) => A_reg_out_28_port, 
                           d_out(27) => A_reg_out_27_port, d_out(26) => 
                           A_reg_out_26_port, d_out(25) => A_reg_out_25_port, 
                           d_out(24) => A_reg_out_24_port, d_out(23) => 
                           A_reg_out_23_port, d_out(22) => A_reg_out_22_port, 
                           d_out(21) => A_reg_out_21_port, d_out(20) => 
                           A_reg_out_20_port, d_out(19) => A_reg_out_19_port, 
                           d_out(18) => A_reg_out_18_port, d_out(17) => 
                           A_reg_out_17_port, d_out(16) => A_reg_out_16_port, 
                           d_out(15) => A_reg_out_15_port, d_out(14) => 
                           A_reg_out_14_port, d_out(13) => A_reg_out_13_port, 
                           d_out(12) => A_reg_out_12_port, d_out(11) => 
                           A_reg_out_11_port, d_out(10) => A_reg_out_10_port, 
                           d_out(9) => A_reg_out_9_port, d_out(8) => 
                           A_reg_out_8_port, d_out(7) => A_reg_out_7_port, 
                           d_out(6) => A_reg_out_6_port, d_out(5) => 
                           A_reg_out_5_port, d_out(4) => A_reg_out_4_port, 
                           d_out(3) => A_reg_out_3_port, d_out(2) => 
                           A_reg_out_2_port, d_out(1) => A_reg_out_1_port, 
                           d_out(0) => A_reg_out_0_port);
   B : reg_N32_12 port map( clk => Clk, rst => n452, d_in(31) => 
                           RF_out_B_31_port, d_in(30) => RF_out_B_30_port, 
                           d_in(29) => RF_out_B_29_port, d_in(28) => 
                           RF_out_B_28_port, d_in(27) => RF_out_B_27_port, 
                           d_in(26) => RF_out_B_26_port, d_in(25) => 
                           RF_out_B_25_port, d_in(24) => RF_out_B_24_port, 
                           d_in(23) => RF_out_B_23_port, d_in(22) => 
                           RF_out_B_22_port, d_in(21) => RF_out_B_21_port, 
                           d_in(20) => RF_out_B_20_port, d_in(19) => 
                           RF_out_B_19_port, d_in(18) => RF_out_B_18_port, 
                           d_in(17) => RF_out_B_17_port, d_in(16) => 
                           RF_out_B_16_port, d_in(15) => RF_out_B_15_port, 
                           d_in(14) => RF_out_B_14_port, d_in(13) => 
                           RF_out_B_13_port, d_in(12) => RF_out_B_12_port, 
                           d_in(11) => RF_out_B_11_port, d_in(10) => 
                           RF_out_B_10_port, d_in(9) => RF_out_B_9_port, 
                           d_in(8) => RF_out_B_8_port, d_in(7) => 
                           RF_out_B_7_port, d_in(6) => RF_out_B_6_port, d_in(5)
                           => RF_out_B_5_port, d_in(4) => RF_out_B_4_port, 
                           d_in(3) => RF_out_B_3_port, d_in(2) => 
                           RF_out_B_2_port, d_in(1) => RF_out_B_1_port, d_in(0)
                           => RF_out_B_0_port, d_out(31) => B_reg_out_31_port, 
                           d_out(30) => B_reg_out_30_port, d_out(29) => 
                           B_reg_out_29_port, d_out(28) => B_reg_out_28_port, 
                           d_out(27) => B_reg_out_27_port, d_out(26) => 
                           B_reg_out_26_port, d_out(25) => B_reg_out_25_port, 
                           d_out(24) => B_reg_out_24_port, d_out(23) => 
                           B_reg_out_23_port, d_out(22) => B_reg_out_22_port, 
                           d_out(21) => B_reg_out_21_port, d_out(20) => 
                           B_reg_out_20_port, d_out(19) => B_reg_out_19_port, 
                           d_out(18) => B_reg_out_18_port, d_out(17) => 
                           B_reg_out_17_port, d_out(16) => B_reg_out_16_port, 
                           d_out(15) => B_reg_out_15_port, d_out(14) => 
                           B_reg_out_14_port, d_out(13) => B_reg_out_13_port, 
                           d_out(12) => B_reg_out_12_port, d_out(11) => 
                           B_reg_out_11_port, d_out(10) => B_reg_out_10_port, 
                           d_out(9) => B_reg_out_9_port, d_out(8) => 
                           B_reg_out_8_port, d_out(7) => B_reg_out_7_port, 
                           d_out(6) => B_reg_out_6_port, d_out(5) => 
                           B_reg_out_5_port, d_out(4) => B_reg_out_4_port, 
                           d_out(3) => B_reg_out_3_port, d_out(2) => 
                           B_reg_out_2_port, d_out(1) => B_reg_out_1_port, 
                           d_out(0) => B_reg_out_0_port);
   Imm16ext : sign_ext_Nstart16_Nend32 port map( Ain(15) => 
                           Instr_reg_out_15_port, Ain(14) => 
                           Instr_reg_out_14_port, Ain(13) => 
                           Instr_reg_out_13_port, Ain(12) => 
                           Instr_reg_out_12_port, Ain(11) => 
                           Instr_reg_out_11_port, Ain(10) => 
                           Instr_reg_out_10_port, Ain(9) => 
                           Instr_reg_out_9_port, Ain(8) => Instr_reg_out_8_port
                           , Ain(7) => Instr_reg_out_7_port, Ain(6) => 
                           Instr_reg_out_6_port, Ain(5) => Instr_reg_out_5_port
                           , Ain(4) => Instr_reg_out_4_port, Ain(3) => 
                           Instr_reg_out_3_port, Ain(2) => Instr_reg_out_2_port
                           , Ain(1) => Instr_reg_out_1_port, Ain(0) => 
                           Instr_reg_out_0_port, Aout(31) => 
                           Immediate_16_extended_31_port, Aout(30) => 
                           Immediate_16_extended_30_port, Aout(29) => 
                           Immediate_16_extended_29_port, Aout(28) => 
                           Immediate_16_extended_28_port, Aout(27) => 
                           Immediate_16_extended_27_port, Aout(26) => 
                           Immediate_16_extended_26_port, Aout(25) => 
                           Immediate_16_extended_25_port, Aout(24) => 
                           Immediate_16_extended_24_port, Aout(23) => 
                           Immediate_16_extended_23_port, Aout(22) => 
                           Immediate_16_extended_22_port, Aout(21) => 
                           Immediate_16_extended_21_port, Aout(20) => 
                           Immediate_16_extended_20_port, Aout(19) => 
                           Immediate_16_extended_19_port, Aout(18) => 
                           Immediate_16_extended_18_port, Aout(17) => 
                           Immediate_16_extended_17_port, Aout(16) => 
                           Immediate_16_extended_16_port, Aout(15) => 
                           Immediate_16_extended_15_port, Aout(14) => 
                           Immediate_16_extended_14_port, Aout(13) => 
                           Immediate_16_extended_13_port, Aout(12) => 
                           Immediate_16_extended_12_port, Aout(11) => 
                           Immediate_16_extended_11_port, Aout(10) => 
                           Immediate_16_extended_10_port, Aout(9) => 
                           Immediate_16_extended_9_port, Aout(8) => 
                           Immediate_16_extended_8_port, Aout(7) => 
                           Immediate_16_extended_7_port, Aout(6) => 
                           Immediate_16_extended_6_port, Aout(5) => 
                           Immediate_16_extended_5_port, Aout(4) => 
                           Immediate_16_extended_4_port, Aout(3) => 
                           Immediate_16_extended_3_port, Aout(2) => 
                           Immediate_16_extended_2_port, Aout(1) => 
                           Immediate_16_extended_1_port, Aout(0) => 
                           Immediate_16_extended_0_port);
   Imm26ext : sign_ext_Nstart26_Nend32 port map( Ain(25) => 
                           Instr_reg_out_25_port, Ain(24) => 
                           Instr_reg_out_24_port, Ain(23) => 
                           Instr_reg_out_23_port, Ain(22) => 
                           Instr_reg_out_22_port, Ain(21) => 
                           Instr_reg_out_21_port, Ain(20) => 
                           Instr_reg_out_20_port, Ain(19) => 
                           Instr_reg_out_19_port, Ain(18) => 
                           Instr_reg_out_18_port, Ain(17) => 
                           Instr_reg_out_17_port, Ain(16) => 
                           Instr_reg_out_16_port, Ain(15) => 
                           Instr_reg_out_15_port, Ain(14) => 
                           Instr_reg_out_14_port, Ain(13) => 
                           Instr_reg_out_13_port, Ain(12) => 
                           Instr_reg_out_12_port, Ain(11) => 
                           Instr_reg_out_11_port, Ain(10) => 
                           Instr_reg_out_10_port, Ain(9) => 
                           Instr_reg_out_9_port, Ain(8) => Instr_reg_out_8_port
                           , Ain(7) => Instr_reg_out_7_port, Ain(6) => 
                           Instr_reg_out_6_port, Ain(5) => Instr_reg_out_5_port
                           , Ain(4) => Instr_reg_out_4_port, Ain(3) => 
                           Instr_reg_out_3_port, Ain(2) => Instr_reg_out_2_port
                           , Ain(1) => Instr_reg_out_1_port, Ain(0) => 
                           Instr_reg_out_0_port, Aout(31) => 
                           Immediate_26_extended_31_port, Aout(30) => 
                           Immediate_26_extended_30_port, Aout(29) => 
                           Immediate_26_extended_29_port, Aout(28) => 
                           Immediate_26_extended_28_port, Aout(27) => 
                           Immediate_26_extended_27_port, Aout(26) => 
                           Immediate_26_extended_26_port, Aout(25) => 
                           Immediate_26_extended_25_port, Aout(24) => 
                           Immediate_26_extended_24_port, Aout(23) => 
                           Immediate_26_extended_23_port, Aout(22) => 
                           Immediate_26_extended_22_port, Aout(21) => 
                           Immediate_26_extended_21_port, Aout(20) => 
                           Immediate_26_extended_20_port, Aout(19) => 
                           Immediate_26_extended_19_port, Aout(18) => 
                           Immediate_26_extended_18_port, Aout(17) => 
                           Immediate_26_extended_17_port, Aout(16) => 
                           Immediate_26_extended_16_port, Aout(15) => 
                           Immediate_26_extended_15_port, Aout(14) => 
                           Immediate_26_extended_14_port, Aout(13) => 
                           Immediate_26_extended_13_port, Aout(12) => 
                           Immediate_26_extended_12_port, Aout(11) => 
                           Immediate_26_extended_11_port, Aout(10) => 
                           Immediate_26_extended_10_port, Aout(9) => 
                           Immediate_26_extended_9_port, Aout(8) => 
                           Immediate_26_extended_8_port, Aout(7) => 
                           Immediate_26_extended_7_port, Aout(6) => 
                           Immediate_26_extended_6_port, Aout(5) => 
                           Immediate_26_extended_5_port, Aout(4) => 
                           Immediate_26_extended_4_port, Aout(3) => 
                           Immediate_26_extended_3_port, Aout(2) => 
                           Immediate_26_extended_2_port, Aout(1) => 
                           Immediate_26_extended_1_port, Aout(0) => 
                           Immediate_26_extended_0_port);
   mux_imm : MUX21_GENERIC_N32_0 port map( A(31) => 
                           Immediate_16_extended_31_port, A(30) => 
                           Immediate_16_extended_30_port, A(29) => 
                           Immediate_16_extended_29_port, A(28) => 
                           Immediate_16_extended_28_port, A(27) => 
                           Immediate_16_extended_27_port, A(26) => 
                           Immediate_16_extended_26_port, A(25) => 
                           Immediate_16_extended_25_port, A(24) => 
                           Immediate_16_extended_24_port, A(23) => 
                           Immediate_16_extended_23_port, A(22) => 
                           Immediate_16_extended_22_port, A(21) => 
                           Immediate_16_extended_21_port, A(20) => 
                           Immediate_16_extended_20_port, A(19) => 
                           Immediate_16_extended_19_port, A(18) => 
                           Immediate_16_extended_18_port, A(17) => 
                           Immediate_16_extended_17_port, A(16) => 
                           Immediate_16_extended_16_port, A(15) => 
                           Immediate_16_extended_15_port, A(14) => 
                           Immediate_16_extended_14_port, A(13) => 
                           Immediate_16_extended_13_port, A(12) => 
                           Immediate_16_extended_12_port, A(11) => 
                           Immediate_16_extended_11_port, A(10) => 
                           Immediate_16_extended_10_port, A(9) => 
                           Immediate_16_extended_9_port, A(8) => 
                           Immediate_16_extended_8_port, A(7) => 
                           Immediate_16_extended_7_port, A(6) => 
                           Immediate_16_extended_6_port, A(5) => 
                           Immediate_16_extended_5_port, A(4) => 
                           Immediate_16_extended_4_port, A(3) => 
                           Immediate_16_extended_3_port, A(2) => 
                           Immediate_16_extended_2_port, A(1) => 
                           Immediate_16_extended_1_port, A(0) => 
                           Immediate_16_extended_0_port, B(31) => 
                           Immediate_26_extended_31_port, B(30) => 
                           Immediate_26_extended_30_port, B(29) => 
                           Immediate_26_extended_29_port, B(28) => 
                           Immediate_26_extended_28_port, B(27) => 
                           Immediate_26_extended_27_port, B(26) => 
                           Immediate_26_extended_26_port, B(25) => 
                           Immediate_26_extended_25_port, B(24) => 
                           Immediate_26_extended_24_port, B(23) => 
                           Immediate_26_extended_23_port, B(22) => 
                           Immediate_26_extended_22_port, B(21) => 
                           Immediate_26_extended_21_port, B(20) => 
                           Immediate_26_extended_20_port, B(19) => 
                           Immediate_26_extended_19_port, B(18) => 
                           Immediate_26_extended_18_port, B(17) => 
                           Immediate_26_extended_17_port, B(16) => 
                           Immediate_26_extended_16_port, B(15) => 
                           Immediate_26_extended_15_port, B(14) => 
                           Immediate_26_extended_14_port, B(13) => 
                           Immediate_26_extended_13_port, B(12) => 
                           Immediate_26_extended_12_port, B(11) => 
                           Immediate_26_extended_11_port, B(10) => 
                           Immediate_26_extended_10_port, B(9) => 
                           Immediate_26_extended_9_port, B(8) => 
                           Immediate_26_extended_8_port, B(7) => 
                           Immediate_26_extended_7_port, B(6) => 
                           Immediate_26_extended_6_port, B(5) => 
                           Immediate_26_extended_5_port, B(4) => 
                           Immediate_26_extended_4_port, B(3) => 
                           Immediate_26_extended_3_port, B(2) => 
                           Immediate_26_extended_2_port, B(1) => 
                           Immediate_26_extended_1_port, B(0) => 
                           Immediate_26_extended_0_port, SEL => IMM_SEL, Y(31) 
                           => Immediate_selected_31_port, Y(30) => 
                           Immediate_selected_30_port, Y(29) => 
                           Immediate_selected_29_port, Y(28) => 
                           Immediate_selected_28_port, Y(27) => 
                           Immediate_selected_27_port, Y(26) => 
                           Immediate_selected_26_port, Y(25) => 
                           Immediate_selected_25_port, Y(24) => 
                           Immediate_selected_24_port, Y(23) => 
                           Immediate_selected_23_port, Y(22) => 
                           Immediate_selected_22_port, Y(21) => 
                           Immediate_selected_21_port, Y(20) => 
                           Immediate_selected_20_port, Y(19) => 
                           Immediate_selected_19_port, Y(18) => 
                           Immediate_selected_18_port, Y(17) => 
                           Immediate_selected_17_port, Y(16) => 
                           Immediate_selected_16_port, Y(15) => 
                           Immediate_selected_15_port, Y(14) => 
                           Immediate_selected_14_port, Y(13) => 
                           Immediate_selected_13_port, Y(12) => 
                           Immediate_selected_12_port, Y(11) => 
                           Immediate_selected_11_port, Y(10) => 
                           Immediate_selected_10_port, Y(9) => 
                           Immediate_selected_9_port, Y(8) => 
                           Immediate_selected_8_port, Y(7) => 
                           Immediate_selected_7_port, Y(6) => 
                           Immediate_selected_6_port, Y(5) => 
                           Immediate_selected_5_port, Y(4) => 
                           Immediate_selected_4_port, Y(3) => 
                           Immediate_selected_3_port, Y(2) => 
                           Immediate_selected_2_port, Y(1) => 
                           Immediate_selected_1_port, Y(0) => 
                           Immediate_selected_0_port);
   Immreg : reg_N32_11 port map( clk => Clk, rst => n452, d_in(31) => 
                           Immediate_selected_31_port, d_in(30) => 
                           Immediate_selected_30_port, d_in(29) => 
                           Immediate_selected_29_port, d_in(28) => 
                           Immediate_selected_28_port, d_in(27) => 
                           Immediate_selected_27_port, d_in(26) => 
                           Immediate_selected_26_port, d_in(25) => 
                           Immediate_selected_25_port, d_in(24) => 
                           Immediate_selected_24_port, d_in(23) => 
                           Immediate_selected_23_port, d_in(22) => 
                           Immediate_selected_22_port, d_in(21) => 
                           Immediate_selected_21_port, d_in(20) => 
                           Immediate_selected_20_port, d_in(19) => 
                           Immediate_selected_19_port, d_in(18) => 
                           Immediate_selected_18_port, d_in(17) => 
                           Immediate_selected_17_port, d_in(16) => 
                           Immediate_selected_16_port, d_in(15) => 
                           Immediate_selected_15_port, d_in(14) => 
                           Immediate_selected_14_port, d_in(13) => 
                           Immediate_selected_13_port, d_in(12) => 
                           Immediate_selected_12_port, d_in(11) => 
                           Immediate_selected_11_port, d_in(10) => 
                           Immediate_selected_10_port, d_in(9) => 
                           Immediate_selected_9_port, d_in(8) => 
                           Immediate_selected_8_port, d_in(7) => 
                           Immediate_selected_7_port, d_in(6) => 
                           Immediate_selected_6_port, d_in(5) => 
                           Immediate_selected_5_port, d_in(4) => 
                           Immediate_selected_4_port, d_in(3) => 
                           Immediate_selected_3_port, d_in(2) => 
                           Immediate_selected_2_port, d_in(1) => 
                           Immediate_selected_1_port, d_in(0) => 
                           Immediate_selected_0_port, d_out(31) => 
                           Immediate_clocked_31_port, d_out(30) => 
                           Immediate_clocked_30_port, d_out(29) => 
                           Immediate_clocked_29_port, d_out(28) => 
                           Immediate_clocked_28_port, d_out(27) => 
                           Immediate_clocked_27_port, d_out(26) => 
                           Immediate_clocked_26_port, d_out(25) => 
                           Immediate_clocked_25_port, d_out(24) => 
                           Immediate_clocked_24_port, d_out(23) => 
                           Immediate_clocked_23_port, d_out(22) => 
                           Immediate_clocked_22_port, d_out(21) => 
                           Immediate_clocked_21_port, d_out(20) => 
                           Immediate_clocked_20_port, d_out(19) => 
                           Immediate_clocked_19_port, d_out(18) => 
                           Immediate_clocked_18_port, d_out(17) => 
                           Immediate_clocked_17_port, d_out(16) => 
                           Immediate_clocked_16_port, d_out(15) => 
                           Immediate_clocked_15_port, d_out(14) => 
                           Immediate_clocked_14_port, d_out(13) => 
                           Immediate_clocked_13_port, d_out(12) => 
                           Immediate_clocked_12_port, d_out(11) => 
                           Immediate_clocked_11_port, d_out(10) => 
                           Immediate_clocked_10_port, d_out(9) => 
                           Immediate_clocked_9_port, d_out(8) => 
                           Immediate_clocked_8_port, d_out(7) => 
                           Immediate_clocked_7_port, d_out(6) => 
                           Immediate_clocked_6_port, d_out(5) => 
                           Immediate_clocked_5_port, d_out(4) => 
                           Immediate_clocked_4_port, d_out(3) => 
                           Immediate_clocked_3_port, d_out(2) => 
                           Immediate_clocked_2_port, d_out(1) => 
                           Immediate_clocked_1_port, d_out(0) => 
                           Immediate_clocked_0_port);
   MUX_A : MUX21_GENERIC_N32_4 port map( A(31) => NPC2_31_port, A(30) => 
                           NPC2_30_port, A(29) => NPC2_29_port, A(28) => 
                           NPC2_28_port, A(27) => NPC2_27_port, A(26) => 
                           NPC2_26_port, A(25) => NPC2_25_port, A(24) => 
                           NPC2_24_port, A(23) => NPC2_23_port, A(22) => 
                           NPC2_22_port, A(21) => NPC2_21_port, A(20) => 
                           NPC2_20_port, A(19) => NPC2_19_port, A(18) => 
                           NPC2_18_port, A(17) => NPC2_17_port, A(16) => 
                           NPC2_16_port, A(15) => NPC2_15_port, A(14) => 
                           NPC2_14_port, A(13) => NPC2_13_port, A(12) => 
                           NPC2_12_port, A(11) => NPC2_11_port, A(10) => 
                           NPC2_10_port, A(9) => NPC2_9_port, A(8) => 
                           NPC2_8_port, A(7) => NPC2_7_port, A(6) => 
                           NPC2_6_port, A(5) => NPC2_5_port, A(4) => 
                           NPC2_4_port, A(3) => NPC2_3_port, A(2) => 
                           NPC2_2_port, A(1) => NPC2_1_port, A(0) => 
                           NPC2_0_port, B(31) => A_reg_out_31_port, B(30) => 
                           A_reg_out_30_port, B(29) => A_reg_out_29_port, B(28)
                           => A_reg_out_28_port, B(27) => A_reg_out_27_port, 
                           B(26) => A_reg_out_26_port, B(25) => 
                           A_reg_out_25_port, B(24) => A_reg_out_24_port, B(23)
                           => A_reg_out_23_port, B(22) => A_reg_out_22_port, 
                           B(21) => A_reg_out_21_port, B(20) => 
                           A_reg_out_20_port, B(19) => A_reg_out_19_port, B(18)
                           => A_reg_out_18_port, B(17) => A_reg_out_17_port, 
                           B(16) => A_reg_out_16_port, B(15) => 
                           A_reg_out_15_port, B(14) => A_reg_out_14_port, B(13)
                           => A_reg_out_13_port, B(12) => A_reg_out_12_port, 
                           B(11) => A_reg_out_11_port, B(10) => 
                           A_reg_out_10_port, B(9) => A_reg_out_9_port, B(8) =>
                           A_reg_out_8_port, B(7) => A_reg_out_7_port, B(6) => 
                           A_reg_out_6_port, B(5) => A_reg_out_5_port, B(4) => 
                           A_reg_out_4_port, B(3) => A_reg_out_3_port, B(2) => 
                           A_reg_out_2_port, B(1) => A_reg_out_1_port, B(0) => 
                           A_reg_out_0_port, SEL => MUXA_SEL, Y(31) => 
                           ALU_operand_1_31_port, Y(30) => 
                           ALU_operand_1_30_port, Y(29) => 
                           ALU_operand_1_29_port, Y(28) => 
                           ALU_operand_1_28_port, Y(27) => 
                           ALU_operand_1_27_port, Y(26) => 
                           ALU_operand_1_26_port, Y(25) => 
                           ALU_operand_1_25_port, Y(24) => 
                           ALU_operand_1_24_port, Y(23) => 
                           ALU_operand_1_23_port, Y(22) => 
                           ALU_operand_1_22_port, Y(21) => 
                           ALU_operand_1_21_port, Y(20) => 
                           ALU_operand_1_20_port, Y(19) => 
                           ALU_operand_1_19_port, Y(18) => 
                           ALU_operand_1_18_port, Y(17) => 
                           ALU_operand_1_17_port, Y(16) => 
                           ALU_operand_1_16_port, Y(15) => 
                           ALU_operand_1_15_port, Y(14) => 
                           ALU_operand_1_14_port, Y(13) => 
                           ALU_operand_1_13_port, Y(12) => 
                           ALU_operand_1_12_port, Y(11) => 
                           ALU_operand_1_11_port, Y(10) => 
                           ALU_operand_1_10_port, Y(9) => ALU_operand_1_9_port,
                           Y(8) => ALU_operand_1_8_port, Y(7) => 
                           ALU_operand_1_7_port, Y(6) => ALU_operand_1_6_port, 
                           Y(5) => ALU_operand_1_5_port, Y(4) => 
                           ALU_operand_1_4_port, Y(3) => ALU_operand_1_3_port, 
                           Y(2) => ALU_operand_1_2_port, Y(1) => 
                           ALU_operand_1_1_port, Y(0) => ALU_operand_1_0_port);
   MUX_B : MUX21_GENERIC_N32_3 port map( A(31) => B_reg_out_31_port, A(30) => 
                           B_reg_out_30_port, A(29) => B_reg_out_29_port, A(28)
                           => B_reg_out_28_port, A(27) => B_reg_out_27_port, 
                           A(26) => B_reg_out_26_port, A(25) => 
                           B_reg_out_25_port, A(24) => B_reg_out_24_port, A(23)
                           => B_reg_out_23_port, A(22) => B_reg_out_22_port, 
                           A(21) => B_reg_out_21_port, A(20) => 
                           B_reg_out_20_port, A(19) => B_reg_out_19_port, A(18)
                           => B_reg_out_18_port, A(17) => B_reg_out_17_port, 
                           A(16) => B_reg_out_16_port, A(15) => 
                           B_reg_out_15_port, A(14) => B_reg_out_14_port, A(13)
                           => B_reg_out_13_port, A(12) => B_reg_out_12_port, 
                           A(11) => B_reg_out_11_port, A(10) => 
                           B_reg_out_10_port, A(9) => B_reg_out_9_port, A(8) =>
                           B_reg_out_8_port, A(7) => B_reg_out_7_port, A(6) => 
                           B_reg_out_6_port, A(5) => B_reg_out_5_port, A(4) => 
                           B_reg_out_4_port, A(3) => B_reg_out_3_port, A(2) => 
                           B_reg_out_2_port, A(1) => B_reg_out_1_port, A(0) => 
                           B_reg_out_0_port, B(31) => Immediate_clocked_31_port
                           , B(30) => Immediate_clocked_30_port, B(29) => 
                           Immediate_clocked_29_port, B(28) => 
                           Immediate_clocked_28_port, B(27) => 
                           Immediate_clocked_27_port, B(26) => 
                           Immediate_clocked_26_port, B(25) => 
                           Immediate_clocked_25_port, B(24) => 
                           Immediate_clocked_24_port, B(23) => 
                           Immediate_clocked_23_port, B(22) => 
                           Immediate_clocked_22_port, B(21) => 
                           Immediate_clocked_21_port, B(20) => 
                           Immediate_clocked_20_port, B(19) => 
                           Immediate_clocked_19_port, B(18) => 
                           Immediate_clocked_18_port, B(17) => 
                           Immediate_clocked_17_port, B(16) => 
                           Immediate_clocked_16_port, B(15) => 
                           Immediate_clocked_15_port, B(14) => 
                           Immediate_clocked_14_port, B(13) => 
                           Immediate_clocked_13_port, B(12) => 
                           Immediate_clocked_12_port, B(11) => 
                           Immediate_clocked_11_port, B(10) => 
                           Immediate_clocked_10_port, B(9) => 
                           Immediate_clocked_9_port, B(8) => 
                           Immediate_clocked_8_port, B(7) => 
                           Immediate_clocked_7_port, B(6) => 
                           Immediate_clocked_6_port, B(5) => 
                           Immediate_clocked_5_port, B(4) => 
                           Immediate_clocked_4_port, B(3) => 
                           Immediate_clocked_3_port, B(2) => 
                           Immediate_clocked_2_port, B(1) => 
                           Immediate_clocked_1_port, B(0) => 
                           Immediate_clocked_0_port, SEL => MUXB_SEL, Y(31) => 
                           ALU_operand_2_31_port, Y(30) => 
                           ALU_operand_2_30_port, Y(29) => 
                           ALU_operand_2_29_port, Y(28) => 
                           ALU_operand_2_28_port, Y(27) => 
                           ALU_operand_2_27_port, Y(26) => 
                           ALU_operand_2_26_port, Y(25) => 
                           ALU_operand_2_25_port, Y(24) => 
                           ALU_operand_2_24_port, Y(23) => 
                           ALU_operand_2_23_port, Y(22) => 
                           ALU_operand_2_22_port, Y(21) => 
                           ALU_operand_2_21_port, Y(20) => 
                           ALU_operand_2_20_port, Y(19) => 
                           ALU_operand_2_19_port, Y(18) => 
                           ALU_operand_2_18_port, Y(17) => 
                           ALU_operand_2_17_port, Y(16) => 
                           ALU_operand_2_16_port, Y(15) => 
                           ALU_operand_2_15_port, Y(14) => 
                           ALU_operand_2_14_port, Y(13) => 
                           ALU_operand_2_13_port, Y(12) => 
                           ALU_operand_2_12_port, Y(11) => 
                           ALU_operand_2_11_port, Y(10) => 
                           ALU_operand_2_10_port, Y(9) => ALU_operand_2_9_port,
                           Y(8) => ALU_operand_2_8_port, Y(7) => 
                           ALU_operand_2_7_port, Y(6) => ALU_operand_2_6_port, 
                           Y(5) => ALU_operand_2_5_port, Y(4) => 
                           ALU_operand_2_4_port, Y(3) => ALU_operand_2_3_port, 
                           Y(2) => ALU_operand_2_2_port, Y(1) => 
                           ALU_operand_2_1_port, Y(0) => ALU_operand_2_0_port);
   ALU_REG : reg_N32_10 port map( clk => Clk, rst => n451, d_in(31) => 
                           ALU_output_FWD_31_port, d_in(30) => 
                           ALU_output_FWD_30_port, d_in(29) => 
                           ALU_output_FWD_29_port, d_in(28) => 
                           ALU_output_FWD_28_port, d_in(27) => 
                           ALU_output_FWD_27_port, d_in(26) => 
                           ALU_output_FWD_26_port, d_in(25) => 
                           ALU_output_FWD_25_port, d_in(24) => 
                           ALU_output_FWD_24_port, d_in(23) => 
                           ALU_output_FWD_23_port, d_in(22) => 
                           ALU_output_FWD_22_port, d_in(21) => 
                           ALU_output_FWD_21_port, d_in(20) => 
                           ALU_output_FWD_20_port, d_in(19) => 
                           ALU_output_FWD_19_port, d_in(18) => 
                           ALU_output_FWD_18_port, d_in(17) => 
                           ALU_output_FWD_17_port, d_in(16) => 
                           ALU_output_FWD_16_port, d_in(15) => 
                           ALU_output_FWD_15_port, d_in(14) => 
                           ALU_output_FWD_14_port, d_in(13) => 
                           ALU_output_FWD_13_port, d_in(12) => 
                           ALU_output_FWD_12_port, d_in(11) => 
                           ALU_output_FWD_11_port, d_in(10) => 
                           ALU_output_FWD_10_port, d_in(9) => 
                           ALU_output_FWD_9_port, d_in(8) => 
                           ALU_output_FWD_8_port, d_in(7) => 
                           ALU_output_FWD_7_port, d_in(6) => 
                           ALU_output_FWD_6_port, d_in(5) => 
                           ALU_output_FWD_5_port, d_in(4) => 
                           ALU_output_FWD_4_port, d_in(3) => 
                           ALU_output_FWD_3_port, d_in(2) => 
                           ALU_output_FWD_2_port, d_in(1) => 
                           ALU_output_FWD_1_port, d_in(0) => 
                           ALU_output_FWD_0_port, d_out(31) => 
                           ALU_reg_out_31_port, d_out(30) => 
                           ALU_reg_out_30_port, d_out(29) => 
                           ALU_reg_out_29_port, d_out(28) => 
                           ALU_reg_out_28_port, d_out(27) => 
                           ALU_reg_out_27_port, d_out(26) => 
                           ALU_reg_out_26_port, d_out(25) => 
                           ALU_reg_out_25_port, d_out(24) => 
                           ALU_reg_out_24_port, d_out(23) => 
                           ALU_reg_out_23_port, d_out(22) => 
                           ALU_reg_out_22_port, d_out(21) => 
                           ALU_reg_out_21_port, d_out(20) => 
                           ALU_reg_out_20_port, d_out(19) => 
                           ALU_reg_out_19_port, d_out(18) => 
                           ALU_reg_out_18_port, d_out(17) => 
                           ALU_reg_out_17_port, d_out(16) => 
                           ALU_reg_out_16_port, d_out(15) => 
                           ALU_reg_out_15_port, d_out(14) => 
                           ALU_reg_out_14_port, d_out(13) => 
                           ALU_reg_out_13_port, d_out(12) => 
                           ALU_reg_out_12_port, d_out(11) => 
                           ALU_reg_out_11_port, d_out(10) => 
                           ALU_reg_out_10_port, d_out(9) => ALU_reg_out_9_port,
                           d_out(8) => ALU_reg_out_8_port, d_out(7) => 
                           ALU_reg_out_7_port, d_out(6) => ALU_reg_out_6_port, 
                           d_out(5) => ALU_reg_out_5_port, d_out(4) => 
                           ALU_reg_out_4_port, d_out(3) => ALU_reg_out_3_port, 
                           d_out(2) => ALU_reg_out_2_port, d_out(1) => 
                           ALU_reg_out_1_port, d_out(0) => ALU_reg_out_0_port);
   BREG : reg_N32_9 port map( clk => Clk, rst => n452, d_in(31) => 
                           B_reg_out_31_port, d_in(30) => B_reg_out_30_port, 
                           d_in(29) => B_reg_out_29_port, d_in(28) => 
                           B_reg_out_28_port, d_in(27) => B_reg_out_27_port, 
                           d_in(26) => B_reg_out_26_port, d_in(25) => 
                           B_reg_out_25_port, d_in(24) => B_reg_out_24_port, 
                           d_in(23) => B_reg_out_23_port, d_in(22) => 
                           B_reg_out_22_port, d_in(21) => B_reg_out_21_port, 
                           d_in(20) => B_reg_out_20_port, d_in(19) => 
                           B_reg_out_19_port, d_in(18) => B_reg_out_18_port, 
                           d_in(17) => B_reg_out_17_port, d_in(16) => 
                           B_reg_out_16_port, d_in(15) => B_reg_out_15_port, 
                           d_in(14) => B_reg_out_14_port, d_in(13) => 
                           B_reg_out_13_port, d_in(12) => B_reg_out_12_port, 
                           d_in(11) => B_reg_out_11_port, d_in(10) => 
                           B_reg_out_10_port, d_in(9) => B_reg_out_9_port, 
                           d_in(8) => B_reg_out_8_port, d_in(7) => 
                           B_reg_out_7_port, d_in(6) => B_reg_out_6_port, 
                           d_in(5) => B_reg_out_5_port, d_in(4) => 
                           B_reg_out_4_port, d_in(3) => B_reg_out_3_port, 
                           d_in(2) => B_reg_out_2_port, d_in(1) => 
                           B_reg_out_1_port, d_in(0) => B_reg_out_0_port, 
                           d_out(31) => DRAM_write_data_31_port, d_out(30) => 
                           DRAM_write_data_30_port, d_out(29) => 
                           DRAM_write_data_29_port, d_out(28) => 
                           DRAM_write_data_28_port, d_out(27) => 
                           DRAM_write_data_27_port, d_out(26) => 
                           DRAM_write_data_26_port, d_out(25) => 
                           DRAM_write_data_25_port, d_out(24) => 
                           DRAM_write_data_24_port, d_out(23) => 
                           DRAM_write_data_23_port, d_out(22) => 
                           DRAM_write_data_22_port, d_out(21) => 
                           DRAM_write_data_21_port, d_out(20) => 
                           DRAM_write_data_20_port, d_out(19) => 
                           DRAM_write_data_19_port, d_out(18) => 
                           DRAM_write_data_18_port, d_out(17) => 
                           DRAM_write_data_17_port, d_out(16) => 
                           DRAM_write_data_16_port, d_out(15) => 
                           DRAM_write_data_15_port, d_out(14) => 
                           DRAM_write_data_14_port, d_out(13) => 
                           DRAM_write_data_13_port, d_out(12) => 
                           DRAM_write_data_12_port, d_out(11) => 
                           DRAM_write_data_11_port, d_out(10) => 
                           DRAM_write_data_10_port, d_out(9) => 
                           DRAM_write_data_9_port, d_out(8) => 
                           DRAM_write_data_8_port, d_out(7) => 
                           DRAM_write_data_7_port, d_out(6) => 
                           DRAM_write_data_6_port, d_out(5) => 
                           DRAM_write_data_5_port, d_out(4) => 
                           DRAM_write_data_4_port, d_out(3) => 
                           DRAM_write_data_3_port, d_out(2) => 
                           DRAM_write_data_2_port, d_out(1) => 
                           DRAM_write_data_1_port, d_out(0) => 
                           DRAM_write_data_0_port);
   dataram : DRAM port map( clk => Clk, rst => n453, WR => DRAM_WR, 
                           sel_store(1) => SEL_STORE1, sel_store(0) => 
                           SEL_STORE0, sel_load(2) => SEL_LOAD2, sel_load(1) =>
                           SEL_LOAD1, sel_load(0) => SEL_LOAD0, addr(11) => 
                           ALU_reg_out_11_port, addr(10) => ALU_reg_out_10_port
                           , addr(9) => ALU_reg_out_9_port, addr(8) => 
                           ALU_reg_out_8_port, addr(7) => ALU_reg_out_7_port, 
                           addr(6) => ALU_reg_out_6_port, addr(5) => 
                           ALU_reg_out_5_port, addr(4) => ALU_reg_out_4_port, 
                           addr(3) => ALU_reg_out_3_port, addr(2) => 
                           ALU_reg_out_2_port, addr(1) => ALU_reg_out_1_port, 
                           addr(0) => ALU_reg_out_0_port, d_in(31) => 
                           DRAM_write_data_FWD_31_port, d_in(30) => 
                           DRAM_write_data_FWD_30_port, d_in(29) => 
                           DRAM_write_data_FWD_29_port, d_in(28) => 
                           DRAM_write_data_FWD_28_port, d_in(27) => 
                           DRAM_write_data_FWD_27_port, d_in(26) => 
                           DRAM_write_data_FWD_26_port, d_in(25) => 
                           DRAM_write_data_FWD_25_port, d_in(24) => 
                           DRAM_write_data_FWD_24_port, d_in(23) => 
                           DRAM_write_data_FWD_23_port, d_in(22) => 
                           DRAM_write_data_FWD_22_port, d_in(21) => 
                           DRAM_write_data_FWD_21_port, d_in(20) => 
                           DRAM_write_data_FWD_20_port, d_in(19) => 
                           DRAM_write_data_FWD_19_port, d_in(18) => 
                           DRAM_write_data_FWD_18_port, d_in(17) => 
                           DRAM_write_data_FWD_17_port, d_in(16) => 
                           DRAM_write_data_FWD_16_port, d_in(15) => 
                           DRAM_write_data_FWD_15_port, d_in(14) => 
                           DRAM_write_data_FWD_14_port, d_in(13) => 
                           DRAM_write_data_FWD_13_port, d_in(12) => 
                           DRAM_write_data_FWD_12_port, d_in(11) => 
                           DRAM_write_data_FWD_11_port, d_in(10) => 
                           DRAM_write_data_FWD_10_port, d_in(9) => 
                           DRAM_write_data_FWD_9_port, d_in(8) => 
                           DRAM_write_data_FWD_8_port, d_in(7) => 
                           DRAM_write_data_FWD_7_port, d_in(6) => 
                           DRAM_write_data_FWD_6_port, d_in(5) => 
                           DRAM_write_data_FWD_5_port, d_in(4) => 
                           DRAM_write_data_FWD_4_port, d_in(3) => 
                           DRAM_write_data_FWD_3_port, d_in(2) => 
                           DRAM_write_data_FWD_2_port, d_in(1) => 
                           DRAM_write_data_FWD_1_port, d_in(0) => 
                           DRAM_write_data_FWD_0_port, d_out(31) => 
                           DRAM_read_data_31_port, d_out(30) => 
                           DRAM_read_data_30_port, d_out(29) => 
                           DRAM_read_data_29_port, d_out(28) => 
                           DRAM_read_data_28_port, d_out(27) => 
                           DRAM_read_data_27_port, d_out(26) => 
                           DRAM_read_data_26_port, d_out(25) => 
                           DRAM_read_data_25_port, d_out(24) => 
                           DRAM_read_data_24_port, d_out(23) => 
                           DRAM_read_data_23_port, d_out(22) => 
                           DRAM_read_data_22_port, d_out(21) => 
                           DRAM_read_data_21_port, d_out(20) => 
                           DRAM_read_data_20_port, d_out(19) => 
                           DRAM_read_data_19_port, d_out(18) => 
                           DRAM_read_data_18_port, d_out(17) => 
                           DRAM_read_data_17_port, d_out(16) => 
                           DRAM_read_data_16_port, d_out(15) => 
                           DRAM_read_data_15_port, d_out(14) => 
                           DRAM_read_data_14_port, d_out(13) => 
                           DRAM_read_data_13_port, d_out(12) => 
                           DRAM_read_data_12_port, d_out(11) => 
                           DRAM_read_data_11_port, d_out(10) => 
                           DRAM_read_data_10_port, d_out(9) => 
                           DRAM_read_data_9_port, d_out(8) => 
                           DRAM_read_data_8_port, d_out(7) => 
                           DRAM_read_data_7_port, d_out(6) => 
                           DRAM_read_data_6_port, d_out(5) => 
                           DRAM_read_data_5_port, d_out(4) => 
                           DRAM_read_data_4_port, d_out(3) => 
                           DRAM_read_data_3_port, d_out(2) => 
                           DRAM_read_data_2_port, d_out(1) => 
                           DRAM_read_data_1_port, d_out(0) => 
                           DRAM_read_data_0_port);
   LMD : reg_N32_8 port map( clk => Clk, rst => n452, d_in(31) => 
                           DRAM_read_data_31_port, d_in(30) => 
                           DRAM_read_data_30_port, d_in(29) => 
                           DRAM_read_data_29_port, d_in(28) => 
                           DRAM_read_data_28_port, d_in(27) => 
                           DRAM_read_data_27_port, d_in(26) => 
                           DRAM_read_data_26_port, d_in(25) => 
                           DRAM_read_data_25_port, d_in(24) => 
                           DRAM_read_data_24_port, d_in(23) => 
                           DRAM_read_data_23_port, d_in(22) => 
                           DRAM_read_data_22_port, d_in(21) => 
                           DRAM_read_data_21_port, d_in(20) => 
                           DRAM_read_data_20_port, d_in(19) => 
                           DRAM_read_data_19_port, d_in(18) => 
                           DRAM_read_data_18_port, d_in(17) => 
                           DRAM_read_data_17_port, d_in(16) => 
                           DRAM_read_data_16_port, d_in(15) => 
                           DRAM_read_data_15_port, d_in(14) => 
                           DRAM_read_data_14_port, d_in(13) => 
                           DRAM_read_data_13_port, d_in(12) => 
                           DRAM_read_data_12_port, d_in(11) => 
                           DRAM_read_data_11_port, d_in(10) => 
                           DRAM_read_data_10_port, d_in(9) => 
                           DRAM_read_data_9_port, d_in(8) => 
                           DRAM_read_data_8_port, d_in(7) => 
                           DRAM_read_data_7_port, d_in(6) => 
                           DRAM_read_data_6_port, d_in(5) => 
                           DRAM_read_data_5_port, d_in(4) => 
                           DRAM_read_data_4_port, d_in(3) => 
                           DRAM_read_data_3_port, d_in(2) => 
                           DRAM_read_data_2_port, d_in(1) => 
                           DRAM_read_data_1_port, d_in(0) => 
                           DRAM_read_data_0_port, d_out(31) => 
                           LMD_reg_out_31_port, d_out(30) => 
                           LMD_reg_out_30_port, d_out(29) => 
                           LMD_reg_out_29_port, d_out(28) => 
                           LMD_reg_out_28_port, d_out(27) => 
                           LMD_reg_out_27_port, d_out(26) => 
                           LMD_reg_out_26_port, d_out(25) => 
                           LMD_reg_out_25_port, d_out(24) => 
                           LMD_reg_out_24_port, d_out(23) => 
                           LMD_reg_out_23_port, d_out(22) => 
                           LMD_reg_out_22_port, d_out(21) => 
                           LMD_reg_out_21_port, d_out(20) => 
                           LMD_reg_out_20_port, d_out(19) => 
                           LMD_reg_out_19_port, d_out(18) => 
                           LMD_reg_out_18_port, d_out(17) => 
                           LMD_reg_out_17_port, d_out(16) => 
                           LMD_reg_out_16_port, d_out(15) => 
                           LMD_reg_out_15_port, d_out(14) => 
                           LMD_reg_out_14_port, d_out(13) => 
                           LMD_reg_out_13_port, d_out(12) => 
                           LMD_reg_out_12_port, d_out(11) => 
                           LMD_reg_out_11_port, d_out(10) => 
                           LMD_reg_out_10_port, d_out(9) => LMD_reg_out_9_port,
                           d_out(8) => LMD_reg_out_8_port, d_out(7) => 
                           LMD_reg_out_7_port, d_out(6) => LMD_reg_out_6_port, 
                           d_out(5) => LMD_reg_out_5_port, d_out(4) => 
                           LMD_reg_out_4_port, d_out(3) => LMD_reg_out_3_port, 
                           d_out(2) => LMD_reg_out_2_port, d_out(1) => 
                           LMD_reg_out_1_port, d_out(0) => LMD_reg_out_0_port);
   LMD1 : reg_N32_7 port map( clk => Clk, rst => n452, d_in(31) => 
                           LMD_reg_out_31_port, d_in(30) => LMD_reg_out_30_port
                           , d_in(29) => LMD_reg_out_29_port, d_in(28) => 
                           LMD_reg_out_28_port, d_in(27) => LMD_reg_out_27_port
                           , d_in(26) => LMD_reg_out_26_port, d_in(25) => 
                           LMD_reg_out_25_port, d_in(24) => LMD_reg_out_24_port
                           , d_in(23) => LMD_reg_out_23_port, d_in(22) => 
                           LMD_reg_out_22_port, d_in(21) => LMD_reg_out_21_port
                           , d_in(20) => LMD_reg_out_20_port, d_in(19) => 
                           LMD_reg_out_19_port, d_in(18) => LMD_reg_out_18_port
                           , d_in(17) => LMD_reg_out_17_port, d_in(16) => 
                           LMD_reg_out_16_port, d_in(15) => LMD_reg_out_15_port
                           , d_in(14) => LMD_reg_out_14_port, d_in(13) => 
                           LMD_reg_out_13_port, d_in(12) => LMD_reg_out_12_port
                           , d_in(11) => LMD_reg_out_11_port, d_in(10) => 
                           LMD_reg_out_10_port, d_in(9) => LMD_reg_out_9_port, 
                           d_in(8) => LMD_reg_out_8_port, d_in(7) => 
                           LMD_reg_out_7_port, d_in(6) => LMD_reg_out_6_port, 
                           d_in(5) => LMD_reg_out_5_port, d_in(4) => 
                           LMD_reg_out_4_port, d_in(3) => LMD_reg_out_3_port, 
                           d_in(2) => LMD_reg_out_2_port, d_in(1) => 
                           LMD_reg_out_1_port, d_in(0) => LMD_reg_out_0_port, 
                           d_out(31) => LMD_reg_out1_31_port, d_out(30) => 
                           LMD_reg_out1_30_port, d_out(29) => 
                           LMD_reg_out1_29_port, d_out(28) => 
                           LMD_reg_out1_28_port, d_out(27) => 
                           LMD_reg_out1_27_port, d_out(26) => 
                           LMD_reg_out1_26_port, d_out(25) => 
                           LMD_reg_out1_25_port, d_out(24) => 
                           LMD_reg_out1_24_port, d_out(23) => 
                           LMD_reg_out1_23_port, d_out(22) => 
                           LMD_reg_out1_22_port, d_out(21) => 
                           LMD_reg_out1_21_port, d_out(20) => 
                           LMD_reg_out1_20_port, d_out(19) => 
                           LMD_reg_out1_19_port, d_out(18) => 
                           LMD_reg_out1_18_port, d_out(17) => 
                           LMD_reg_out1_17_port, d_out(16) => 
                           LMD_reg_out1_16_port, d_out(15) => 
                           LMD_reg_out1_15_port, d_out(14) => 
                           LMD_reg_out1_14_port, d_out(13) => 
                           LMD_reg_out1_13_port, d_out(12) => 
                           LMD_reg_out1_12_port, d_out(11) => 
                           LMD_reg_out1_11_port, d_out(10) => 
                           LMD_reg_out1_10_port, d_out(9) => 
                           LMD_reg_out1_9_port, d_out(8) => LMD_reg_out1_8_port
                           , d_out(7) => LMD_reg_out1_7_port, d_out(6) => 
                           LMD_reg_out1_6_port, d_out(5) => LMD_reg_out1_5_port
                           , d_out(4) => LMD_reg_out1_4_port, d_out(3) => 
                           LMD_reg_out1_3_port, d_out(2) => LMD_reg_out1_2_port
                           , d_out(1) => LMD_reg_out1_1_port, d_out(0) => 
                           LMD_reg_out1_0_port);
   ALUWB : reg_N32_6 port map( clk => Clk, rst => n451, d_in(31) => 
                           ALU_reg_out_31_port, d_in(30) => ALU_reg_out_30_port
                           , d_in(29) => ALU_reg_out_29_port, d_in(28) => 
                           ALU_reg_out_28_port, d_in(27) => ALU_reg_out_27_port
                           , d_in(26) => ALU_reg_out_26_port, d_in(25) => 
                           ALU_reg_out_25_port, d_in(24) => ALU_reg_out_24_port
                           , d_in(23) => ALU_reg_out_23_port, d_in(22) => 
                           ALU_reg_out_22_port, d_in(21) => ALU_reg_out_21_port
                           , d_in(20) => ALU_reg_out_20_port, d_in(19) => 
                           ALU_reg_out_19_port, d_in(18) => ALU_reg_out_18_port
                           , d_in(17) => ALU_reg_out_17_port, d_in(16) => 
                           ALU_reg_out_16_port, d_in(15) => ALU_reg_out_15_port
                           , d_in(14) => ALU_reg_out_14_port, d_in(13) => 
                           ALU_reg_out_13_port, d_in(12) => ALU_reg_out_12_port
                           , d_in(11) => ALU_reg_out_11_port, d_in(10) => 
                           ALU_reg_out_10_port, d_in(9) => ALU_reg_out_9_port, 
                           d_in(8) => ALU_reg_out_8_port, d_in(7) => 
                           ALU_reg_out_7_port, d_in(6) => ALU_reg_out_6_port, 
                           d_in(5) => ALU_reg_out_5_port, d_in(4) => 
                           ALU_reg_out_4_port, d_in(3) => ALU_reg_out_3_port, 
                           d_in(2) => ALU_reg_out_2_port, d_in(1) => 
                           ALU_reg_out_1_port, d_in(0) => ALU_reg_out_0_port, 
                           d_out(31) => ALU_WB_out_31_port, d_out(30) => 
                           ALU_WB_out_30_port, d_out(29) => ALU_WB_out_29_port,
                           d_out(28) => ALU_WB_out_28_port, d_out(27) => 
                           ALU_WB_out_27_port, d_out(26) => ALU_WB_out_26_port,
                           d_out(25) => ALU_WB_out_25_port, d_out(24) => 
                           ALU_WB_out_24_port, d_out(23) => ALU_WB_out_23_port,
                           d_out(22) => ALU_WB_out_22_port, d_out(21) => 
                           ALU_WB_out_21_port, d_out(20) => ALU_WB_out_20_port,
                           d_out(19) => ALU_WB_out_19_port, d_out(18) => 
                           ALU_WB_out_18_port, d_out(17) => ALU_WB_out_17_port,
                           d_out(16) => ALU_WB_out_16_port, d_out(15) => 
                           ALU_WB_out_15_port, d_out(14) => ALU_WB_out_14_port,
                           d_out(13) => ALU_WB_out_13_port, d_out(12) => 
                           ALU_WB_out_12_port, d_out(11) => ALU_WB_out_11_port,
                           d_out(10) => ALU_WB_out_10_port, d_out(9) => 
                           ALU_WB_out_9_port, d_out(8) => ALU_WB_out_8_port, 
                           d_out(7) => ALU_WB_out_7_port, d_out(6) => 
                           ALU_WB_out_6_port, d_out(5) => ALU_WB_out_5_port, 
                           d_out(4) => ALU_WB_out_4_port, d_out(3) => 
                           ALU_WB_out_3_port, d_out(2) => ALU_WB_out_2_port, 
                           d_out(1) => ALU_WB_out_1_port, d_out(0) => 
                           ALU_WB_out_0_port);
   ALUWB1 : reg_N32_5 port map( clk => Clk, rst => n451, d_in(31) => 
                           ALU_WB_out_31_port, d_in(30) => ALU_WB_out_30_port, 
                           d_in(29) => ALU_WB_out_29_port, d_in(28) => 
                           ALU_WB_out_28_port, d_in(27) => ALU_WB_out_27_port, 
                           d_in(26) => ALU_WB_out_26_port, d_in(25) => 
                           ALU_WB_out_25_port, d_in(24) => ALU_WB_out_24_port, 
                           d_in(23) => ALU_WB_out_23_port, d_in(22) => 
                           ALU_WB_out_22_port, d_in(21) => ALU_WB_out_21_port, 
                           d_in(20) => ALU_WB_out_20_port, d_in(19) => 
                           ALU_WB_out_19_port, d_in(18) => ALU_WB_out_18_port, 
                           d_in(17) => ALU_WB_out_17_port, d_in(16) => 
                           ALU_WB_out_16_port, d_in(15) => ALU_WB_out_15_port, 
                           d_in(14) => ALU_WB_out_14_port, d_in(13) => 
                           ALU_WB_out_13_port, d_in(12) => ALU_WB_out_12_port, 
                           d_in(11) => ALU_WB_out_11_port, d_in(10) => 
                           ALU_WB_out_10_port, d_in(9) => ALU_WB_out_9_port, 
                           d_in(8) => ALU_WB_out_8_port, d_in(7) => 
                           ALU_WB_out_7_port, d_in(6) => ALU_WB_out_6_port, 
                           d_in(5) => ALU_WB_out_5_port, d_in(4) => 
                           ALU_WB_out_4_port, d_in(3) => ALU_WB_out_3_port, 
                           d_in(2) => ALU_WB_out_2_port, d_in(1) => 
                           ALU_WB_out_1_port, d_in(0) => ALU_WB_out_0_port, 
                           d_out(31) => ALU_WB_out1_31_port, d_out(30) => 
                           ALU_WB_out1_30_port, d_out(29) => 
                           ALU_WB_out1_29_port, d_out(28) => 
                           ALU_WB_out1_28_port, d_out(27) => 
                           ALU_WB_out1_27_port, d_out(26) => 
                           ALU_WB_out1_26_port, d_out(25) => 
                           ALU_WB_out1_25_port, d_out(24) => 
                           ALU_WB_out1_24_port, d_out(23) => 
                           ALU_WB_out1_23_port, d_out(22) => 
                           ALU_WB_out1_22_port, d_out(21) => 
                           ALU_WB_out1_21_port, d_out(20) => 
                           ALU_WB_out1_20_port, d_out(19) => 
                           ALU_WB_out1_19_port, d_out(18) => 
                           ALU_WB_out1_18_port, d_out(17) => 
                           ALU_WB_out1_17_port, d_out(16) => 
                           ALU_WB_out1_16_port, d_out(15) => 
                           ALU_WB_out1_15_port, d_out(14) => 
                           ALU_WB_out1_14_port, d_out(13) => 
                           ALU_WB_out1_13_port, d_out(12) => 
                           ALU_WB_out1_12_port, d_out(11) => 
                           ALU_WB_out1_11_port, d_out(10) => 
                           ALU_WB_out1_10_port, d_out(9) => ALU_WB_out1_9_port,
                           d_out(8) => ALU_WB_out1_8_port, d_out(7) => 
                           ALU_WB_out1_7_port, d_out(6) => ALU_WB_out1_6_port, 
                           d_out(5) => ALU_WB_out1_5_port, d_out(4) => 
                           ALU_WB_out1_4_port, d_out(3) => ALU_WB_out1_3_port, 
                           d_out(2) => ALU_WB_out1_2_port, d_out(1) => 
                           ALU_WB_out1_1_port, d_out(0) => ALU_WB_out1_0_port);
   mux_WB : MUX21_GENERIC_N32_2 port map( A(31) => LMD_reg_out_31_port, A(30) 
                           => LMD_reg_out_30_port, A(29) => LMD_reg_out_29_port
                           , A(28) => LMD_reg_out_28_port, A(27) => 
                           LMD_reg_out_27_port, A(26) => LMD_reg_out_26_port, 
                           A(25) => LMD_reg_out_25_port, A(24) => 
                           LMD_reg_out_24_port, A(23) => LMD_reg_out_23_port, 
                           A(22) => LMD_reg_out_22_port, A(21) => 
                           LMD_reg_out_21_port, A(20) => LMD_reg_out_20_port, 
                           A(19) => LMD_reg_out_19_port, A(18) => 
                           LMD_reg_out_18_port, A(17) => LMD_reg_out_17_port, 
                           A(16) => LMD_reg_out_16_port, A(15) => 
                           LMD_reg_out_15_port, A(14) => LMD_reg_out_14_port, 
                           A(13) => LMD_reg_out_13_port, A(12) => 
                           LMD_reg_out_12_port, A(11) => LMD_reg_out_11_port, 
                           A(10) => LMD_reg_out_10_port, A(9) => 
                           LMD_reg_out_9_port, A(8) => LMD_reg_out_8_port, A(7)
                           => LMD_reg_out_7_port, A(6) => LMD_reg_out_6_port, 
                           A(5) => LMD_reg_out_5_port, A(4) => 
                           LMD_reg_out_4_port, A(3) => LMD_reg_out_3_port, A(2)
                           => LMD_reg_out_2_port, A(1) => LMD_reg_out_1_port, 
                           A(0) => LMD_reg_out_0_port, B(31) => 
                           ALU_WB_out_31_port, B(30) => ALU_WB_out_30_port, 
                           B(29) => ALU_WB_out_29_port, B(28) => 
                           ALU_WB_out_28_port, B(27) => ALU_WB_out_27_port, 
                           B(26) => ALU_WB_out_26_port, B(25) => 
                           ALU_WB_out_25_port, B(24) => ALU_WB_out_24_port, 
                           B(23) => ALU_WB_out_23_port, B(22) => 
                           ALU_WB_out_22_port, B(21) => ALU_WB_out_21_port, 
                           B(20) => ALU_WB_out_20_port, B(19) => 
                           ALU_WB_out_19_port, B(18) => ALU_WB_out_18_port, 
                           B(17) => ALU_WB_out_17_port, B(16) => 
                           ALU_WB_out_16_port, B(15) => ALU_WB_out_15_port, 
                           B(14) => ALU_WB_out_14_port, B(13) => 
                           ALU_WB_out_13_port, B(12) => ALU_WB_out_12_port, 
                           B(11) => ALU_WB_out_11_port, B(10) => 
                           ALU_WB_out_10_port, B(9) => ALU_WB_out_9_port, B(8) 
                           => ALU_WB_out_8_port, B(7) => ALU_WB_out_7_port, 
                           B(6) => ALU_WB_out_6_port, B(5) => ALU_WB_out_5_port
                           , B(4) => ALU_WB_out_4_port, B(3) => 
                           ALU_WB_out_3_port, B(2) => ALU_WB_out_2_port, B(1) 
                           => ALU_WB_out_1_port, B(0) => ALU_WB_out_0_port, SEL
                           => WB_MUX_SEL, Y(31) => WB_mux_out_31_port, Y(30) =>
                           WB_mux_out_30_port, Y(29) => WB_mux_out_29_port, 
                           Y(28) => WB_mux_out_28_port, Y(27) => 
                           WB_mux_out_27_port, Y(26) => WB_mux_out_26_port, 
                           Y(25) => WB_mux_out_25_port, Y(24) => 
                           WB_mux_out_24_port, Y(23) => WB_mux_out_23_port, 
                           Y(22) => WB_mux_out_22_port, Y(21) => 
                           WB_mux_out_21_port, Y(20) => WB_mux_out_20_port, 
                           Y(19) => WB_mux_out_19_port, Y(18) => 
                           WB_mux_out_18_port, Y(17) => WB_mux_out_17_port, 
                           Y(16) => WB_mux_out_16_port, Y(15) => 
                           WB_mux_out_15_port, Y(14) => WB_mux_out_14_port, 
                           Y(13) => WB_mux_out_13_port, Y(12) => 
                           WB_mux_out_12_port, Y(11) => WB_mux_out_11_port, 
                           Y(10) => WB_mux_out_10_port, Y(9) => 
                           WB_mux_out_9_port, Y(8) => WB_mux_out_8_port, Y(7) 
                           => WB_mux_out_7_port, Y(6) => WB_mux_out_6_port, 
                           Y(5) => WB_mux_out_5_port, Y(4) => WB_mux_out_4_port
                           , Y(3) => WB_mux_out_3_port, Y(2) => 
                           WB_mux_out_2_port, Y(1) => WB_mux_out_1_port, Y(0) 
                           => WB_mux_out_0_port);
   RFin_mux : MUX21_GENERIC_N32_1 port map( A(31) => NPC4_31_port, A(30) => 
                           NPC4_30_port, A(29) => NPC4_29_port, A(28) => 
                           NPC4_28_port, A(27) => NPC4_27_port, A(26) => 
                           NPC4_26_port, A(25) => NPC4_25_port, A(24) => 
                           NPC4_24_port, A(23) => NPC4_23_port, A(22) => 
                           NPC4_22_port, A(21) => NPC4_21_port, A(20) => 
                           NPC4_20_port, A(19) => NPC4_19_port, A(18) => 
                           NPC4_18_port, A(17) => NPC4_17_port, A(16) => 
                           NPC4_16_port, A(15) => NPC4_15_port, A(14) => 
                           NPC4_14_port, A(13) => NPC4_13_port, A(12) => 
                           NPC4_12_port, A(11) => NPC4_11_port, A(10) => 
                           NPC4_10_port, A(9) => NPC4_9_port, A(8) => 
                           NPC4_8_port, A(7) => NPC4_7_port, A(6) => 
                           NPC4_6_port, A(5) => NPC4_5_port, A(4) => 
                           NPC4_4_port, A(3) => NPC4_3_port, A(2) => 
                           NPC4_2_port, A(1) => NPC4_1_port, A(0) => 
                           NPC4_0_port, B(31) => WB_mux_out_31_port, B(30) => 
                           WB_mux_out_30_port, B(29) => WB_mux_out_29_port, 
                           B(28) => WB_mux_out_28_port, B(27) => 
                           WB_mux_out_27_port, B(26) => WB_mux_out_26_port, 
                           B(25) => WB_mux_out_25_port, B(24) => 
                           WB_mux_out_24_port, B(23) => WB_mux_out_23_port, 
                           B(22) => WB_mux_out_22_port, B(21) => 
                           WB_mux_out_21_port, B(20) => WB_mux_out_20_port, 
                           B(19) => WB_mux_out_19_port, B(18) => 
                           WB_mux_out_18_port, B(17) => WB_mux_out_17_port, 
                           B(16) => WB_mux_out_16_port, B(15) => 
                           WB_mux_out_15_port, B(14) => WB_mux_out_14_port, 
                           B(13) => WB_mux_out_13_port, B(12) => 
                           WB_mux_out_12_port, B(11) => WB_mux_out_11_port, 
                           B(10) => WB_mux_out_10_port, B(9) => 
                           WB_mux_out_9_port, B(8) => WB_mux_out_8_port, B(7) 
                           => WB_mux_out_7_port, B(6) => WB_mux_out_6_port, 
                           B(5) => WB_mux_out_5_port, B(4) => WB_mux_out_4_port
                           , B(3) => WB_mux_out_3_port, B(2) => 
                           WB_mux_out_2_port, B(1) => WB_mux_out_1_port, B(0) 
                           => WB_mux_out_0_port, SEL => JAL_op4, Y(31) => 
                           RF_write_data_31_port, Y(30) => 
                           RF_write_data_30_port, Y(29) => 
                           RF_write_data_29_port, Y(28) => 
                           RF_write_data_28_port, Y(27) => 
                           RF_write_data_27_port, Y(26) => 
                           RF_write_data_26_port, Y(25) => 
                           RF_write_data_25_port, Y(24) => 
                           RF_write_data_24_port, Y(23) => 
                           RF_write_data_23_port, Y(22) => 
                           RF_write_data_22_port, Y(21) => 
                           RF_write_data_21_port, Y(20) => 
                           RF_write_data_20_port, Y(19) => 
                           RF_write_data_19_port, Y(18) => 
                           RF_write_data_18_port, Y(17) => 
                           RF_write_data_17_port, Y(16) => 
                           RF_write_data_16_port, Y(15) => 
                           RF_write_data_15_port, Y(14) => 
                           RF_write_data_14_port, Y(13) => 
                           RF_write_data_13_port, Y(12) => 
                           RF_write_data_12_port, Y(11) => 
                           RF_write_data_11_port, Y(10) => 
                           RF_write_data_10_port, Y(9) => RF_write_data_9_port,
                           Y(8) => RF_write_data_8_port, Y(7) => 
                           RF_write_data_7_port, Y(6) => RF_write_data_6_port, 
                           Y(5) => RF_write_data_5_port, Y(4) => 
                           RF_write_data_4_port, Y(3) => RF_write_data_3_port, 
                           Y(2) => RF_write_data_2_port, Y(1) => 
                           RF_write_data_1_port, Y(0) => RF_write_data_0_port);
   PC : reg_en_N32 port map( clk => Clk, rst => n451, en => PC_enable_fixed, 
                           d_in(31) => PC_reg_in_31_port, d_in(30) => 
                           PC_reg_in_30_port, d_in(29) => PC_reg_in_29_port, 
                           d_in(28) => PC_reg_in_28_port, d_in(27) => 
                           PC_reg_in_27_port, d_in(26) => PC_reg_in_26_port, 
                           d_in(25) => PC_reg_in_25_port, d_in(24) => 
                           PC_reg_in_24_port, d_in(23) => PC_reg_in_23_port, 
                           d_in(22) => PC_reg_in_22_port, d_in(21) => 
                           PC_reg_in_21_port, d_in(20) => PC_reg_in_20_port, 
                           d_in(19) => PC_reg_in_19_port, d_in(18) => 
                           PC_reg_in_18_port, d_in(17) => PC_reg_in_17_port, 
                           d_in(16) => PC_reg_in_16_port, d_in(15) => 
                           PC_reg_in_15_port, d_in(14) => PC_reg_in_14_port, 
                           d_in(13) => PC_reg_in_13_port, d_in(12) => 
                           PC_reg_in_12_port, d_in(11) => PC_reg_in_11_port, 
                           d_in(10) => PC_reg_in_10_port, d_in(9) => 
                           PC_reg_in_9_port, d_in(8) => PC_reg_in_8_port, 
                           d_in(7) => PC_reg_in_7_port, d_in(6) => 
                           PC_reg_in_6_port, d_in(5) => PC_reg_in_5_port, 
                           d_in(4) => PC_reg_in_4_port, d_in(3) => 
                           PC_reg_in_3_port, d_in(2) => PC_reg_in_2_port, 
                           d_in(1) => PC_reg_in_1_port, d_in(0) => 
                           PC_reg_in_0_port, d_out(31) => PC_out_31, d_out(30) 
                           => PC_out_28_port, d_out(29) => PC_out_27_port, 
                           d_out(28) => PC_out_26_port, d_out(27) => 
                           PC_out_25_port, d_out(26) => PC_out_24_port, 
                           d_out(25) => PC_out_23_port, d_out(24) => 
                           PC_out_22_port, d_out(23) => PC_out_21_port, 
                           d_out(22) => PC_out_20_port, d_out(21) => 
                           PC_out_19_port, d_out(20) => PC_out_18_port, 
                           d_out(19) => PC_out_17_port, d_out(18) => 
                           PC_out_16_port, d_out(17) => PC_out_15_port, 
                           d_out(16) => PC_out_14_port, d_out(15) => 
                           PC_out_13_port, d_out(14) => PC_out_12_port, 
                           d_out(13) => PC_out_11_port, d_out(12) => 
                           PC_out_10_port, d_out(11) => PC_out_9_port, 
                           d_out(10) => PC_out_8_port, d_out(9) => 
                           PC_out_7_port, d_out(8) => PC_out_6_port, d_out(7) 
                           => PC_out_5_port, d_out(6) => PC_out_4_port, 
                           d_out(5) => PC_out_3_port, d_out(4) => PC_out_2_port
                           , d_out(3) => PC_out_1_port, d_out(2) => 
                           PC_out_0_port, d_out(1) => PC_reg_out_1_port, 
                           d_out(0) => PC_reg_out_0_port);
   PCi : PC_incr port map( PC(31) => PC_out_31, PC(30) => PC_out_28_port, 
                           PC(29) => PC_out_27_port, PC(28) => PC_out_26_port, 
                           PC(27) => PC_out_25_port, PC(26) => PC_out_24_port, 
                           PC(25) => PC_out_23_port, PC(24) => PC_out_22_port, 
                           PC(23) => PC_out_21_port, PC(22) => PC_out_20_port, 
                           PC(21) => PC_out_19_port, PC(20) => PC_out_18_port, 
                           PC(19) => PC_out_17_port, PC(18) => PC_out_16_port, 
                           PC(17) => PC_out_15_port, PC(16) => PC_out_14_port, 
                           PC(15) => PC_out_13_port, PC(14) => PC_out_12_port, 
                           PC(13) => PC_out_11_port, PC(12) => PC_out_10_port, 
                           PC(11) => PC_out_9_port, PC(10) => PC_out_8_port, 
                           PC(9) => PC_out_7_port, PC(8) => PC_out_6_port, 
                           PC(7) => PC_out_5_port, PC(6) => PC_out_4_port, 
                           PC(5) => PC_out_3_port, PC(4) => PC_out_2_port, 
                           PC(3) => PC_out_1_port, PC(2) => PC_out_0_port, 
                           PC(1) => PC_reg_out_1_port, PC(0) => 
                           PC_reg_out_0_port, NPC(31) => NPC_31_port, NPC(30) 
                           => NPC_30_port, NPC(29) => NPC_29_port, NPC(28) => 
                           NPC_28_port, NPC(27) => NPC_27_port, NPC(26) => 
                           NPC_26_port, NPC(25) => NPC_25_port, NPC(24) => 
                           NPC_24_port, NPC(23) => NPC_23_port, NPC(22) => 
                           NPC_22_port, NPC(21) => NPC_21_port, NPC(20) => 
                           NPC_20_port, NPC(19) => NPC_19_port, NPC(18) => 
                           NPC_18_port, NPC(17) => NPC_17_port, NPC(16) => 
                           NPC_16_port, NPC(15) => NPC_15_port, NPC(14) => 
                           NPC_14_port, NPC(13) => NPC_13_port, NPC(12) => 
                           NPC_12_port, NPC(11) => NPC_11_port, NPC(10) => 
                           NPC_10_port, NPC(9) => NPC_9_port, NPC(8) => 
                           NPC_8_port, NPC(7) => NPC_7_port, NPC(6) => 
                           NPC_6_port, NPC(5) => NPC_5_port, NPC(4) => 
                           NPC_4_port, NPC(3) => NPC_3_port, NPC(2) => 
                           NPC_2_port, NPC(1) => NPC_1_port, NPC(0) => 
                           NPC_0_port);
   NPCreg1 : reg_N32_4 port map( clk => Clk, rst => n451, d_in(31) => 
                           NPC_31_port, d_in(30) => NPC_30_port, d_in(29) => 
                           NPC_29_port, d_in(28) => NPC_28_port, d_in(27) => 
                           NPC_27_port, d_in(26) => NPC_26_port, d_in(25) => 
                           NPC_25_port, d_in(24) => NPC_24_port, d_in(23) => 
                           NPC_23_port, d_in(22) => NPC_22_port, d_in(21) => 
                           NPC_21_port, d_in(20) => NPC_20_port, d_in(19) => 
                           NPC_19_port, d_in(18) => NPC_18_port, d_in(17) => 
                           NPC_17_port, d_in(16) => NPC_16_port, d_in(15) => 
                           NPC_15_port, d_in(14) => NPC_14_port, d_in(13) => 
                           NPC_13_port, d_in(12) => NPC_12_port, d_in(11) => 
                           NPC_11_port, d_in(10) => NPC_10_port, d_in(9) => 
                           NPC_9_port, d_in(8) => NPC_8_port, d_in(7) => 
                           NPC_7_port, d_in(6) => NPC_6_port, d_in(5) => 
                           NPC_5_port, d_in(4) => NPC_4_port, d_in(3) => 
                           NPC_3_port, d_in(2) => NPC_2_port, d_in(1) => 
                           NPC_1_port, d_in(0) => NPC_0_port, d_out(31) => 
                           NPC1_31_port, d_out(30) => NPC1_30_port, d_out(29) 
                           => NPC1_29_port, d_out(28) => NPC1_28_port, 
                           d_out(27) => NPC1_27_port, d_out(26) => NPC1_26_port
                           , d_out(25) => NPC1_25_port, d_out(24) => 
                           NPC1_24_port, d_out(23) => NPC1_23_port, d_out(22) 
                           => NPC1_22_port, d_out(21) => NPC1_21_port, 
                           d_out(20) => NPC1_20_port, d_out(19) => NPC1_19_port
                           , d_out(18) => NPC1_18_port, d_out(17) => 
                           NPC1_17_port, d_out(16) => NPC1_16_port, d_out(15) 
                           => NPC1_15_port, d_out(14) => NPC1_14_port, 
                           d_out(13) => NPC1_13_port, d_out(12) => NPC1_12_port
                           , d_out(11) => NPC1_11_port, d_out(10) => 
                           NPC1_10_port, d_out(9) => NPC1_9_port, d_out(8) => 
                           NPC1_8_port, d_out(7) => NPC1_7_port, d_out(6) => 
                           NPC1_6_port, d_out(5) => NPC1_5_port, d_out(4) => 
                           NPC1_4_port, d_out(3) => NPC1_3_port, d_out(2) => 
                           NPC1_2_port, d_out(1) => NPC1_1_port, d_out(0) => 
                           NPC1_0_port);
   NPCreg2 : reg_N32_3 port map( clk => Clk, rst => n452, d_in(31) => 
                           NPC1_31_port, d_in(30) => NPC1_30_port, d_in(29) => 
                           NPC1_29_port, d_in(28) => NPC1_28_port, d_in(27) => 
                           NPC1_27_port, d_in(26) => NPC1_26_port, d_in(25) => 
                           NPC1_25_port, d_in(24) => NPC1_24_port, d_in(23) => 
                           NPC1_23_port, d_in(22) => NPC1_22_port, d_in(21) => 
                           NPC1_21_port, d_in(20) => NPC1_20_port, d_in(19) => 
                           NPC1_19_port, d_in(18) => NPC1_18_port, d_in(17) => 
                           NPC1_17_port, d_in(16) => NPC1_16_port, d_in(15) => 
                           NPC1_15_port, d_in(14) => NPC1_14_port, d_in(13) => 
                           NPC1_13_port, d_in(12) => NPC1_12_port, d_in(11) => 
                           NPC1_11_port, d_in(10) => NPC1_10_port, d_in(9) => 
                           NPC1_9_port, d_in(8) => NPC1_8_port, d_in(7) => 
                           NPC1_7_port, d_in(6) => NPC1_6_port, d_in(5) => 
                           NPC1_5_port, d_in(4) => NPC1_4_port, d_in(3) => 
                           NPC1_3_port, d_in(2) => NPC1_2_port, d_in(1) => 
                           NPC1_1_port, d_in(0) => NPC1_0_port, d_out(31) => 
                           NPC2_31_port, d_out(30) => NPC2_30_port, d_out(29) 
                           => NPC2_29_port, d_out(28) => NPC2_28_port, 
                           d_out(27) => NPC2_27_port, d_out(26) => NPC2_26_port
                           , d_out(25) => NPC2_25_port, d_out(24) => 
                           NPC2_24_port, d_out(23) => NPC2_23_port, d_out(22) 
                           => NPC2_22_port, d_out(21) => NPC2_21_port, 
                           d_out(20) => NPC2_20_port, d_out(19) => NPC2_19_port
                           , d_out(18) => NPC2_18_port, d_out(17) => 
                           NPC2_17_port, d_out(16) => NPC2_16_port, d_out(15) 
                           => NPC2_15_port, d_out(14) => NPC2_14_port, 
                           d_out(13) => NPC2_13_port, d_out(12) => NPC2_12_port
                           , d_out(11) => NPC2_11_port, d_out(10) => 
                           NPC2_10_port, d_out(9) => NPC2_9_port, d_out(8) => 
                           NPC2_8_port, d_out(7) => NPC2_7_port, d_out(6) => 
                           NPC2_6_port, d_out(5) => NPC2_5_port, d_out(4) => 
                           NPC2_4_port, d_out(3) => NPC2_3_port, d_out(2) => 
                           NPC2_2_port, d_out(1) => NPC2_1_port, d_out(0) => 
                           NPC2_0_port);
   NPCreg3 : reg_N32_2 port map( clk => Clk, rst => n452, d_in(31) => 
                           NPC2_31_port, d_in(30) => NPC2_30_port, d_in(29) => 
                           NPC2_29_port, d_in(28) => NPC2_28_port, d_in(27) => 
                           NPC2_27_port, d_in(26) => NPC2_26_port, d_in(25) => 
                           NPC2_25_port, d_in(24) => NPC2_24_port, d_in(23) => 
                           NPC2_23_port, d_in(22) => NPC2_22_port, d_in(21) => 
                           NPC2_21_port, d_in(20) => NPC2_20_port, d_in(19) => 
                           NPC2_19_port, d_in(18) => NPC2_18_port, d_in(17) => 
                           NPC2_17_port, d_in(16) => NPC2_16_port, d_in(15) => 
                           NPC2_15_port, d_in(14) => NPC2_14_port, d_in(13) => 
                           NPC2_13_port, d_in(12) => NPC2_12_port, d_in(11) => 
                           NPC2_11_port, d_in(10) => NPC2_10_port, d_in(9) => 
                           NPC2_9_port, d_in(8) => NPC2_8_port, d_in(7) => 
                           NPC2_7_port, d_in(6) => NPC2_6_port, d_in(5) => 
                           NPC2_5_port, d_in(4) => NPC2_4_port, d_in(3) => 
                           NPC2_3_port, d_in(2) => NPC2_2_port, d_in(1) => 
                           NPC2_1_port, d_in(0) => NPC2_0_port, d_out(31) => 
                           NPC3_31_port, d_out(30) => NPC3_30_port, d_out(29) 
                           => NPC3_29_port, d_out(28) => NPC3_28_port, 
                           d_out(27) => NPC3_27_port, d_out(26) => NPC3_26_port
                           , d_out(25) => NPC3_25_port, d_out(24) => 
                           NPC3_24_port, d_out(23) => NPC3_23_port, d_out(22) 
                           => NPC3_22_port, d_out(21) => NPC3_21_port, 
                           d_out(20) => NPC3_20_port, d_out(19) => NPC3_19_port
                           , d_out(18) => NPC3_18_port, d_out(17) => 
                           NPC3_17_port, d_out(16) => NPC3_16_port, d_out(15) 
                           => NPC3_15_port, d_out(14) => NPC3_14_port, 
                           d_out(13) => NPC3_13_port, d_out(12) => NPC3_12_port
                           , d_out(11) => NPC3_11_port, d_out(10) => 
                           NPC3_10_port, d_out(9) => NPC3_9_port, d_out(8) => 
                           NPC3_8_port, d_out(7) => NPC3_7_port, d_out(6) => 
                           NPC3_6_port, d_out(5) => NPC3_5_port, d_out(4) => 
                           NPC3_4_port, d_out(3) => NPC3_3_port, d_out(2) => 
                           NPC3_2_port, d_out(1) => NPC3_1_port, d_out(0) => 
                           NPC3_0_port);
   NPCreg4 : reg_N32_1 port map( clk => Clk, rst => n452, d_in(31) => 
                           NPC3_31_port, d_in(30) => NPC3_30_port, d_in(29) => 
                           NPC3_29_port, d_in(28) => NPC3_28_port, d_in(27) => 
                           NPC3_27_port, d_in(26) => NPC3_26_port, d_in(25) => 
                           NPC3_25_port, d_in(24) => NPC3_24_port, d_in(23) => 
                           NPC3_23_port, d_in(22) => NPC3_22_port, d_in(21) => 
                           NPC3_21_port, d_in(20) => NPC3_20_port, d_in(19) => 
                           NPC3_19_port, d_in(18) => NPC3_18_port, d_in(17) => 
                           NPC3_17_port, d_in(16) => NPC3_16_port, d_in(15) => 
                           NPC3_15_port, d_in(14) => NPC3_14_port, d_in(13) => 
                           NPC3_13_port, d_in(12) => NPC3_12_port, d_in(11) => 
                           NPC3_11_port, d_in(10) => NPC3_10_port, d_in(9) => 
                           NPC3_9_port, d_in(8) => NPC3_8_port, d_in(7) => 
                           NPC3_7_port, d_in(6) => NPC3_6_port, d_in(5) => 
                           NPC3_5_port, d_in(4) => NPC3_4_port, d_in(3) => 
                           NPC3_3_port, d_in(2) => NPC3_2_port, d_in(1) => 
                           NPC3_1_port, d_in(0) => NPC3_0_port, d_out(31) => 
                           NPC4_31_port, d_out(30) => NPC4_30_port, d_out(29) 
                           => NPC4_29_port, d_out(28) => NPC4_28_port, 
                           d_out(27) => NPC4_27_port, d_out(26) => NPC4_26_port
                           , d_out(25) => NPC4_25_port, d_out(24) => 
                           NPC4_24_port, d_out(23) => NPC4_23_port, d_out(22) 
                           => NPC4_22_port, d_out(21) => NPC4_21_port, 
                           d_out(20) => NPC4_20_port, d_out(19) => NPC4_19_port
                           , d_out(18) => NPC4_18_port, d_out(17) => 
                           NPC4_17_port, d_out(16) => NPC4_16_port, d_out(15) 
                           => NPC4_15_port, d_out(14) => NPC4_14_port, 
                           d_out(13) => NPC4_13_port, d_out(12) => NPC4_12_port
                           , d_out(11) => NPC4_11_port, d_out(10) => 
                           NPC4_10_port, d_out(9) => NPC4_9_port, d_out(8) => 
                           NPC4_8_port, d_out(7) => NPC4_7_port, d_out(6) => 
                           NPC4_6_port, d_out(5) => NPC4_5_port, d_out(4) => 
                           NPC4_4_port, d_out(3) => NPC4_3_port, d_out(2) => 
                           NPC4_2_port, d_out(1) => NPC4_1_port, d_out(0) => 
                           NPC4_0_port);
   JUMPENREG1 : ff_0 port map( clk => Clk, rst => n452, d_in => JUMP_EN, d_out 
                           => JUMP_EN1);
   JUMPENREG2 : ff_31 port map( clk => Clk, rst => n452, d_in => JUMP_EN1, 
                           d_out => JUMP_EN2);
   forward_branchREG1 : ff_30 port map( clk => Clk, rst => n453, d_in => 
                           forward_branch, d_out => forward_branch1);
   forward_branchREG2 : ff_29 port map( clk => Clk, rst => n453, d_in => 
                           forward_branch1, d_out => forward_branch2);
   pc_mux : mux_pc port map( A(31) => NPC_31_port, A(30) => NPC_30_port, A(29) 
                           => NPC_29_port, A(28) => NPC_28_port, A(27) => 
                           NPC_27_port, A(26) => NPC_26_port, A(25) => 
                           NPC_25_port, A(24) => NPC_24_port, A(23) => 
                           NPC_23_port, A(22) => NPC_22_port, A(21) => 
                           NPC_21_port, A(20) => NPC_20_port, A(19) => 
                           NPC_19_port, A(18) => NPC_18_port, A(17) => 
                           NPC_17_port, A(16) => NPC_16_port, A(15) => 
                           NPC_15_port, A(14) => NPC_14_port, A(13) => 
                           NPC_13_port, A(12) => NPC_12_port, A(11) => 
                           NPC_11_port, A(10) => NPC_10_port, A(9) => 
                           NPC_9_port, A(8) => NPC_8_port, A(7) => NPC_7_port, 
                           A(6) => NPC_6_port, A(5) => NPC_5_port, A(4) => 
                           NPC_4_port, A(3) => NPC_3_port, A(2) => NPC_2_port, 
                           A(1) => NPC_1_port, A(0) => NPC_0_port, B(31) => 
                           PC_displaced_31_port, B(30) => PC_displaced_30_port,
                           B(29) => PC_displaced_29_port, B(28) => 
                           PC_displaced_28_port, B(27) => PC_displaced_27_port,
                           B(26) => PC_displaced_26_port, B(25) => 
                           PC_displaced_25_port, B(24) => PC_displaced_24_port,
                           B(23) => PC_displaced_23_port, B(22) => 
                           PC_displaced_22_port, B(21) => PC_displaced_21_port,
                           B(20) => PC_displaced_20_port, B(19) => 
                           PC_displaced_19_port, B(18) => PC_displaced_18_port,
                           B(17) => PC_displaced_17_port, B(16) => 
                           PC_displaced_16_port, B(15) => PC_displaced_15_port,
                           B(14) => PC_displaced_14_port, B(13) => 
                           PC_displaced_13_port, B(12) => PC_displaced_12_port,
                           B(11) => PC_displaced_11_port, B(10) => 
                           PC_displaced_10_port, B(9) => PC_displaced_9_port, 
                           B(8) => PC_displaced_8_port, B(7) => 
                           PC_displaced_7_port, B(6) => PC_displaced_6_port, 
                           B(5) => PC_displaced_5_port, B(4) => 
                           PC_displaced_4_port, B(3) => PC_displaced_3_port, 
                           B(2) => PC_displaced_2_port, B(1) => 
                           PC_displaced_1_port, B(0) => PC_displaced_0_port, 
                           C(31) => RF_out_A_FWD_31_port, C(30) => 
                           RF_out_A_FWD_30_port, C(29) => RF_out_A_FWD_29_port,
                           C(28) => RF_out_A_FWD_28_port, C(27) => 
                           RF_out_A_FWD_27_port, C(26) => RF_out_A_FWD_26_port,
                           C(25) => RF_out_A_FWD_25_port, C(24) => 
                           RF_out_A_FWD_24_port, C(23) => RF_out_A_FWD_23_port,
                           C(22) => RF_out_A_FWD_22_port, C(21) => 
                           RF_out_A_FWD_21_port, C(20) => RF_out_A_FWD_20_port,
                           C(19) => RF_out_A_FWD_19_port, C(18) => 
                           RF_out_A_FWD_18_port, C(17) => RF_out_A_FWD_17_port,
                           C(16) => RF_out_A_FWD_16_port, C(15) => 
                           RF_out_A_FWD_15_port, C(14) => RF_out_A_FWD_14_port,
                           C(13) => RF_out_A_FWD_13_port, C(12) => 
                           RF_out_A_FWD_12_port, C(11) => RF_out_A_FWD_11_port,
                           C(10) => RF_out_A_FWD_10_port, C(9) => 
                           RF_out_A_FWD_9_port, C(8) => RF_out_A_FWD_8_port, 
                           C(7) => RF_out_A_FWD_7_port, C(6) => 
                           RF_out_A_FWD_6_port, C(5) => RF_out_A_FWD_5_port, 
                           C(4) => RF_out_A_FWD_4_port, C(3) => 
                           RF_out_A_FWD_3_port, C(2) => RF_out_A_FWD_2_port, 
                           C(1) => RF_out_A_FWD_1_port, C(0) => 
                           RF_out_A_FWD_0_port, D(31) => NPC2_31_port, D(30) =>
                           NPC2_30_port, D(29) => NPC2_29_port, D(28) => 
                           NPC2_28_port, D(27) => NPC2_27_port, D(26) => 
                           NPC2_26_port, D(25) => NPC2_25_port, D(24) => 
                           NPC2_24_port, D(23) => NPC2_23_port, D(22) => 
                           NPC2_22_port, D(21) => NPC2_21_port, D(20) => 
                           NPC2_20_port, D(19) => NPC2_19_port, D(18) => 
                           NPC2_18_port, D(17) => NPC2_17_port, D(16) => 
                           NPC2_16_port, D(15) => NPC2_15_port, D(14) => 
                           NPC2_14_port, D(13) => NPC2_13_port, D(12) => 
                           NPC2_12_port, D(11) => NPC2_11_port, D(10) => 
                           NPC2_10_port, D(9) => NPC2_9_port, D(8) => 
                           NPC2_8_port, D(7) => NPC2_7_port, D(6) => 
                           NPC2_6_port, D(5) => NPC2_5_port, D(4) => 
                           NPC2_4_port, D(3) => NPC2_3_port, D(2) => 
                           NPC2_2_port, D(1) => NPC2_1_port, D(0) => 
                           NPC2_0_port, E(31) => ALU_output_FWD_31_port, E(30) 
                           => ALU_output_FWD_30_port, E(29) => 
                           ALU_output_FWD_29_port, E(28) => 
                           ALU_output_FWD_28_port, E(27) => 
                           ALU_output_FWD_27_port, E(26) => 
                           ALU_output_FWD_26_port, E(25) => 
                           ALU_output_FWD_25_port, E(24) => 
                           ALU_output_FWD_24_port, E(23) => 
                           ALU_output_FWD_23_port, E(22) => 
                           ALU_output_FWD_22_port, E(21) => 
                           ALU_output_FWD_21_port, E(20) => 
                           ALU_output_FWD_20_port, E(19) => 
                           ALU_output_FWD_19_port, E(18) => 
                           ALU_output_FWD_18_port, E(17) => 
                           ALU_output_FWD_17_port, E(16) => 
                           ALU_output_FWD_16_port, E(15) => 
                           ALU_output_FWD_15_port, E(14) => 
                           ALU_output_FWD_14_port, E(13) => 
                           ALU_output_FWD_13_port, E(12) => 
                           ALU_output_FWD_12_port, E(11) => 
                           ALU_output_FWD_11_port, E(10) => 
                           ALU_output_FWD_10_port, E(9) => 
                           ALU_output_FWD_9_port, E(8) => ALU_output_FWD_8_port
                           , E(7) => ALU_output_FWD_7_port, E(6) => 
                           ALU_output_FWD_6_port, E(5) => ALU_output_FWD_5_port
                           , E(4) => ALU_output_FWD_4_port, E(3) => 
                           ALU_output_FWD_3_port, E(2) => ALU_output_FWD_2_port
                           , E(1) => ALU_output_FWD_1_port, E(0) => 
                           ALU_output_FWD_0_port, F(31) => NPC2_31_port, F(30) 
                           => NPC2_30_port, F(29) => NPC2_29_port, F(28) => 
                           NPC2_28_port, F(27) => NPC2_27_port, F(26) => 
                           NPC2_26_port, F(25) => NPC2_25_port, F(24) => 
                           NPC2_24_port, F(23) => NPC2_23_port, F(22) => 
                           NPC2_22_port, F(21) => NPC2_21_port, F(20) => 
                           NPC2_20_port, F(19) => NPC2_19_port, F(18) => 
                           NPC2_18_port, F(17) => NPC2_17_port, F(16) => 
                           NPC2_16_port, F(15) => NPC2_15_port, F(14) => 
                           NPC2_14_port, F(13) => NPC2_13_port, F(12) => 
                           NPC2_12_port, F(11) => NPC2_11_port, F(10) => 
                           NPC2_10_port, F(9) => NPC2_9_port, F(8) => 
                           NPC2_8_port, F(7) => NPC2_7_port, F(6) => 
                           NPC2_6_port, F(5) => NPC2_5_port, F(4) => 
                           NPC2_4_port, F(3) => NPC2_3_port, F(2) => 
                           NPC2_2_port, F(1) => NPC2_1_port, F(0) => 
                           NPC2_0_port, sel(2) => PC_mux_sel_2_port, sel(1) => 
                           flush0_0_port, sel(0) => PC_mux_sel_0_port, Y(31) =>
                           PC_reg_in_31_port, Y(30) => PC_reg_in_30_port, Y(29)
                           => PC_reg_in_29_port, Y(28) => PC_reg_in_28_port, 
                           Y(27) => PC_reg_in_27_port, Y(26) => 
                           PC_reg_in_26_port, Y(25) => PC_reg_in_25_port, Y(24)
                           => PC_reg_in_24_port, Y(23) => PC_reg_in_23_port, 
                           Y(22) => PC_reg_in_22_port, Y(21) => 
                           PC_reg_in_21_port, Y(20) => PC_reg_in_20_port, Y(19)
                           => PC_reg_in_19_port, Y(18) => PC_reg_in_18_port, 
                           Y(17) => PC_reg_in_17_port, Y(16) => 
                           PC_reg_in_16_port, Y(15) => PC_reg_in_15_port, Y(14)
                           => PC_reg_in_14_port, Y(13) => PC_reg_in_13_port, 
                           Y(12) => PC_reg_in_12_port, Y(11) => 
                           PC_reg_in_11_port, Y(10) => PC_reg_in_10_port, Y(9) 
                           => PC_reg_in_9_port, Y(8) => PC_reg_in_8_port, Y(7) 
                           => PC_reg_in_7_port, Y(6) => PC_reg_in_6_port, Y(5) 
                           => PC_reg_in_5_port, Y(4) => PC_reg_in_4_port, Y(3) 
                           => PC_reg_in_3_port, Y(2) => PC_reg_in_2_port, Y(1) 
                           => PC_reg_in_1_port, Y(0) => PC_reg_in_0_port);
   flushreg1 : reg_N2_0 port map( clk => Clk, rst => n452, d_in(1) => 
                           flush0_1_port, d_in(0) => flush0_0_port, d_out(1) =>
                           flush_1_port, d_out(0) => flush_0_port);
   flushreg2 : reg_N2_1 port map( clk => Clk, rst => n452, d_in(1) => 
                           flush_1_port, d_in(0) => flush_0_port, d_out(1) => 
                           flush2_1_port, d_out(0) => flush2_0_port);
   pcen1 : ff_28 port map( clk => Clk, rst => n453, d_in => PC_enable, d_out =>
                           PC_enable1);
   cnt : counter port map( clk => Clk, rst => n452, tc => bootstrap);
   JALreg1 : ff_27 port map( clk => Clk, rst => n453, d_in => JAL_op, d_out => 
                           JAL_op1);
   JALreg2 : ff_26 port map( clk => Clk, rst => n453, d_in => JAL_op1, d_out =>
                           JAL_op2);
   JALreg3 : ff_25 port map( clk => Clk, rst => n453, d_in => JAL_op2, d_out =>
                           JAL_op3);
   JALreg4 : ff_24 port map( clk => Clk, rst => n453, d_in => JAL_op3, d_out =>
                           JAL_op4);
   JRreg1 : ff_23 port map( clk => Clk, rst => n453, d_in => JR_op, d_out => 
                           JR_op1);
   BRANCH_opREG1 : ff_22 port map( clk => Clk, rst => n453, d_in => BRANCH_op, 
                           d_out => BRANCH_op1);
   BRANCH_opREG2 : ff_21 port map( clk => Clk, rst => n453, d_in => BRANCH_op1,
                           d_out => BRANCH_op2);
   LOADREG1 : ff_20 port map( clk => Clk, rst => n452, d_in => LOAD_op, d_out 
                           => LOAD_op1);
   LOADREG2 : ff_19 port map( clk => Clk, rst => n452, d_in => LOAD_op1, d_out 
                           => LOAD_op2);
   STOREREG1 : ff_18 port map( clk => Clk, rst => n452, d_in => STORE_op, d_out
                           => STORE_op1);
   STOREREG2 : ff_17 port map( clk => Clk, rst => n452, d_in => STORE_op1, 
                           d_out => STORE_op2);
   FWDAREG3 : ff_16 port map( clk => Clk, rst => n452, d_in => FWD_A_mem_dec, 
                           d_out => FWD_A_sel_0_port);
   FWDAREG : ff_15 port map( clk => Clk, rst => n452, d_in => FWD_A_exe_dec, 
                           d_out => FWD_A_sel_2_port);
   FWDAREG2 : ff_14 port map( clk => Clk, rst => n452, d_in => FWD_A_wb_dec, 
                           d_out => FWD_A_sel_1_port);
   FWDAMUX : mux_fwd_0 port map( OP(31) => ALU_operand_1_31_port, OP(30) => 
                           ALU_operand_1_30_port, OP(29) => 
                           ALU_operand_1_29_port, OP(28) => 
                           ALU_operand_1_28_port, OP(27) => 
                           ALU_operand_1_27_port, OP(26) => 
                           ALU_operand_1_26_port, OP(25) => 
                           ALU_operand_1_25_port, OP(24) => 
                           ALU_operand_1_24_port, OP(23) => 
                           ALU_operand_1_23_port, OP(22) => 
                           ALU_operand_1_22_port, OP(21) => 
                           ALU_operand_1_21_port, OP(20) => 
                           ALU_operand_1_20_port, OP(19) => 
                           ALU_operand_1_19_port, OP(18) => 
                           ALU_operand_1_18_port, OP(17) => 
                           ALU_operand_1_17_port, OP(16) => 
                           ALU_operand_1_16_port, OP(15) => 
                           ALU_operand_1_15_port, OP(14) => 
                           ALU_operand_1_14_port, OP(13) => 
                           ALU_operand_1_13_port, OP(12) => 
                           ALU_operand_1_12_port, OP(11) => 
                           ALU_operand_1_11_port, OP(10) => 
                           ALU_operand_1_10_port, OP(9) => ALU_operand_1_9_port
                           , OP(8) => ALU_operand_1_8_port, OP(7) => 
                           ALU_operand_1_7_port, OP(6) => ALU_operand_1_6_port,
                           OP(5) => ALU_operand_1_5_port, OP(4) => 
                           ALU_operand_1_4_port, OP(3) => ALU_operand_1_3_port,
                           OP(2) => ALU_operand_1_2_port, OP(1) => 
                           ALU_operand_1_1_port, OP(0) => ALU_operand_1_0_port,
                           alu_out(31) => ALU_reg_out_31_port, alu_out(30) => 
                           ALU_reg_out_30_port, alu_out(29) => 
                           ALU_reg_out_29_port, alu_out(28) => 
                           ALU_reg_out_28_port, alu_out(27) => 
                           ALU_reg_out_27_port, alu_out(26) => 
                           ALU_reg_out_26_port, alu_out(25) => 
                           ALU_reg_out_25_port, alu_out(24) => 
                           ALU_reg_out_24_port, alu_out(23) => 
                           ALU_reg_out_23_port, alu_out(22) => 
                           ALU_reg_out_22_port, alu_out(21) => 
                           ALU_reg_out_21_port, alu_out(20) => 
                           ALU_reg_out_20_port, alu_out(19) => 
                           ALU_reg_out_19_port, alu_out(18) => 
                           ALU_reg_out_18_port, alu_out(17) => 
                           ALU_reg_out_17_port, alu_out(16) => 
                           ALU_reg_out_16_port, alu_out(15) => 
                           ALU_reg_out_15_port, alu_out(14) => 
                           ALU_reg_out_14_port, alu_out(13) => 
                           ALU_reg_out_13_port, alu_out(12) => 
                           ALU_reg_out_12_port, alu_out(11) => 
                           ALU_reg_out_11_port, alu_out(10) => 
                           ALU_reg_out_10_port, alu_out(9) => 
                           ALU_reg_out_9_port, alu_out(8) => ALU_reg_out_8_port
                           , alu_out(7) => ALU_reg_out_7_port, alu_out(6) => 
                           ALU_reg_out_6_port, alu_out(5) => ALU_reg_out_5_port
                           , alu_out(4) => ALU_reg_out_4_port, alu_out(3) => 
                           ALU_reg_out_3_port, alu_out(2) => ALU_reg_out_2_port
                           , alu_out(1) => ALU_reg_out_1_port, alu_out(0) => 
                           ALU_reg_out_0_port, alu_wb_in(31) => 
                           ALU_WB_out_31_port, alu_wb_in(30) => 
                           ALU_WB_out_30_port, alu_wb_in(29) => 
                           ALU_WB_out_29_port, alu_wb_in(28) => 
                           ALU_WB_out_28_port, alu_wb_in(27) => 
                           ALU_WB_out_27_port, alu_wb_in(26) => 
                           ALU_WB_out_26_port, alu_wb_in(25) => 
                           ALU_WB_out_25_port, alu_wb_in(24) => 
                           ALU_WB_out_24_port, alu_wb_in(23) => 
                           ALU_WB_out_23_port, alu_wb_in(22) => 
                           ALU_WB_out_22_port, alu_wb_in(21) => 
                           ALU_WB_out_21_port, alu_wb_in(20) => 
                           ALU_WB_out_20_port, alu_wb_in(19) => 
                           ALU_WB_out_19_port, alu_wb_in(18) => 
                           ALU_WB_out_18_port, alu_wb_in(17) => 
                           ALU_WB_out_17_port, alu_wb_in(16) => 
                           ALU_WB_out_16_port, alu_wb_in(15) => 
                           ALU_WB_out_15_port, alu_wb_in(14) => 
                           ALU_WB_out_14_port, alu_wb_in(13) => 
                           ALU_WB_out_13_port, alu_wb_in(12) => 
                           ALU_WB_out_12_port, alu_wb_in(11) => 
                           ALU_WB_out_11_port, alu_wb_in(10) => 
                           ALU_WB_out_10_port, alu_wb_in(9) => 
                           ALU_WB_out_9_port, alu_wb_in(8) => ALU_WB_out_8_port
                           , alu_wb_in(7) => ALU_WB_out_7_port, alu_wb_in(6) =>
                           ALU_WB_out_6_port, alu_wb_in(5) => ALU_WB_out_5_port
                           , alu_wb_in(4) => ALU_WB_out_4_port, alu_wb_in(3) =>
                           ALU_WB_out_3_port, alu_wb_in(2) => ALU_WB_out_2_port
                           , alu_wb_in(1) => ALU_WB_out_1_port, alu_wb_in(0) =>
                           ALU_WB_out_0_port, lmd_out(31) => 
                           LMD_reg_out_31_port, lmd_out(30) => 
                           LMD_reg_out_30_port, lmd_out(29) => 
                           LMD_reg_out_29_port, lmd_out(28) => 
                           LMD_reg_out_28_port, lmd_out(27) => 
                           LMD_reg_out_27_port, lmd_out(26) => 
                           LMD_reg_out_26_port, lmd_out(25) => 
                           LMD_reg_out_25_port, lmd_out(24) => 
                           LMD_reg_out_24_port, lmd_out(23) => 
                           LMD_reg_out_23_port, lmd_out(22) => 
                           LMD_reg_out_22_port, lmd_out(21) => 
                           LMD_reg_out_21_port, lmd_out(20) => 
                           LMD_reg_out_20_port, lmd_out(19) => 
                           LMD_reg_out_19_port, lmd_out(18) => 
                           LMD_reg_out_18_port, lmd_out(17) => 
                           LMD_reg_out_17_port, lmd_out(16) => 
                           LMD_reg_out_16_port, lmd_out(15) => 
                           LMD_reg_out_15_port, lmd_out(14) => 
                           LMD_reg_out_14_port, lmd_out(13) => 
                           LMD_reg_out_13_port, lmd_out(12) => 
                           LMD_reg_out_12_port, lmd_out(11) => 
                           LMD_reg_out_11_port, lmd_out(10) => 
                           LMD_reg_out_10_port, lmd_out(9) => 
                           LMD_reg_out_9_port, lmd_out(8) => LMD_reg_out_8_port
                           , lmd_out(7) => LMD_reg_out_7_port, lmd_out(6) => 
                           LMD_reg_out_6_port, lmd_out(5) => LMD_reg_out_5_port
                           , lmd_out(4) => LMD_reg_out_4_port, lmd_out(3) => 
                           LMD_reg_out_3_port, lmd_out(2) => LMD_reg_out_2_port
                           , lmd_out(1) => LMD_reg_out_1_port, lmd_out(0) => 
                           LMD_reg_out_0_port, OPF(31) => 
                           ALU_operand_1_FWD_31_port, OPF(30) => 
                           ALU_operand_1_FWD_30_port, OPF(29) => 
                           ALU_operand_1_FWD_29_port, OPF(28) => 
                           ALU_operand_1_FWD_28_port, OPF(27) => 
                           ALU_operand_1_FWD_27_port, OPF(26) => 
                           ALU_operand_1_FWD_26_port, OPF(25) => 
                           ALU_operand_1_FWD_25_port, OPF(24) => 
                           ALU_operand_1_FWD_24_port, OPF(23) => 
                           ALU_operand_1_FWD_23_port, OPF(22) => 
                           ALU_operand_1_FWD_22_port, OPF(21) => 
                           ALU_operand_1_FWD_21_port, OPF(20) => 
                           ALU_operand_1_FWD_20_port, OPF(19) => 
                           ALU_operand_1_FWD_19_port, OPF(18) => 
                           ALU_operand_1_FWD_18_port, OPF(17) => 
                           ALU_operand_1_FWD_17_port, OPF(16) => 
                           ALU_operand_1_FWD_16_port, OPF(15) => 
                           ALU_operand_1_FWD_15_port, OPF(14) => 
                           ALU_operand_1_FWD_14_port, OPF(13) => 
                           ALU_operand_1_FWD_13_port, OPF(12) => 
                           ALU_operand_1_FWD_12_port, OPF(11) => 
                           ALU_operand_1_FWD_11_port, OPF(10) => 
                           ALU_operand_1_FWD_10_port, OPF(9) => 
                           ALU_operand_1_FWD_9_port, OPF(8) => 
                           ALU_operand_1_FWD_8_port, OPF(7) => 
                           ALU_operand_1_FWD_7_port, OPF(6) => 
                           ALU_operand_1_FWD_6_port, OPF(5) => 
                           ALU_operand_1_FWD_5_port, OPF(4) => 
                           ALU_operand_1_FWD_4_port, OPF(3) => 
                           ALU_operand_1_FWD_3_port, OPF(2) => 
                           ALU_operand_1_FWD_2_port, OPF(1) => 
                           ALU_operand_1_FWD_1_port, OPF(0) => 
                           ALU_operand_1_FWD_0_port, sel(2) => FWD_A_sel_2_port
                           , sel(1) => FWD_A_sel_1_port, sel(0) => 
                           FWD_A_sel_0_port);
   FWDBREG3a : ff_13 port map( clk => Clk, rst => n452, d_in => FWD_B_mem_exe, 
                           d_out => FWD_B_sel_0_port);
   FWDBREG : ff_12 port map( clk => Clk, rst => n452, d_in => FWD_B_exe_dec, 
                           d_out => FWD_B_sel_2_port);
   FWDBREG2 : ff_11 port map( clk => Clk, rst => n452, d_in => FWD_B_wb_dec, 
                           d_out => FWD_B_sel_1_port);
   FWDBMUX : mux_fwd_1 port map( OP(31) => ALU_operand_2_31_port, OP(30) => 
                           ALU_operand_2_30_port, OP(29) => 
                           ALU_operand_2_29_port, OP(28) => 
                           ALU_operand_2_28_port, OP(27) => 
                           ALU_operand_2_27_port, OP(26) => 
                           ALU_operand_2_26_port, OP(25) => 
                           ALU_operand_2_25_port, OP(24) => 
                           ALU_operand_2_24_port, OP(23) => 
                           ALU_operand_2_23_port, OP(22) => 
                           ALU_operand_2_22_port, OP(21) => 
                           ALU_operand_2_21_port, OP(20) => 
                           ALU_operand_2_20_port, OP(19) => 
                           ALU_operand_2_19_port, OP(18) => 
                           ALU_operand_2_18_port, OP(17) => 
                           ALU_operand_2_17_port, OP(16) => 
                           ALU_operand_2_16_port, OP(15) => 
                           ALU_operand_2_15_port, OP(14) => 
                           ALU_operand_2_14_port, OP(13) => 
                           ALU_operand_2_13_port, OP(12) => 
                           ALU_operand_2_12_port, OP(11) => 
                           ALU_operand_2_11_port, OP(10) => 
                           ALU_operand_2_10_port, OP(9) => ALU_operand_2_9_port
                           , OP(8) => ALU_operand_2_8_port, OP(7) => 
                           ALU_operand_2_7_port, OP(6) => ALU_operand_2_6_port,
                           OP(5) => ALU_operand_2_5_port, OP(4) => 
                           ALU_operand_2_4_port, OP(3) => ALU_operand_2_3_port,
                           OP(2) => ALU_operand_2_2_port, OP(1) => 
                           ALU_operand_2_1_port, OP(0) => ALU_operand_2_0_port,
                           alu_out(31) => ALU_reg_out_31_port, alu_out(30) => 
                           ALU_reg_out_30_port, alu_out(29) => 
                           ALU_reg_out_29_port, alu_out(28) => 
                           ALU_reg_out_28_port, alu_out(27) => 
                           ALU_reg_out_27_port, alu_out(26) => 
                           ALU_reg_out_26_port, alu_out(25) => 
                           ALU_reg_out_25_port, alu_out(24) => 
                           ALU_reg_out_24_port, alu_out(23) => 
                           ALU_reg_out_23_port, alu_out(22) => 
                           ALU_reg_out_22_port, alu_out(21) => 
                           ALU_reg_out_21_port, alu_out(20) => 
                           ALU_reg_out_20_port, alu_out(19) => 
                           ALU_reg_out_19_port, alu_out(18) => 
                           ALU_reg_out_18_port, alu_out(17) => 
                           ALU_reg_out_17_port, alu_out(16) => 
                           ALU_reg_out_16_port, alu_out(15) => 
                           ALU_reg_out_15_port, alu_out(14) => 
                           ALU_reg_out_14_port, alu_out(13) => 
                           ALU_reg_out_13_port, alu_out(12) => 
                           ALU_reg_out_12_port, alu_out(11) => 
                           ALU_reg_out_11_port, alu_out(10) => 
                           ALU_reg_out_10_port, alu_out(9) => 
                           ALU_reg_out_9_port, alu_out(8) => ALU_reg_out_8_port
                           , alu_out(7) => ALU_reg_out_7_port, alu_out(6) => 
                           ALU_reg_out_6_port, alu_out(5) => ALU_reg_out_5_port
                           , alu_out(4) => ALU_reg_out_4_port, alu_out(3) => 
                           ALU_reg_out_3_port, alu_out(2) => ALU_reg_out_2_port
                           , alu_out(1) => ALU_reg_out_1_port, alu_out(0) => 
                           ALU_reg_out_0_port, alu_wb_in(31) => 
                           ALU_WB_out_31_port, alu_wb_in(30) => 
                           ALU_WB_out_30_port, alu_wb_in(29) => 
                           ALU_WB_out_29_port, alu_wb_in(28) => 
                           ALU_WB_out_28_port, alu_wb_in(27) => 
                           ALU_WB_out_27_port, alu_wb_in(26) => 
                           ALU_WB_out_26_port, alu_wb_in(25) => 
                           ALU_WB_out_25_port, alu_wb_in(24) => 
                           ALU_WB_out_24_port, alu_wb_in(23) => 
                           ALU_WB_out_23_port, alu_wb_in(22) => 
                           ALU_WB_out_22_port, alu_wb_in(21) => 
                           ALU_WB_out_21_port, alu_wb_in(20) => 
                           ALU_WB_out_20_port, alu_wb_in(19) => 
                           ALU_WB_out_19_port, alu_wb_in(18) => 
                           ALU_WB_out_18_port, alu_wb_in(17) => 
                           ALU_WB_out_17_port, alu_wb_in(16) => 
                           ALU_WB_out_16_port, alu_wb_in(15) => 
                           ALU_WB_out_15_port, alu_wb_in(14) => 
                           ALU_WB_out_14_port, alu_wb_in(13) => 
                           ALU_WB_out_13_port, alu_wb_in(12) => 
                           ALU_WB_out_12_port, alu_wb_in(11) => 
                           ALU_WB_out_11_port, alu_wb_in(10) => 
                           ALU_WB_out_10_port, alu_wb_in(9) => 
                           ALU_WB_out_9_port, alu_wb_in(8) => ALU_WB_out_8_port
                           , alu_wb_in(7) => ALU_WB_out_7_port, alu_wb_in(6) =>
                           ALU_WB_out_6_port, alu_wb_in(5) => ALU_WB_out_5_port
                           , alu_wb_in(4) => ALU_WB_out_4_port, alu_wb_in(3) =>
                           ALU_WB_out_3_port, alu_wb_in(2) => ALU_WB_out_2_port
                           , alu_wb_in(1) => ALU_WB_out_1_port, alu_wb_in(0) =>
                           ALU_WB_out_0_port, lmd_out(31) => 
                           LMD_reg_out_31_port, lmd_out(30) => 
                           LMD_reg_out_30_port, lmd_out(29) => 
                           LMD_reg_out_29_port, lmd_out(28) => 
                           LMD_reg_out_28_port, lmd_out(27) => 
                           LMD_reg_out_27_port, lmd_out(26) => 
                           LMD_reg_out_26_port, lmd_out(25) => 
                           LMD_reg_out_25_port, lmd_out(24) => 
                           LMD_reg_out_24_port, lmd_out(23) => 
                           LMD_reg_out_23_port, lmd_out(22) => 
                           LMD_reg_out_22_port, lmd_out(21) => 
                           LMD_reg_out_21_port, lmd_out(20) => 
                           LMD_reg_out_20_port, lmd_out(19) => 
                           LMD_reg_out_19_port, lmd_out(18) => 
                           LMD_reg_out_18_port, lmd_out(17) => 
                           LMD_reg_out_17_port, lmd_out(16) => 
                           LMD_reg_out_16_port, lmd_out(15) => 
                           LMD_reg_out_15_port, lmd_out(14) => 
                           LMD_reg_out_14_port, lmd_out(13) => 
                           LMD_reg_out_13_port, lmd_out(12) => 
                           LMD_reg_out_12_port, lmd_out(11) => 
                           LMD_reg_out_11_port, lmd_out(10) => 
                           LMD_reg_out_10_port, lmd_out(9) => 
                           LMD_reg_out_9_port, lmd_out(8) => LMD_reg_out_8_port
                           , lmd_out(7) => LMD_reg_out_7_port, lmd_out(6) => 
                           LMD_reg_out_6_port, lmd_out(5) => LMD_reg_out_5_port
                           , lmd_out(4) => LMD_reg_out_4_port, lmd_out(3) => 
                           LMD_reg_out_3_port, lmd_out(2) => LMD_reg_out_2_port
                           , lmd_out(1) => LMD_reg_out_1_port, lmd_out(0) => 
                           LMD_reg_out_0_port, OPF(31) => 
                           ALU_operand_2_FWD_31_port, OPF(30) => 
                           ALU_operand_2_FWD_30_port, OPF(29) => 
                           ALU_operand_2_FWD_29_port, OPF(28) => 
                           ALU_operand_2_FWD_28_port, OPF(27) => 
                           ALU_operand_2_FWD_27_port, OPF(26) => 
                           ALU_operand_2_FWD_26_port, OPF(25) => 
                           ALU_operand_2_FWD_25_port, OPF(24) => 
                           ALU_operand_2_FWD_24_port, OPF(23) => 
                           ALU_operand_2_FWD_23_port, OPF(22) => 
                           ALU_operand_2_FWD_22_port, OPF(21) => 
                           ALU_operand_2_FWD_21_port, OPF(20) => 
                           ALU_operand_2_FWD_20_port, OPF(19) => 
                           ALU_operand_2_FWD_19_port, OPF(18) => 
                           ALU_operand_2_FWD_18_port, OPF(17) => 
                           ALU_operand_2_FWD_17_port, OPF(16) => 
                           ALU_operand_2_FWD_16_port, OPF(15) => 
                           ALU_operand_2_FWD_15_port, OPF(14) => 
                           ALU_operand_2_FWD_14_port, OPF(13) => 
                           ALU_operand_2_FWD_13_port, OPF(12) => 
                           ALU_operand_2_FWD_12_port, OPF(11) => 
                           ALU_operand_2_FWD_11_port, OPF(10) => 
                           ALU_operand_2_FWD_10_port, OPF(9) => 
                           ALU_operand_2_FWD_9_port, OPF(8) => 
                           ALU_operand_2_FWD_8_port, OPF(7) => 
                           ALU_operand_2_FWD_7_port, OPF(6) => 
                           ALU_operand_2_FWD_6_port, OPF(5) => 
                           ALU_operand_2_FWD_5_port, OPF(4) => 
                           ALU_operand_2_FWD_4_port, OPF(3) => 
                           ALU_operand_2_FWD_3_port, OPF(2) => 
                           ALU_operand_2_FWD_2_port, OPF(1) => 
                           ALU_operand_2_FWD_1_port, OPF(0) => 
                           ALU_operand_2_FWD_0_port, sel(2) => FWD_B_sel_2_port
                           , sel(1) => FWD_B_sel_1_port, sel(0) => 
                           FWD_B_sel_0_port);
   FWDBREG3 : ff_10 port map( clk => Clk, rst => n452, d_in => FWD_B_exe_mem, 
                           d_out => FWD_B_exe_mem1);
   FWDBREG4 : ff_9 port map( clk => Clk, rst => n452, d_in => FWD_B_exe_mem1, 
                           d_out => FWD_B_exe_mem2);
   FWDBREG5 : ff_8 port map( clk => Clk, rst => n452, d_in => FWD_B_wb_mem, 
                           d_out => FWD_B_wb_mem1);
   FWDBREG6 : ff_7 port map( clk => Clk, rst => n452, d_in => FWD_B_wb_mem1, 
                           d_out => FWD_B_wb_mem2);
   FWDBREG7 : ff_6 port map( clk => Clk, rst => n452, d_in => FWD_B_mem_mem, 
                           d_out => FWD_B_mem_mem1);
   FWDBREG8 : ff_5 port map( clk => Clk, rst => n452, d_in => FWD_B_mem_mem1, 
                           d_out => FWD_B_mem_mem2);
   FWDBREG9 : ff_4 port map( clk => Clk, rst => n452, d_in => FWD_B_lmd1_mem, 
                           d_out => FWD_B_lmd1_mem1);
   FWDBREG10 : ff_3 port map( clk => Clk, rst => n452, d_in => FWD_B_lmd1_mem1,
                           d_out => FWD_B_lmd1_mem2);
   FWDBRANCH1 : ff_2 port map( clk => Clk, rst => n452, d_in => FWD_exe_branch,
                           d_out => FWD_exe_branch1);
   FWDBRANCH2 : ff_1 port map( clk => Clk, rst => n452, d_in => FWD_wb_branch, 
                           d_out => FWD_wb_branch1);
   U3 : NOR4_X1 port map( A1 => RD2_3_port, A2 => RD2_4_port, A3 => RD2_2_port,
                           A4 => n342, ZN => n290);
   U4 : BUF_X1 port map( A => n110, Z => n434);
   U5 : BUF_X1 port map( A => n110, Z => n435);
   U6 : INV_X1 port map( A => n449, ZN => n440);
   U7 : BUF_X1 port map( A => n110, Z => n436);
   U8 : BUF_X1 port map( A => n115, Z => n429);
   U9 : BUF_X1 port map( A => n115, Z => n430);
   U10 : BUF_X1 port map( A => n115, Z => n431);
   U11 : BUF_X1 port map( A => n450, Z => n449);
   U12 : NAND2_X1 port map( A1 => n209, A2 => n432, ZN => n110);
   U13 : BUF_X1 port map( A => n446, Z => n447);
   U14 : BUF_X1 port map( A => n445, Z => n448);
   U15 : BUF_X1 port map( A => n450, Z => n445);
   U16 : BUF_X1 port map( A => n450, Z => n446);
   U17 : BUF_X1 port map( A => n450, Z => n444);
   U18 : BUF_X1 port map( A => n450, Z => n441);
   U19 : BUF_X1 port map( A => n450, Z => n443);
   U20 : BUF_X1 port map( A => n450, Z => n442);
   U21 : BUF_X1 port map( A => n355, Z => n210);
   U22 : BUF_X1 port map( A => n355, Z => n312);
   U23 : BUF_X1 port map( A => n355, Z => n313);
   U24 : AOI21_X1 port map( B1 => n106, B2 => n107, A => n108, ZN => 
                           flush0_0_port);
   U25 : INV_X1 port map( A => n97, ZN => n432);
   U26 : INV_X1 port map( A => n97, ZN => n433);
   U27 : NOR2_X1 port map( A1 => n209, A2 => n97, ZN => n115);
   U28 : OAI21_X1 port map( B1 => n218, B2 => PC_enable, A => n107, ZN => n103)
                           ;
   U29 : NOR2_X1 port map( A1 => n212, A2 => n106, ZN => n209);
   U30 : INV_X1 port map( A => n221, ZN => PC_mux_sel_0_port);
   U31 : AOI21_X1 port map( B1 => n106, B2 => n103, A => n108, ZN => n221);
   U32 : INV_X1 port map( A => n104, ZN => PC_mux_sel_2_port);
   U33 : INV_X1 port map( A => n230, ZN => n211);
   U34 : INV_X1 port map( A => n120, ZN => ALU_output_FWD_7_port);
   U35 : INV_X1 port map( A => n162, ZN => ALU_output_FWD_23_port);
   U36 : INV_X1 port map( A => n168, ZN => ALU_output_FWD_21_port);
   U37 : INV_X1 port map( A => n180, ZN => ALU_output_FWD_18_port);
   U38 : INV_X1 port map( A => n186, ZN => ALU_output_FWD_16_port);
   U39 : INV_X1 port map( A => n189, ZN => ALU_output_FWD_15_port);
   U40 : INV_X1 port map( A => n192, ZN => ALU_output_FWD_14_port);
   U41 : INV_X1 port map( A => n195, ZN => ALU_output_FWD_13_port);
   U42 : INV_X1 port map( A => n198, ZN => ALU_output_FWD_12_port);
   U43 : INV_X1 port map( A => n201, ZN => ALU_output_FWD_11_port);
   U44 : INV_X1 port map( A => n204, ZN => ALU_output_FWD_10_port);
   U45 : INV_X1 port map( A => n174, ZN => ALU_output_FWD_1_port);
   U46 : INV_X1 port map( A => n207, ZN => ALU_output_FWD_0_port);
   U47 : INV_X1 port map( A => n147, ZN => ALU_output_FWD_28_port);
   U48 : INV_X1 port map( A => n153, ZN => ALU_output_FWD_26_port);
   U49 : INV_X1 port map( A => n159, ZN => ALU_output_FWD_24_port);
   U50 : INV_X1 port map( A => n165, ZN => ALU_output_FWD_22_port);
   U51 : INV_X1 port map( A => n171, ZN => ALU_output_FWD_20_port);
   U52 : INV_X1 port map( A => n177, ZN => ALU_output_FWD_19_port);
   U53 : INV_X1 port map( A => n183, ZN => ALU_output_FWD_17_port);
   U54 : INV_X1 port map( A => n117, ZN => ALU_output_FWD_8_port);
   U55 : INV_X1 port map( A => n123, ZN => ALU_output_FWD_6_port);
   U56 : INV_X1 port map( A => n129, ZN => ALU_output_FWD_4_port);
   U57 : INV_X1 port map( A => n141, ZN => ALU_output_FWD_2_port);
   U58 : INV_X1 port map( A => n150, ZN => ALU_output_FWD_27_port);
   U59 : INV_X1 port map( A => n156, ZN => ALU_output_FWD_25_port);
   U60 : INV_X1 port map( A => n112, ZN => ALU_output_FWD_9_port);
   U61 : INV_X1 port map( A => n126, ZN => ALU_output_FWD_5_port);
   U62 : INV_X1 port map( A => n132, ZN => ALU_output_FWD_3_port);
   U63 : INV_X1 port map( A => n138, ZN => ALU_output_FWD_30_port);
   U64 : INV_X1 port map( A => n144, ZN => ALU_output_FWD_29_port);
   U65 : INV_X1 port map( A => n135, ZN => ALU_output_FWD_31_port);
   U66 : OAI21_X1 port map( B1 => n103, B2 => n104, A => n105, ZN => 
                           flush0_1_port);
   U67 : INV_X1 port map( A => flush0_0_port, ZN => n105);
   U68 : INV_X1 port map( A => n304, ZN => n303);
   U69 : INV_X1 port map( A => n216, ZN => RD_1_port);
   U70 : INV_X1 port map( A => n215, ZN => RD_2_port);
   U71 : INV_X1 port map( A => n109, ZN => STORE_op);
   U72 : NOR3_X1 port map( A1 => n335, A2 => n290, A3 => n212, ZN => 
                           FWD_A_mem_dec);
   U73 : NOR3_X1 port map( A1 => n327, A2 => n304, A3 => n328, ZN => 
                           FWD_B_exe_dec);
   U74 : INV_X1 port map( A => n308, ZN => FWD_B_lmd1_mem);
   U75 : NOR2_X1 port map( A1 => n230, A2 => n284, ZN => FWD_exe_branch);
   U76 : NOR2_X1 port map( A1 => n212, A2 => n284, ZN => FWD_wb_branch);
   U77 : INV_X1 port map( A => n213, ZN => RD_4_port);
   U78 : INV_X1 port map( A => n217, ZN => RD_0_port);
   U79 : INV_X1 port map( A => n214, ZN => RD_3_port);
   U80 : INV_X1 port map( A => JAL_op2, ZN => n450);
   U81 : BUF_X1 port map( A => n353, Z => n332);
   U82 : BUF_X1 port map( A => n353, Z => n424);
   U83 : NOR2_X1 port map( A1 => n420, A2 => n418, ZN => n355);
   U84 : BUF_X1 port map( A => n354, Z => n314);
   U85 : BUF_X1 port map( A => n354, Z => n330);
   U86 : BUF_X1 port map( A => n352, Z => n426);
   U87 : BUF_X1 port map( A => n352, Z => n427);
   U88 : BUF_X1 port map( A => n353, Z => n425);
   U89 : BUF_X1 port map( A => n354, Z => n331);
   U90 : BUF_X1 port map( A => n352, Z => n428);
   U91 : INV_X1 port map( A => n419, ZN => n418);
   U92 : OAI22_X1 port map( A1 => Instr_reg_out_20_port, A2 => n322, B1 => 
                           Instr_reg_out_15_port, B2 => n304, ZN => n213);
   U93 : OAI22_X1 port map( A1 => Instr_reg_out_19_port, A2 => n322, B1 => 
                           Instr_reg_out_14_port, B2 => n304, ZN => n214);
   U94 : OAI22_X1 port map( A1 => Instr_reg_out_18_port, A2 => n322, B1 => 
                           Instr_reg_out_13_port, B2 => n304, ZN => n215);
   U95 : OAI22_X1 port map( A1 => Instr_reg_out_16_port, A2 => n322, B1 => 
                           Instr_reg_out_11_port, B2 => n304, ZN => n217);
   U96 : OAI22_X1 port map( A1 => Instr_reg_out_17_port, A2 => n322, B1 => 
                           Instr_reg_out_12_port, B2 => n304, ZN => n216);
   U97 : NOR3_X1 port map( A1 => n222, A2 => JR_op, A3 => n223, ZN => n108);
   U98 : AOI21_X1 port map( B1 => Instr(15), B2 => BRANCH_op, A => JUMP_EN, ZN 
                           => n222);
   U99 : INV_X1 port map( A => n224, ZN => n223);
   U100 : OAI221_X1 port map( B1 => n435, B2 => n137, C1 => n138, C2 => n433, A
                           => n139, ZN => RF_out_A_FWD_30_port);
   U101 : OAI221_X1 port map( B1 => n435, B2 => n143, C1 => n144, C2 => n433, A
                           => n145, ZN => RF_out_A_FWD_29_port);
   U102 : OAI221_X1 port map( B1 => n435, B2 => n161, C1 => n162, C2 => n433, A
                           => n163, ZN => RF_out_A_FWD_23_port);
   U103 : OAI221_X1 port map( B1 => n435, B2 => n146, C1 => n147, C2 => n433, A
                           => n148, ZN => RF_out_A_FWD_28_port);
   U104 : OAI221_X1 port map( B1 => n435, B2 => n152, C1 => n153, C2 => n433, A
                           => n154, ZN => RF_out_A_FWD_26_port);
   U105 : OAI221_X1 port map( B1 => n435, B2 => n158, C1 => n159, C2 => n433, A
                           => n160, ZN => RF_out_A_FWD_24_port);
   U106 : OAI221_X1 port map( B1 => n435, B2 => n149, C1 => n150, C2 => n433, A
                           => n151, ZN => RF_out_A_FWD_27_port);
   U107 : OAI221_X1 port map( B1 => n435, B2 => n155, C1 => n156, C2 => n433, A
                           => n157, ZN => RF_out_A_FWD_25_port);
   U108 : NOR4_X1 port map( A1 => ALU_reg_out_22_port, A2 => 
                           ALU_reg_out_21_port, A3 => ALU_reg_out_20_port, A4 
                           => ALU_reg_out_1_port, ZN => n244);
   U109 : NOR4_X1 port map( A1 => A_reg_out_9_port, A2 => A_reg_out_8_port, A3 
                           => A_reg_out_7_port, A4 => A_reg_out_6_port, ZN => 
                           n261);
   U110 : NOR4_X1 port map( A1 => A_reg_out_23_port, A2 => A_reg_out_22_port, 
                           A3 => A_reg_out_21_port, A4 => A_reg_out_20_port, ZN
                           => n265);
   U111 : NOR4_X1 port map( A1 => A_reg_out_5_port, A2 => A_reg_out_4_port, A3 
                           => A_reg_out_3_port, A4 => A_reg_out_31_port, ZN => 
                           n260);
   U112 : NOR4_X1 port map( A1 => A_reg_out_1_port, A2 => A_reg_out_19_port, A3
                           => A_reg_out_18_port, A4 => A_reg_out_17_port, ZN =>
                           n264);
   U113 : AOI21_X1 port map( B1 => n245, B2 => n246, A => n247, ZN => n233);
   U114 : INV_X1 port map( A => FWD_wb_branch1, ZN => n247);
   U115 : NOR4_X1 port map( A1 => n252, A2 => n253, A3 => n254, A4 => n255, ZN 
                           => n245);
   U116 : NOR4_X1 port map( A1 => n248, A2 => n249, A3 => n250, A4 => n251, ZN 
                           => n246);
   U117 : NOR4_X1 port map( A1 => ALU_reg_out_19_port, A2 => 
                           ALU_reg_out_18_port, A3 => ALU_reg_out_17_port, A4 
                           => ALU_reg_out_16_port, ZN => n243);
   U118 : NOR4_X1 port map( A1 => ALU_reg_out_2_port, A2 => ALU_reg_out_29_port
                           , A3 => ALU_reg_out_28_port, A4 => 
                           ALU_reg_out_27_port, ZN => n238);
   U119 : NOR4_X1 port map( A1 => ALU_reg_out_15_port, A2 => 
                           ALU_reg_out_14_port, A3 => ALU_reg_out_13_port, A4 
                           => ALU_reg_out_12_port, ZN => n242);
   U120 : NOR4_X1 port map( A1 => A_reg_out_30_port, A2 => A_reg_out_2_port, A3
                           => A_reg_out_29_port, A4 => A_reg_out_28_port, ZN =>
                           n259);
   U121 : NOR4_X1 port map( A1 => A_reg_out_16_port, A2 => A_reg_out_15_port, 
                           A3 => A_reg_out_14_port, A4 => A_reg_out_13_port, ZN
                           => n263);
   U122 : NOR4_X1 port map( A1 => ALU_reg_out_26_port, A2 => 
                           ALU_reg_out_25_port, A3 => ALU_reg_out_24_port, A4 
                           => ALU_reg_out_23_port, ZN => n237);
   U123 : NOR4_X1 port map( A1 => A_reg_out_27_port, A2 => A_reg_out_26_port, 
                           A3 => A_reg_out_25_port, A4 => A_reg_out_24_port, ZN
                           => n258);
   U124 : BUF_X2 port map( A => Rst, Z => n451);
   U125 : NAND4_X1 port map( A1 => n336, A2 => n337, A3 => n338, A4 => n339, ZN
                           => n212);
   U126 : XNOR2_X1 port map( A => Instr_reg_out_23_port, B => RD2_2_port, ZN =>
                           n336);
   U127 : XNOR2_X1 port map( A => Instr_reg_out_24_port, B => RD2_3_port, ZN =>
                           n338);
   U128 : NOR2_X1 port map( A1 => n340, A2 => n341, ZN => n339);
   U129 : NOR3_X1 port map( A1 => Instr(31), A2 => Instr(29), A3 => n423, ZN =>
                           n282);
   U130 : INV_X1 port map( A => PC_enable1, ZN => n423);
   U131 : NAND2_X1 port map( A1 => n304, A2 => n326, ZN => n322);
   U132 : OR3_X1 port map( A1 => Instr_reg_out_28_port, A2 => 
                           Instr_reg_out_29_port, A3 => n311, ZN => n326);
   U133 : AND2_X1 port map( A1 => ALU_OPCODE(2), A2 => PC_enable1, ZN => 
                           ALU_OPCODE_in_2_port);
   U134 : AOI22_X1 port map( A1 => ALU_output_16_port, A2 => n447, B1 => 
                           NPC2_16_port, B2 => JAL_op2, ZN => n186);
   U135 : AOI22_X1 port map( A1 => ALU_output_15_port, A2 => n447, B1 => 
                           NPC2_15_port, B2 => JAL_op2, ZN => n189);
   U136 : AOI22_X1 port map( A1 => ALU_output_14_port, A2 => n447, B1 => 
                           NPC2_14_port, B2 => JAL_op2, ZN => n192);
   U137 : AOI22_X1 port map( A1 => ALU_output_13_port, A2 => n447, B1 => 
                           NPC2_13_port, B2 => n440, ZN => n195);
   U138 : AOI22_X1 port map( A1 => ALU_output_12_port, A2 => n448, B1 => 
                           NPC2_12_port, B2 => JAL_op2, ZN => n198);
   U139 : AOI22_X1 port map( A1 => ALU_output_11_port, A2 => n448, B1 => 
                           NPC2_11_port, B2 => n440, ZN => n201);
   U140 : AOI22_X1 port map( A1 => ALU_output_10_port, A2 => n448, B1 => 
                           NPC2_10_port, B2 => JAL_op2, ZN => n204);
   U141 : AOI22_X1 port map( A1 => ALU_output_0_port, A2 => n448, B1 => 
                           NPC2_0_port, B2 => n440, ZN => n207);
   U142 : AOI22_X1 port map( A1 => ALU_output_23_port, A2 => n445, B1 => 
                           NPC2_23_port, B2 => n440, ZN => n162);
   U143 : AOI22_X1 port map( A1 => ALU_output_21_port, A2 => n445, B1 => 
                           NPC2_21_port, B2 => n440, ZN => n168);
   U144 : AOI22_X1 port map( A1 => ALU_output_18_port, A2 => n446, B1 => 
                           NPC2_18_port, B2 => n440, ZN => n180);
   U145 : AOI22_X1 port map( A1 => ALU_output_1_port, A2 => n446, B1 => 
                           NPC2_1_port, B2 => n440, ZN => n174);
   U146 : AOI22_X1 port map( A1 => ALU_output_28_port, A2 => n443, B1 => 
                           NPC2_28_port, B2 => JAL_op2, ZN => n147);
   U147 : AOI22_X1 port map( A1 => ALU_output_26_port, A2 => n444, B1 => 
                           NPC2_26_port, B2 => n440, ZN => n153);
   U148 : AOI22_X1 port map( A1 => ALU_output_24_port, A2 => n444, B1 => 
                           NPC2_24_port, B2 => n440, ZN => n159);
   U149 : AOI22_X1 port map( A1 => ALU_output_22_port, A2 => n445, B1 => 
                           NPC2_22_port, B2 => n440, ZN => n165);
   U150 : AOI22_X1 port map( A1 => ALU_output_20_port, A2 => n445, B1 => 
                           NPC2_20_port, B2 => n440, ZN => n171);
   U151 : AOI22_X1 port map( A1 => ALU_output_19_port, A2 => n446, B1 => 
                           NPC2_19_port, B2 => n440, ZN => n177);
   U152 : AOI22_X1 port map( A1 => ALU_output_17_port, A2 => n446, B1 => 
                           NPC2_17_port, B2 => n440, ZN => n183);
   U153 : AOI22_X1 port map( A1 => ALU_output_8_port, A2 => n441, B1 => 
                           NPC2_8_port, B2 => n440, ZN => n117);
   U154 : AOI22_X1 port map( A1 => ALU_output_6_port, A2 => n441, B1 => 
                           NPC2_6_port, B2 => JAL_op2, ZN => n123);
   U155 : AOI22_X1 port map( A1 => ALU_output_4_port, A2 => n442, B1 => 
                           NPC2_4_port, B2 => JAL_op2, ZN => n129);
   U156 : AOI22_X1 port map( A1 => ALU_output_2_port, A2 => n443, B1 => 
                           NPC2_2_port, B2 => JAL_op2, ZN => n141);
   U157 : AOI22_X1 port map( A1 => ALU_output_27_port, A2 => n444, B1 => 
                           NPC2_27_port, B2 => n440, ZN => n150);
   U158 : AOI22_X1 port map( A1 => ALU_output_25_port, A2 => n444, B1 => 
                           NPC2_25_port, B2 => n440, ZN => n156);
   U159 : AOI22_X1 port map( A1 => ALU_output_9_port, A2 => n441, B1 => 
                           NPC2_9_port, B2 => n440, ZN => n112);
   U160 : AOI22_X1 port map( A1 => ALU_output_7_port, A2 => n441, B1 => 
                           NPC2_7_port, B2 => JAL_op2, ZN => n120);
   U161 : AOI22_X1 port map( A1 => ALU_output_5_port, A2 => n442, B1 => 
                           NPC2_5_port, B2 => JAL_op2, ZN => n126);
   U162 : AOI22_X1 port map( A1 => ALU_output_3_port, A2 => n442, B1 => 
                           NPC2_3_port, B2 => JAL_op2, ZN => n132);
   U163 : AOI22_X1 port map( A1 => ALU_output_30_port, A2 => n443, B1 => 
                           NPC2_30_port, B2 => JAL_op2, ZN => n138);
   U164 : AOI22_X1 port map( A1 => ALU_output_29_port, A2 => n443, B1 => 
                           NPC2_29_port, B2 => JAL_op2, ZN => n144);
   U165 : AOI22_X1 port map( A1 => ALU_output_31_port, A2 => n442, B1 => 
                           NPC2_31_port, B2 => n440, ZN => n135);
   U166 : AND2_X1 port map( A1 => ALU_OPCODE(4), A2 => PC_enable1, ZN => 
                           ALU_OPCODE_in_0_port);
   U167 : NAND4_X1 port map( A1 => n280, A2 => n279, A3 => n229, A4 => n329, ZN
                           => n304);
   U168 : NOR3_X1 port map( A1 => Instr_reg_out_29_port, A2 => 
                           Instr_reg_out_31_port, A3 => Instr_reg_out_30_port, 
                           ZN => n329);
   U169 : OAI211_X1 port map( C1 => n218, C2 => n219, A => n107, B => n220, ZN 
                           => n104);
   U170 : INV_X1 port map( A => PC_enable, ZN => n219);
   U171 : NOR2_X1 port map( A1 => JR_op1, A2 => n108, ZN => n220);
   U172 : AOI22_X1 port map( A1 => LOAD_op1, A2 => n211, B1 => n109, B2 => 
                           FWD_B_mem_mem, ZN => n224);
   U173 : NAND4_X1 port map( A1 => n344, A2 => n345, A3 => n346, A4 => n347, ZN
                           => n230);
   U174 : XNOR2_X1 port map( A => Instr_reg_out_23_port, B => RD1_2_port, ZN =>
                           n344);
   U175 : XNOR2_X1 port map( A => Instr_reg_out_24_port, B => RD1_3_port, ZN =>
                           n346);
   U176 : XNOR2_X1 port map( A => Instr_reg_out_25_port, B => RD1_4_port, ZN =>
                           n345);
   U177 : NOR2_X1 port map( A1 => SPILL, A2 => FILL, ZN => PC_enable);
   U178 : XNOR2_X1 port map( A => Instr_reg_out_25_port, B => RD2_4_port, ZN =>
                           n337);
   U179 : NOR3_X1 port map( A1 => n289, A2 => n290, A3 => n291, ZN => n286);
   U180 : XNOR2_X1 port map( A => RD2_2_port, B => n215, ZN => n289);
   U181 : XNOR2_X1 port map( A => RD2_3_port, B => n214, ZN => n291);
   U182 : NOR3_X1 port map( A1 => n319, A2 => n320, A3 => n321, ZN => n316);
   U183 : XNOR2_X1 port map( A => RD1_4_port, B => n213, ZN => n319);
   U184 : XNOR2_X1 port map( A => RD1_3_port, B => n214, ZN => n321);
   U185 : NOR3_X1 port map( A1 => n292, A2 => n293, A3 => n294, ZN => n285);
   U186 : XNOR2_X1 port map( A => RD2_1_port, B => n216, ZN => n292);
   U187 : XNOR2_X1 port map( A => RD2_0_port, B => n217, ZN => n293);
   U188 : XNOR2_X1 port map( A => RD2_4_port, B => n213, ZN => n294);
   U189 : XNOR2_X1 port map( A => Instr_reg_out_20_port, B => RD1_4_port, ZN =>
                           n307);
   U190 : XNOR2_X1 port map( A => Instr_reg_out_19_port, B => RD1_3_port, ZN =>
                           n306);
   U191 : AOI211_X1 port map( C1 => Instr_reg_out_27_port, C2 => n229, A => 
                           Instr_reg_out_30_port, B => Instr_reg_out_28_port, 
                           ZN => n228);
   U192 : AND2_X1 port map( A1 => JR_op1, A2 => n211, ZN => n97);
   U193 : XNOR2_X1 port map( A => n231, B => EQ_COND, ZN => n226);
   U194 : NAND2_X1 port map( A1 => n237, A2 => n238, ZN => n236);
   U195 : NAND4_X1 port map( A1 => n241, A2 => n242, A3 => n243, A4 => n244, ZN
                           => n234);
   U196 : AND2_X1 port map( A1 => ALU_OPCODE(3), A2 => PC_enable1, ZN => 
                           ALU_OPCODE_in_1_port);
   U197 : NOR3_X1 port map( A1 => n323, A2 => n324, A3 => n325, ZN => n315);
   U198 : XNOR2_X1 port map( A => RD1_1_port, B => n216, ZN => n323);
   U199 : XNOR2_X1 port map( A => RD1_0_port, B => n217, ZN => n324);
   U200 : XNOR2_X1 port map( A => RD1_2_port, B => n215, ZN => n325);
   U201 : AND2_X1 port map( A1 => ALU_OPCODE(0), A2 => PC_enable1, ZN => 
                           ALU_OPCODE_in_4_port);
   U202 : AND2_X1 port map( A1 => ALU_OPCODE(1), A2 => PC_enable1, ZN => 
                           ALU_OPCODE_in_3_port);
   U203 : AOI21_X1 port map( B1 => n256, B2 => n257, A => FWD_wb_branch1, ZN =>
                           n232);
   U204 : AND4_X1 port map( A1 => n262, A2 => n263, A3 => n264, A4 => n265, ZN 
                           => n256);
   U205 : AND4_X1 port map( A1 => n258, A2 => n259, A3 => n260, A4 => n261, ZN 
                           => n257);
   U206 : NOR4_X1 port map( A1 => A_reg_out_12_port, A2 => A_reg_out_11_port, 
                           A3 => A_reg_out_10_port, A4 => A_reg_out_0_port, ZN 
                           => n262);
   U207 : NOR2_X1 port map( A1 => n348, A2 => n349, ZN => n347);
   U208 : AND2_X1 port map( A1 => n224, A2 => n225, ZN => n107);
   U209 : OR3_X1 port map( A1 => n226, A2 => forward_branch2, A3 => n227, ZN =>
                           n225);
   U210 : INV_X1 port map( A => BRANCH_op2, ZN => n227);
   U211 : OR4_X1 port map( A1 => ALU_WB_out_24_port, A2 => ALU_WB_out_25_port, 
                           A3 => ALU_WB_out_26_port, A4 => ALU_WB_out_27_port, 
                           ZN => n251);
   U212 : OR4_X1 port map( A1 => ALU_WB_out_0_port, A2 => ALU_WB_out_10_port, 
                           A3 => ALU_WB_out_11_port, A4 => ALU_WB_out_12_port, 
                           ZN => n255);
   U213 : OR4_X1 port map( A1 => ALU_WB_out_28_port, A2 => ALU_WB_out_29_port, 
                           A3 => ALU_WB_out_2_port, A4 => ALU_WB_out_30_port, 
                           ZN => n250);
   U214 : OR4_X1 port map( A1 => ALU_WB_out_13_port, A2 => ALU_WB_out_14_port, 
                           A3 => ALU_WB_out_15_port, A4 => ALU_WB_out_16_port, 
                           ZN => n254);
   U215 : OR4_X1 port map( A1 => ALU_WB_out_31_port, A2 => ALU_WB_out_3_port, 
                           A3 => ALU_WB_out_4_port, A4 => ALU_WB_out_5_port, ZN
                           => n249);
   U216 : OR4_X1 port map( A1 => ALU_WB_out_17_port, A2 => ALU_WB_out_18_port, 
                           A3 => ALU_WB_out_19_port, A4 => ALU_WB_out_1_port, 
                           ZN => n253);
   U217 : OR4_X1 port map( A1 => ALU_WB_out_6_port, A2 => ALU_WB_out_7_port, A3
                           => ALU_WB_out_8_port, A4 => ALU_WB_out_9_port, ZN =>
                           n248);
   U218 : OR4_X1 port map( A1 => ALU_WB_out_20_port, A2 => ALU_WB_out_21_port, 
                           A3 => ALU_WB_out_22_port, A4 => ALU_WB_out_23_port, 
                           ZN => n252);
   U219 : INV_X1 port map( A => Instr_reg_out_28_port, ZN => n279);
   U220 : NAND4_X1 port map( A1 => n125, A2 => n122, A3 => n239, A4 => n240, ZN
                           => n235);
   U221 : NOR3_X1 port map( A1 => ALU_reg_out_7_port, A2 => ALU_reg_out_9_port,
                           A3 => ALU_reg_out_8_port, ZN => n239);
   U222 : NOR4_X1 port map( A1 => ALU_reg_out_4_port, A2 => ALU_reg_out_3_port,
                           A3 => ALU_reg_out_31_port, A4 => ALU_reg_out_30_port
                           , ZN => n240);
   U223 : INV_X1 port map( A => JR_op1, ZN => n106);
   U224 : OAI221_X1 port map( B1 => n434, B2 => n173, C1 => n174, C2 => n432, A
                           => n175, ZN => RF_out_A_FWD_1_port);
   U225 : OAI221_X1 port map( B1 => n434, B2 => n206, C1 => n207, C2 => n432, A
                           => n208, ZN => RF_out_A_FWD_0_port);
   U226 : OAI221_X1 port map( B1 => n436, B2 => n122, C1 => n123, C2 => n433, A
                           => n124, ZN => RF_out_A_FWD_6_port);
   U227 : OAI221_X1 port map( B1 => n436, B2 => n128, C1 => n129, C2 => n433, A
                           => n130, ZN => RF_out_A_FWD_4_port);
   U228 : OAI221_X1 port map( B1 => n435, B2 => n140, C1 => n141, C2 => n433, A
                           => n142, ZN => RF_out_A_FWD_2_port);
   U229 : OAI221_X1 port map( B1 => n436, B2 => n119, C1 => n120, C2 => n433, A
                           => n121, ZN => RF_out_A_FWD_7_port);
   U230 : OAI221_X1 port map( B1 => n436, B2 => n125, C1 => n126, C2 => n433, A
                           => n127, ZN => RF_out_A_FWD_5_port);
   U231 : OAI221_X1 port map( B1 => n436, B2 => n131, C1 => n132, C2 => n433, A
                           => n133, ZN => RF_out_A_FWD_3_port);
   U232 : OAI221_X1 port map( B1 => n436, B2 => n134, C1 => n135, C2 => n433, A
                           => n136, ZN => RF_out_A_FWD_31_port);
   U233 : OAI221_X1 port map( B1 => n435, B2 => n167, C1 => n168, C2 => n433, A
                           => n169, ZN => RF_out_A_FWD_21_port);
   U234 : OAI221_X1 port map( B1 => n434, B2 => n179, C1 => n180, C2 => n432, A
                           => n181, ZN => RF_out_A_FWD_18_port);
   U235 : OAI221_X1 port map( B1 => n434, B2 => n185, C1 => n186, C2 => n432, A
                           => n187, ZN => RF_out_A_FWD_16_port);
   U236 : OAI221_X1 port map( B1 => n434, B2 => n188, C1 => n189, C2 => n432, A
                           => n190, ZN => RF_out_A_FWD_15_port);
   U237 : OAI221_X1 port map( B1 => n434, B2 => n191, C1 => n192, C2 => n432, A
                           => n193, ZN => RF_out_A_FWD_14_port);
   U238 : OAI221_X1 port map( B1 => n434, B2 => n194, C1 => n195, C2 => n432, A
                           => n196, ZN => RF_out_A_FWD_13_port);
   U239 : OAI221_X1 port map( B1 => n434, B2 => n197, C1 => n198, C2 => n432, A
                           => n199, ZN => RF_out_A_FWD_12_port);
   U240 : OAI221_X1 port map( B1 => n434, B2 => n200, C1 => n201, C2 => n432, A
                           => n202, ZN => RF_out_A_FWD_11_port);
   U241 : OAI221_X1 port map( B1 => n434, B2 => n203, C1 => n204, C2 => n432, A
                           => n205, ZN => RF_out_A_FWD_10_port);
   U242 : OAI221_X1 port map( B1 => n435, B2 => n164, C1 => n165, C2 => n433, A
                           => n166, ZN => RF_out_A_FWD_22_port);
   U243 : OAI221_X1 port map( B1 => n435, B2 => n170, C1 => n171, C2 => n433, A
                           => n172, ZN => RF_out_A_FWD_20_port);
   U244 : OAI221_X1 port map( B1 => n434, B2 => n176, C1 => n177, C2 => n432, A
                           => n178, ZN => RF_out_A_FWD_19_port);
   U245 : OAI221_X1 port map( B1 => n434, B2 => n182, C1 => n183, C2 => n432, A
                           => n184, ZN => RF_out_A_FWD_17_port);
   U246 : OAI221_X1 port map( B1 => n436, B2 => n116, C1 => n117, C2 => n433, A
                           => n118, ZN => RF_out_A_FWD_8_port);
   U247 : OAI221_X1 port map( B1 => n436, B2 => n111, C1 => n112, C2 => n433, A
                           => n114, ZN => RF_out_A_FWD_9_port);
   U248 : AND3_X1 port map( A1 => BRANCH_op2, A2 => n226, A3 => forward_branch2
                           , ZN => n218);
   U249 : NAND2_X1 port map( A1 => RF_out_A_8_port, A2 => n431, ZN => n118);
   U250 : NAND2_X1 port map( A1 => RF_out_A_6_port, A2 => n431, ZN => n124);
   U251 : NAND2_X1 port map( A1 => RF_out_A_4_port, A2 => n431, ZN => n130);
   U252 : NAND2_X1 port map( A1 => RF_out_A_9_port, A2 => n431, ZN => n114);
   U253 : NAND2_X1 port map( A1 => RF_out_A_7_port, A2 => n431, ZN => n121);
   U254 : NAND2_X1 port map( A1 => RF_out_A_5_port, A2 => n431, ZN => n127);
   U255 : NAND2_X1 port map( A1 => RF_out_A_3_port, A2 => n431, ZN => n133);
   U256 : NAND2_X1 port map( A1 => RF_out_A_31_port, A2 => n431, ZN => n136);
   U257 : NOR3_X1 port map( A1 => n98, A2 => n99, A3 => n100, ZN => n305);
   U258 : XOR2_X1 port map( A => Instr_reg_out_18_port, B => RD1_2_port, Z => 
                           n98);
   U259 : XOR2_X1 port map( A => Instr_reg_out_16_port, B => RD1_0_port, Z => 
                           n99);
   U260 : XOR2_X1 port map( A => Instr_reg_out_17_port, B => RD1_1_port, Z => 
                           n100);
   U261 : INV_X1 port map( A => Instr_reg_out_26_port, ZN => n229);
   U262 : INV_X1 port map( A => ALU_reg_out_0_port, ZN => n206);
   U263 : INV_X1 port map( A => ALU_reg_out_6_port, ZN => n122);
   U264 : INV_X1 port map( A => ALU_reg_out_10_port, ZN => n203);
   U265 : INV_X1 port map( A => ALU_reg_out_11_port, ZN => n200);
   U266 : INV_X1 port map( A => ALU_reg_out_5_port, ZN => n125);
   U267 : AND3_X1 port map( A1 => n282, A2 => n283, A3 => Instr(27), ZN => n281
                           );
   U268 : INV_X1 port map( A => Instr_reg_out_27_port, ZN => n280);
   U269 : AND4_X1 port map( A1 => LOAD_op1, A2 => n305, A3 => n306, A4 => n307,
                           ZN => FWD_B_mem_mem);
   U270 : AND2_X1 port map( A1 => n281, A2 => Instr(30), ZN => JR_op);
   U271 : INV_X1 port map( A => Instr_reg_out_31_port, ZN => n278);
   U272 : NAND2_X1 port map( A1 => RF_out_A_23_port, A2 => n430, ZN => n163);
   U273 : NAND2_X1 port map( A1 => RF_out_A_21_port, A2 => n430, ZN => n169);
   U274 : NAND2_X1 port map( A1 => RF_out_A_18_port, A2 => n429, ZN => n181);
   U275 : NAND2_X1 port map( A1 => RF_out_A_16_port, A2 => n429, ZN => n187);
   U276 : NAND2_X1 port map( A1 => RF_out_A_15_port, A2 => n429, ZN => n190);
   U277 : NAND2_X1 port map( A1 => RF_out_A_14_port, A2 => n429, ZN => n193);
   U278 : NAND2_X1 port map( A1 => RF_out_A_13_port, A2 => n429, ZN => n196);
   U279 : NAND2_X1 port map( A1 => RF_out_A_12_port, A2 => n429, ZN => n199);
   U280 : NAND2_X1 port map( A1 => RF_out_A_11_port, A2 => n429, ZN => n202);
   U281 : NAND2_X1 port map( A1 => RF_out_A_10_port, A2 => n429, ZN => n205);
   U282 : NAND2_X1 port map( A1 => RF_out_A_1_port, A2 => n429, ZN => n175);
   U283 : NAND2_X1 port map( A1 => RF_out_A_0_port, A2 => n429, ZN => n208);
   U284 : NAND2_X1 port map( A1 => RF_out_A_28_port, A2 => n430, ZN => n148);
   U285 : NAND2_X1 port map( A1 => RF_out_A_26_port, A2 => n430, ZN => n154);
   U286 : NAND2_X1 port map( A1 => RF_out_A_24_port, A2 => n430, ZN => n160);
   U287 : NAND2_X1 port map( A1 => RF_out_A_22_port, A2 => n430, ZN => n166);
   U288 : NAND2_X1 port map( A1 => RF_out_A_20_port, A2 => n430, ZN => n172);
   U289 : NAND2_X1 port map( A1 => RF_out_A_19_port, A2 => n429, ZN => n178);
   U290 : NAND2_X1 port map( A1 => RF_out_A_17_port, A2 => n429, ZN => n184);
   U291 : NAND2_X1 port map( A1 => RF_out_A_2_port, A2 => n430, ZN => n142);
   U292 : NAND2_X1 port map( A1 => RF_out_A_27_port, A2 => n430, ZN => n151);
   U293 : NAND2_X1 port map( A1 => RF_out_A_25_port, A2 => n430, ZN => n157);
   U294 : NAND2_X1 port map( A1 => RF_out_A_30_port, A2 => n430, ZN => n139);
   U295 : NAND2_X1 port map( A1 => RF_out_A_29_port, A2 => n430, ZN => n145);
   U296 : NOR4_X1 port map( A1 => n283, A2 => n422, A3 => Instr(27), A4 => 
                           Instr(30), ZN => BRANCH_op);
   U297 : INV_X1 port map( A => n282, ZN => n422);
   U298 : AND4_X1 port map( A1 => n200, A2 => n203, A3 => n206, A4 => 
                           FWD_exe_branch1, ZN => n241);
   U299 : INV_X1 port map( A => Instr(28), ZN => n283);
   U300 : AND4_X1 port map( A1 => n315, A2 => n316, A3 => n317, A4 => n318, ZN 
                           => FWD_B_exe_mem);
   U301 : NOR3_X1 port map( A1 => OPCODE1_0_port, A2 => OPCODE1_2_port, A3 => 
                           OPCODE1_1_port, ZN => n317);
   U302 : NOR3_X1 port map( A1 => OPCODE1_3_port, A2 => OPCODE1_5_port, A3 => 
                           OPCODE1_4_port, ZN => n318);
   U303 : AND4_X1 port map( A1 => n285, A2 => n286, A3 => n287, A4 => n288, ZN 
                           => FWD_B_wb_mem);
   U304 : NOR3_X1 port map( A1 => OPCODE2_0_port, A2 => OPCODE2_2_port, A3 => 
                           OPCODE2_1_port, ZN => n287);
   U305 : NOR3_X1 port map( A1 => OPCODE2_3_port, A2 => OPCODE2_5_port, A3 => 
                           OPCODE2_4_port, ZN => n288);
   U306 : NOR4_X1 port map( A1 => RD1_3_port, A2 => RD1_4_port, A3 => 
                           RD1_2_port, A4 => n343, ZN => n320);
   U307 : OR2_X1 port map( A1 => RD1_1_port, A2 => RD1_0_port, ZN => n343);
   U308 : NAND2_X1 port map( A1 => n266, A2 => n267, ZN => 
                           PC_Immediate_displacement_31_port);
   U309 : NAND2_X1 port map( A1 => JUMP_EN, A2 => Instr(25), ZN => n267);
   U310 : BUF_X2 port map( A => Rst, Z => n452);
   U311 : XNOR2_X1 port map( A => Instr_reg_out_20_port, B => RD2_4_port, ZN =>
                           n302);
   U312 : XNOR2_X1 port map( A => Instr_reg_out_19_port, B => RD2_3_port, ZN =>
                           n300);
   U313 : NAND4_X1 port map( A1 => LOAD_op2, A2 => n301, A3 => n300, A4 => n302
                           , ZN => n308);
   U314 : OR2_X1 port map( A1 => forward_branch, A2 => JUMP_EN, ZN => n266);
   U315 : OR2_X1 port map( A1 => PC_enable1, A2 => bootstrap, ZN => 
                           PC_enable_fixed);
   U316 : BUF_X1 port map( A => Rst, Z => n453);
   U317 : NOR3_X1 port map( A1 => n101, A2 => n102, A3 => n113, ZN => n301);
   U318 : XOR2_X1 port map( A => Instr_reg_out_18_port, B => RD2_2_port, Z => 
                           n101);
   U319 : XOR2_X1 port map( A => Instr_reg_out_16_port, B => RD2_0_port, Z => 
                           n102);
   U320 : XOR2_X1 port map( A => Instr_reg_out_17_port, B => RD2_1_port, Z => 
                           n113);
   U321 : OR3_X1 port map( A1 => STORE_op1, A2 => LOAD_op1, A3 => n320, ZN => 
                           n328);
   U322 : INV_X1 port map( A => BRANCH_op1, ZN => n284);
   U323 : INV_X1 port map( A => LOAD_op2, ZN => n335);
   U324 : INV_X1 port map( A => ALU_reg_out_9_port, ZN => n111);
   U325 : INV_X1 port map( A => ALU_reg_out_1_port, ZN => n173);
   U326 : INV_X1 port map( A => ALU_reg_out_8_port, ZN => n116);
   U327 : INV_X1 port map( A => ALU_reg_out_7_port, ZN => n119);
   U328 : INV_X1 port map( A => ALU_reg_out_3_port, ZN => n131);
   U329 : INV_X1 port map( A => ALU_reg_out_4_port, ZN => n128);
   U330 : INV_X1 port map( A => ALU_reg_out_2_port, ZN => n140);
   U331 : INV_X1 port map( A => ALU_reg_out_23_port, ZN => n161);
   U332 : INV_X1 port map( A => ALU_reg_out_16_port, ZN => n185);
   U333 : INV_X1 port map( A => ALU_reg_out_12_port, ZN => n197);
   U334 : INV_X1 port map( A => ALU_reg_out_27_port, ZN => n149);
   U335 : INV_X1 port map( A => ALU_reg_out_30_port, ZN => n137);
   U336 : INV_X1 port map( A => ALU_reg_out_13_port, ZN => n194);
   U337 : INV_X1 port map( A => ALU_reg_out_28_port, ZN => n146);
   U338 : INV_X1 port map( A => ALU_reg_out_24_port, ZN => n158);
   U339 : INV_X1 port map( A => ALU_reg_out_20_port, ZN => n170);
   U340 : INV_X1 port map( A => ALU_reg_out_17_port, ZN => n182);
   U341 : INV_X1 port map( A => ALU_reg_out_31_port, ZN => n134);
   U342 : INV_X1 port map( A => ALU_reg_out_21_port, ZN => n167);
   U343 : INV_X1 port map( A => ALU_reg_out_18_port, ZN => n179);
   U344 : INV_X1 port map( A => ALU_reg_out_14_port, ZN => n191);
   U345 : INV_X1 port map( A => ALU_reg_out_25_port, ZN => n155);
   U346 : INV_X1 port map( A => ALU_reg_out_29_port, ZN => n143);
   U347 : INV_X1 port map( A => ALU_reg_out_15_port, ZN => n188);
   U348 : INV_X1 port map( A => ALU_reg_out_26_port, ZN => n152);
   U349 : INV_X1 port map( A => ALU_reg_out_22_port, ZN => n164);
   U350 : INV_X1 port map( A => ALU_reg_out_19_port, ZN => n176);
   U351 : NAND2_X1 port map( A1 => n266, A2 => n268, ZN => 
                           PC_Immediate_displacement_24_port);
   U352 : NAND2_X1 port map( A1 => Instr(24), A2 => JUMP_EN, ZN => n268);
   U353 : NAND2_X1 port map( A1 => n266, A2 => n269, ZN => 
                           PC_Immediate_displacement_23_port);
   U354 : NAND2_X1 port map( A1 => Instr(23), A2 => JUMP_EN, ZN => n269);
   U355 : NAND2_X1 port map( A1 => n266, A2 => n270, ZN => 
                           PC_Immediate_displacement_22_port);
   U356 : NAND2_X1 port map( A1 => Instr(22), A2 => JUMP_EN, ZN => n270);
   U357 : NAND2_X1 port map( A1 => n266, A2 => n271, ZN => 
                           PC_Immediate_displacement_21_port);
   U358 : NAND2_X1 port map( A1 => Instr(21), A2 => JUMP_EN, ZN => n271);
   U359 : NAND2_X1 port map( A1 => n266, A2 => n272, ZN => 
                           PC_Immediate_displacement_20_port);
   U360 : NAND2_X1 port map( A1 => Instr(20), A2 => JUMP_EN, ZN => n272);
   U361 : NAND2_X1 port map( A1 => n266, A2 => n273, ZN => 
                           PC_Immediate_displacement_19_port);
   U362 : NAND2_X1 port map( A1 => Instr(19), A2 => JUMP_EN, ZN => n273);
   U363 : NAND2_X1 port map( A1 => n266, A2 => n274, ZN => 
                           PC_Immediate_displacement_18_port);
   U364 : NAND2_X1 port map( A1 => Instr(18), A2 => JUMP_EN, ZN => n274);
   U365 : NAND2_X1 port map( A1 => n266, A2 => n275, ZN => 
                           PC_Immediate_displacement_17_port);
   U366 : NAND2_X1 port map( A1 => Instr(17), A2 => JUMP_EN, ZN => n275);
   U367 : NAND2_X1 port map( A1 => n266, A2 => n276, ZN => 
                           PC_Immediate_displacement_16_port);
   U368 : NAND2_X1 port map( A1 => Instr(16), A2 => JUMP_EN, ZN => n276);
   U369 : INV_X1 port map( A => flush2_1_port, ZN => n298);
   U370 : INV_X1 port map( A => flush2_0_port, ZN => n297);
   U371 : INV_X1 port map( A => STORE_op2, ZN => n299);
   U372 : INV_X1 port map( A => Instr(15), ZN => forward_branch);
   U373 : OR2_X1 port map( A1 => RD2_1_port, A2 => RD2_0_port, ZN => n342);
   U374 : NOR4_X1 port map( A1 => Instr_reg_out_30_port, A2 => 
                           Instr_reg_out_29_port, A3 => n277, A4 => n278, ZN =>
                           LOAD_op);
   U375 : AOI21_X1 port map( B1 => Instr_reg_out_26_port, B2 => n279, A => n280
                           , ZN => n277);
   U376 : NOR4_X1 port map( A1 => JUMP_EN2, A2 => BRANCH_op1, A3 => n230, A4 =>
                           n328, ZN => FWD_A_exe_dec);
   U377 : NOR4_X1 port map( A1 => n333, A2 => n334, A3 => n290, A4 => n212, ZN 
                           => FWD_A_wb_dec);
   U378 : OR2_X1 port map( A1 => BRANCH_op1, A2 => JUMP_EN2, ZN => n334);
   U379 : NAND4_X1 port map( A1 => n335, A2 => n299, A3 => n297, A4 => n298, ZN
                           => n333);
   U380 : NOR3_X1 port map( A1 => n308, A2 => n290, A3 => n309, ZN => 
                           FWD_B_mem_exe);
   U381 : NOR4_X1 port map( A1 => Instr_reg_out_30_port, A2 => n310, A3 => n311
                           , A4 => n279, ZN => n309);
   U382 : INV_X1 port map( A => Instr_reg_out_29_port, ZN => n310);
   U383 : NOR4_X1 port map( A1 => n295, A2 => n296, A3 => LOAD_op2, A4 => n290,
                           ZN => FWD_B_wb_dec);
   U384 : NAND4_X1 port map( A1 => n300, A2 => n301, A3 => n302, A4 => n303, ZN
                           => n295);
   U385 : AND2_X1 port map( A1 => Instr(26), A2 => n281, ZN => JAL_op);
   U386 : NOR3_X1 port map( A1 => FWD_B_lmd1_mem2, A2 => FWD_B_mem_mem2, A3 => 
                           n418, ZN => n354);
   U387 : BUF_X1 port map( A => FWD_B_exe_mem2, Z => n439);
   U388 : NOR2_X1 port map( A1 => n421, A2 => n439, ZN => n352);
   U389 : INV_X1 port map( A => FWD_B_wb_mem2, ZN => n421);
   U390 : BUF_X1 port map( A => FWD_B_exe_mem2, Z => n438);
   U391 : BUF_X1 port map( A => FWD_B_exe_mem2, Z => n437);
   U392 : NOR2_X1 port map( A1 => n439, A2 => FWD_B_wb_mem2, ZN => n419);
   U393 : AND3_X1 port map( A1 => n419, A2 => n420, A3 => FWD_B_lmd1_mem2, ZN 
                           => n353);
   U394 : INV_X1 port map( A => FWD_B_mem_mem2, ZN => n420);
   U395 : NAND2_X1 port map( A1 => n366, A2 => n367, ZN => 
                           DRAM_write_data_FWD_3_port);
   U396 : AOI22_X1 port map( A1 => LMD_reg_out_3_port, A2 => n313, B1 => 
                           ALU_WB_out_3_port, B2 => n437, ZN => n366);
   U397 : AOI222_X1 port map( A1 => ALU_WB_out1_3_port, A2 => n428, B1 => 
                           LMD_reg_out1_3_port, B2 => n425, C1 => 
                           DRAM_write_data_3_port, C2 => n331, ZN => n367);
   U398 : NAND2_X1 port map( A1 => n364, A2 => n365, ZN => 
                           DRAM_write_data_FWD_4_port);
   U399 : AOI22_X1 port map( A1 => LMD_reg_out_4_port, A2 => n313, B1 => 
                           ALU_WB_out_4_port, B2 => n437, ZN => n364);
   U400 : AOI222_X1 port map( A1 => ALU_WB_out1_4_port, A2 => n428, B1 => 
                           LMD_reg_out1_4_port, B2 => n425, C1 => 
                           DRAM_write_data_4_port, C2 => n331, ZN => n365);
   U401 : NAND2_X1 port map( A1 => n362, A2 => n363, ZN => 
                           DRAM_write_data_FWD_5_port);
   U402 : AOI22_X1 port map( A1 => LMD_reg_out_5_port, A2 => n313, B1 => 
                           ALU_WB_out_5_port, B2 => n437, ZN => n362);
   U403 : AOI222_X1 port map( A1 => ALU_WB_out1_5_port, A2 => n428, B1 => 
                           LMD_reg_out1_5_port, B2 => n425, C1 => 
                           DRAM_write_data_5_port, C2 => n331, ZN => n363);
   U404 : NAND2_X1 port map( A1 => n360, A2 => n361, ZN => 
                           DRAM_write_data_FWD_6_port);
   U405 : AOI22_X1 port map( A1 => LMD_reg_out_6_port, A2 => n313, B1 => 
                           ALU_WB_out_6_port, B2 => n437, ZN => n360);
   U406 : AOI222_X1 port map( A1 => ALU_WB_out1_6_port, A2 => n428, B1 => 
                           LMD_reg_out1_6_port, B2 => n425, C1 => 
                           DRAM_write_data_6_port, C2 => n331, ZN => n361);
   U407 : NAND2_X1 port map( A1 => n358, A2 => n359, ZN => 
                           DRAM_write_data_FWD_7_port);
   U408 : AOI22_X1 port map( A1 => LMD_reg_out_7_port, A2 => n313, B1 => 
                           ALU_WB_out_7_port, B2 => n437, ZN => n358);
   U409 : AOI222_X1 port map( A1 => ALU_WB_out1_7_port, A2 => n428, B1 => 
                           LMD_reg_out1_7_port, B2 => n425, C1 => 
                           DRAM_write_data_7_port, C2 => n331, ZN => n359);
   U410 : NAND2_X1 port map( A1 => n356, A2 => n357, ZN => 
                           DRAM_write_data_FWD_8_port);
   U411 : AOI22_X1 port map( A1 => LMD_reg_out_8_port, A2 => n313, B1 => 
                           ALU_WB_out_8_port, B2 => n437, ZN => n356);
   U412 : AOI222_X1 port map( A1 => ALU_WB_out1_8_port, A2 => n428, B1 => 
                           LMD_reg_out1_8_port, B2 => n425, C1 => 
                           DRAM_write_data_8_port, C2 => n331, ZN => n357);
   U413 : NAND2_X1 port map( A1 => n350, A2 => n351, ZN => 
                           DRAM_write_data_FWD_9_port);
   U414 : AOI22_X1 port map( A1 => LMD_reg_out_9_port, A2 => n313, B1 => n439, 
                           B2 => ALU_WB_out_9_port, ZN => n350);
   U415 : AOI222_X1 port map( A1 => ALU_WB_out1_9_port, A2 => n428, B1 => 
                           LMD_reg_out1_9_port, B2 => n425, C1 => 
                           DRAM_write_data_9_port, C2 => n331, ZN => n351);
   U416 : NAND2_X1 port map( A1 => n368, A2 => n369, ZN => 
                           DRAM_write_data_FWD_31_port);
   U417 : AOI22_X1 port map( A1 => LMD_reg_out_31_port, A2 => n313, B1 => 
                           ALU_WB_out_31_port, B2 => n437, ZN => n368);
   U418 : AOI222_X1 port map( A1 => ALU_WB_out1_31_port, A2 => n428, B1 => 
                           LMD_reg_out1_31_port, B2 => n425, C1 => 
                           DRAM_write_data_31_port, C2 => n331, ZN => n369);
   U419 : NAND2_X1 port map( A1 => n416, A2 => n417, ZN => 
                           DRAM_write_data_FWD_0_port);
   U420 : AOI22_X1 port map( A1 => LMD_reg_out_0_port, A2 => n210, B1 => 
                           ALU_WB_out_0_port, B2 => n439, ZN => n416);
   U421 : AOI222_X1 port map( A1 => ALU_WB_out1_0_port, A2 => n426, B1 => 
                           LMD_reg_out1_0_port, B2 => n332, C1 => 
                           DRAM_write_data_0_port, C2 => n314, ZN => n417);
   U422 : NAND2_X1 port map( A1 => n394, A2 => n395, ZN => 
                           DRAM_write_data_FWD_1_port);
   U423 : AOI22_X1 port map( A1 => LMD_reg_out_1_port, A2 => n210, B1 => 
                           ALU_WB_out_1_port, B2 => n438, ZN => n394);
   U424 : AOI222_X1 port map( A1 => ALU_WB_out1_1_port, A2 => n426, B1 => 
                           LMD_reg_out1_1_port, B2 => n332, C1 => 
                           DRAM_write_data_1_port, C2 => n314, ZN => n395);
   U425 : NAND2_X1 port map( A1 => n372, A2 => n373, ZN => 
                           DRAM_write_data_FWD_2_port);
   U426 : AOI22_X1 port map( A1 => LMD_reg_out_2_port, A2 => n312, B1 => 
                           ALU_WB_out_2_port, B2 => n437, ZN => n372);
   U427 : AOI222_X1 port map( A1 => ALU_WB_out1_2_port, A2 => n427, B1 => 
                           LMD_reg_out1_2_port, B2 => n424, C1 => 
                           DRAM_write_data_2_port, C2 => n330, ZN => n373);
   U428 : NAND2_X1 port map( A1 => n414, A2 => n415, ZN => 
                           DRAM_write_data_FWD_10_port);
   U429 : AOI22_X1 port map( A1 => LMD_reg_out_10_port, A2 => n210, B1 => 
                           ALU_WB_out_10_port, B2 => n439, ZN => n414);
   U430 : AOI222_X1 port map( A1 => ALU_WB_out1_10_port, A2 => n426, B1 => 
                           LMD_reg_out1_10_port, B2 => n332, C1 => 
                           DRAM_write_data_10_port, C2 => n314, ZN => n415);
   U431 : NAND2_X1 port map( A1 => n412, A2 => n413, ZN => 
                           DRAM_write_data_FWD_11_port);
   U432 : AOI22_X1 port map( A1 => LMD_reg_out_11_port, A2 => n210, B1 => 
                           ALU_WB_out_11_port, B2 => n439, ZN => n412);
   U433 : AOI222_X1 port map( A1 => ALU_WB_out1_11_port, A2 => n426, B1 => 
                           LMD_reg_out1_11_port, B2 => n332, C1 => 
                           DRAM_write_data_11_port, C2 => n314, ZN => n413);
   U434 : NAND2_X1 port map( A1 => n410, A2 => n411, ZN => 
                           DRAM_write_data_FWD_12_port);
   U435 : AOI22_X1 port map( A1 => LMD_reg_out_12_port, A2 => n210, B1 => 
                           ALU_WB_out_12_port, B2 => n439, ZN => n410);
   U436 : AOI222_X1 port map( A1 => ALU_WB_out1_12_port, A2 => n426, B1 => 
                           LMD_reg_out1_12_port, B2 => n332, C1 => 
                           DRAM_write_data_12_port, C2 => n314, ZN => n411);
   U437 : NAND2_X1 port map( A1 => n408, A2 => n409, ZN => 
                           DRAM_write_data_FWD_13_port);
   U438 : AOI22_X1 port map( A1 => LMD_reg_out_13_port, A2 => n210, B1 => 
                           ALU_WB_out_13_port, B2 => n439, ZN => n408);
   U439 : AOI222_X1 port map( A1 => ALU_WB_out1_13_port, A2 => n426, B1 => 
                           LMD_reg_out1_13_port, B2 => n332, C1 => 
                           DRAM_write_data_13_port, C2 => n314, ZN => n409);
   U440 : NAND2_X1 port map( A1 => n406, A2 => n407, ZN => 
                           DRAM_write_data_FWD_14_port);
   U441 : AOI22_X1 port map( A1 => LMD_reg_out_14_port, A2 => n210, B1 => 
                           ALU_WB_out_14_port, B2 => n439, ZN => n406);
   U442 : AOI222_X1 port map( A1 => ALU_WB_out1_14_port, A2 => n426, B1 => 
                           LMD_reg_out1_14_port, B2 => n332, C1 => 
                           DRAM_write_data_14_port, C2 => n314, ZN => n407);
   U443 : NAND2_X1 port map( A1 => n404, A2 => n405, ZN => 
                           DRAM_write_data_FWD_15_port);
   U444 : AOI22_X1 port map( A1 => LMD_reg_out_15_port, A2 => n210, B1 => 
                           ALU_WB_out_15_port, B2 => n439, ZN => n404);
   U445 : AOI222_X1 port map( A1 => ALU_WB_out1_15_port, A2 => n426, B1 => 
                           LMD_reg_out1_15_port, B2 => n332, C1 => 
                           DRAM_write_data_15_port, C2 => n314, ZN => n405);
   U446 : NAND2_X1 port map( A1 => n402, A2 => n403, ZN => 
                           DRAM_write_data_FWD_16_port);
   U447 : AOI22_X1 port map( A1 => LMD_reg_out_16_port, A2 => n210, B1 => 
                           ALU_WB_out_16_port, B2 => n438, ZN => n402);
   U448 : AOI222_X1 port map( A1 => ALU_WB_out1_16_port, A2 => n426, B1 => 
                           LMD_reg_out1_16_port, B2 => n332, C1 => 
                           DRAM_write_data_16_port, C2 => n314, ZN => n403);
   U449 : NAND2_X1 port map( A1 => n400, A2 => n401, ZN => 
                           DRAM_write_data_FWD_17_port);
   U450 : AOI22_X1 port map( A1 => LMD_reg_out_17_port, A2 => n210, B1 => 
                           ALU_WB_out_17_port, B2 => n438, ZN => n400);
   U451 : AOI222_X1 port map( A1 => ALU_WB_out1_17_port, A2 => n426, B1 => 
                           LMD_reg_out1_17_port, B2 => n332, C1 => 
                           DRAM_write_data_17_port, C2 => n314, ZN => n401);
   U452 : NAND2_X1 port map( A1 => n398, A2 => n399, ZN => 
                           DRAM_write_data_FWD_18_port);
   U453 : AOI22_X1 port map( A1 => LMD_reg_out_18_port, A2 => n210, B1 => 
                           ALU_WB_out_18_port, B2 => n438, ZN => n398);
   U454 : AOI222_X1 port map( A1 => ALU_WB_out1_18_port, A2 => n426, B1 => 
                           LMD_reg_out1_18_port, B2 => n332, C1 => 
                           DRAM_write_data_18_port, C2 => n314, ZN => n399);
   U455 : NAND2_X1 port map( A1 => n396, A2 => n397, ZN => 
                           DRAM_write_data_FWD_19_port);
   U465 : AOI22_X1 port map( A1 => LMD_reg_out_19_port, A2 => n210, B1 => 
                           ALU_WB_out_19_port, B2 => n438, ZN => n396);
   U466 : AOI222_X1 port map( A1 => ALU_WB_out1_19_port, A2 => n426, B1 => 
                           LMD_reg_out1_19_port, B2 => n332, C1 => 
                           DRAM_write_data_19_port, C2 => n314, ZN => n397);
   U467 : NAND2_X1 port map( A1 => n392, A2 => n393, ZN => 
                           DRAM_write_data_FWD_20_port);
   U468 : AOI22_X1 port map( A1 => LMD_reg_out_20_port, A2 => n312, B1 => 
                           ALU_WB_out_20_port, B2 => n438, ZN => n392);
   U469 : AOI222_X1 port map( A1 => ALU_WB_out1_20_port, A2 => n427, B1 => 
                           LMD_reg_out1_20_port, B2 => n424, C1 => 
                           DRAM_write_data_20_port, C2 => n330, ZN => n393);
   U470 : NAND2_X1 port map( A1 => n390, A2 => n391, ZN => 
                           DRAM_write_data_FWD_21_port);
   U471 : AOI22_X1 port map( A1 => LMD_reg_out_21_port, A2 => n312, B1 => 
                           ALU_WB_out_21_port, B2 => n438, ZN => n390);
   U472 : AOI222_X1 port map( A1 => ALU_WB_out1_21_port, A2 => n427, B1 => 
                           LMD_reg_out1_21_port, B2 => n424, C1 => 
                           DRAM_write_data_21_port, C2 => n330, ZN => n391);
   U473 : NAND2_X1 port map( A1 => n388, A2 => n389, ZN => 
                           DRAM_write_data_FWD_22_port);
   U474 : AOI22_X1 port map( A1 => LMD_reg_out_22_port, A2 => n312, B1 => 
                           ALU_WB_out_22_port, B2 => n438, ZN => n388);
   U475 : AOI222_X1 port map( A1 => ALU_WB_out1_22_port, A2 => n427, B1 => 
                           LMD_reg_out1_22_port, B2 => n424, C1 => 
                           DRAM_write_data_22_port, C2 => n330, ZN => n389);
   U476 : NAND2_X1 port map( A1 => n386, A2 => n387, ZN => 
                           DRAM_write_data_FWD_23_port);
   U477 : AOI22_X1 port map( A1 => LMD_reg_out_23_port, A2 => n312, B1 => 
                           ALU_WB_out_23_port, B2 => n438, ZN => n386);
   U478 : AOI222_X1 port map( A1 => ALU_WB_out1_23_port, A2 => n427, B1 => 
                           LMD_reg_out1_23_port, B2 => n424, C1 => 
                           DRAM_write_data_23_port, C2 => n330, ZN => n387);
   U479 : NAND2_X1 port map( A1 => n384, A2 => n385, ZN => 
                           DRAM_write_data_FWD_24_port);
   U480 : AOI22_X1 port map( A1 => LMD_reg_out_24_port, A2 => n312, B1 => 
                           ALU_WB_out_24_port, B2 => n438, ZN => n384);
   U481 : AOI222_X1 port map( A1 => ALU_WB_out1_24_port, A2 => n427, B1 => 
                           LMD_reg_out1_24_port, B2 => n424, C1 => 
                           DRAM_write_data_24_port, C2 => n330, ZN => n385);
   U482 : NAND2_X1 port map( A1 => n382, A2 => n383, ZN => 
                           DRAM_write_data_FWD_25_port);
   U483 : AOI22_X1 port map( A1 => LMD_reg_out_25_port, A2 => n312, B1 => 
                           ALU_WB_out_25_port, B2 => n438, ZN => n382);
   U484 : AOI222_X1 port map( A1 => ALU_WB_out1_25_port, A2 => n427, B1 => 
                           LMD_reg_out1_25_port, B2 => n424, C1 => 
                           DRAM_write_data_25_port, C2 => n330, ZN => n383);
   U485 : NAND2_X1 port map( A1 => n380, A2 => n381, ZN => 
                           DRAM_write_data_FWD_26_port);
   U486 : AOI22_X1 port map( A1 => LMD_reg_out_26_port, A2 => n312, B1 => 
                           ALU_WB_out_26_port, B2 => n437, ZN => n380);
   U487 : AOI222_X1 port map( A1 => ALU_WB_out1_26_port, A2 => n427, B1 => 
                           LMD_reg_out1_26_port, B2 => n424, C1 => 
                           DRAM_write_data_26_port, C2 => n330, ZN => n381);
   U488 : NAND2_X1 port map( A1 => n378, A2 => n379, ZN => 
                           DRAM_write_data_FWD_27_port);
   U489 : AOI22_X1 port map( A1 => LMD_reg_out_27_port, A2 => n312, B1 => 
                           ALU_WB_out_27_port, B2 => n437, ZN => n378);
   U490 : AOI222_X1 port map( A1 => ALU_WB_out1_27_port, A2 => n427, B1 => 
                           LMD_reg_out1_27_port, B2 => n424, C1 => 
                           DRAM_write_data_27_port, C2 => n330, ZN => n379);
   U491 : NAND2_X1 port map( A1 => n376, A2 => n377, ZN => 
                           DRAM_write_data_FWD_28_port);
   U492 : AOI22_X1 port map( A1 => LMD_reg_out_28_port, A2 => n312, B1 => 
                           ALU_WB_out_28_port, B2 => n437, ZN => n376);
   U493 : AOI222_X1 port map( A1 => ALU_WB_out1_28_port, A2 => n427, B1 => 
                           LMD_reg_out1_28_port, B2 => n424, C1 => 
                           DRAM_write_data_28_port, C2 => n330, ZN => n377);
   U494 : NAND2_X1 port map( A1 => n374, A2 => n375, ZN => 
                           DRAM_write_data_FWD_29_port);
   U495 : AOI22_X1 port map( A1 => LMD_reg_out_29_port, A2 => n312, B1 => 
                           ALU_WB_out_29_port, B2 => n437, ZN => n374);
   U496 : AOI222_X1 port map( A1 => ALU_WB_out1_29_port, A2 => n427, B1 => 
                           LMD_reg_out1_29_port, B2 => n424, C1 => 
                           DRAM_write_data_29_port, C2 => n330, ZN => n375);
   U497 : NAND2_X1 port map( A1 => n370, A2 => n371, ZN => 
                           DRAM_write_data_FWD_30_port);
   U498 : AOI22_X1 port map( A1 => LMD_reg_out_30_port, A2 => n312, B1 => 
                           ALU_WB_out_30_port, B2 => n438, ZN => n370);
   U499 : AOI222_X1 port map( A1 => ALU_WB_out1_30_port, A2 => n427, B1 => 
                           LMD_reg_out1_30_port, B2 => n424, C1 => 
                           DRAM_write_data_30_port, C2 => n330, ZN => n371);
   n454 <= '1';

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dlx.all;

entity dlx is

   port( Clk, Rst : in std_logic;  IR : in bus32;  PC : out bus32);

end dlx;

architecture SYN_struct of dlx is

   component CU_HW
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  flush : in std_logic_vector (1 downto 0);  JUMP_EN, RF_RD1_EN, 
            RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, MUXA_SEL, MUXB_SEL, EQ_COND :
            out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 4);  
            SEL_STORE1, SEL_STORE0, SEL_LOAD2, SEL_LOAD1, SEL_LOAD0, DRAM_WR, 
            WB_MUX_SEL, RF_WR : out std_logic);
   end component;
   
   component datapath
      port( Clk, Rst : in std_logic;  Instr : in std_logic_vector (31 downto 0)
            ;  JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, 
            MUXA_SEL, MUXB_SEL, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 4);  SEL_STORE1, SEL_STORE0, SEL_LOAD2, 
            SEL_LOAD1, SEL_LOAD0, DRAM_WR, WB_MUX_SEL, RF_WR : in std_logic;  
            flush : out std_logic_vector (1 downto 0);  PC_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, MUXA_SEL, 
      MUXB_SEL, EQ_COND, ALU_OPCODE_4_port, ALU_OPCODE_3_port, 
      ALU_OPCODE_2_port, ALU_OPCODE_1_port, ALU_OPCODE_0_port, SEL_STORE1, 
      SEL_STORE0, SEL_LOAD2, SEL_LOAD1, SEL_LOAD0, DRAM_WR, WB_MUX_SEL, RF_WR, 
      flush_1_port, flush_0_port, net271204, net271205, net271206, net271207, 
      net271208, net271209, net271210, net271211, net271212, net271213, 
      net271214, net271215, net271216, net271217, net271218, net271219, 
      net271220, net271221, net271222, net271223, net271224, net271225, 
      net271226 : std_logic;

begin
   
   RF_WR <= '0';
   WB_MUX_SEL <= '0';
   DRAM_WR <= '0';
   SEL_LOAD0 <= '0';
   SEL_LOAD1 <= '0';
   SEL_LOAD2 <= '0';
   SEL_STORE0 <= '0';
   SEL_STORE1 <= '0';
   ALU_OPCODE_0_port <= '0';
   ALU_OPCODE_1_port <= '0';
   ALU_OPCODE_2_port <= '0';
   ALU_OPCODE_3_port <= '0';
   ALU_OPCODE_4_port <= '0';
   EQ_COND <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   IMM_SEL <= '0';
   RET <= '0';
   CALL <= '0';
   RF_EN <= '0';
   RF_RD2_EN <= '0';
   RF_RD1_EN <= '0';
   JUMP_EN <= '0';
   DTP : datapath port map( Clk => Clk, Rst => Rst, Instr(31) => IR(31), 
                           Instr(30) => IR(30), Instr(29) => IR(29), Instr(28) 
                           => IR(28), Instr(27) => IR(27), Instr(26) => IR(26),
                           Instr(25) => IR(25), Instr(24) => IR(24), Instr(23) 
                           => IR(23), Instr(22) => IR(22), Instr(21) => IR(21),
                           Instr(20) => IR(20), Instr(19) => IR(19), Instr(18) 
                           => IR(18), Instr(17) => IR(17), Instr(16) => IR(16),
                           Instr(15) => IR(15), Instr(14) => IR(14), Instr(13) 
                           => IR(13), Instr(12) => IR(12), Instr(11) => IR(11),
                           Instr(10) => IR(10), Instr(9) => IR(9), Instr(8) => 
                           IR(8), Instr(7) => IR(7), Instr(6) => IR(6), 
                           Instr(5) => IR(5), Instr(4) => IR(4), Instr(3) => 
                           IR(3), Instr(2) => IR(2), Instr(1) => IR(1), 
                           Instr(0) => IR(0), JUMP_EN => JUMP_EN, RF_RD1_EN => 
                           RF_RD1_EN, RF_RD2_EN => RF_RD2_EN, RF_EN => RF_EN, 
                           CALL => CALL, RET => RET, IMM_SEL => IMM_SEL, 
                           MUXA_SEL => MUXA_SEL, MUXB_SEL => MUXB_SEL, EQ_COND 
                           => EQ_COND, ALU_OPCODE(0) => ALU_OPCODE_4_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_3_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_0_port, SEL_STORE1 => SEL_STORE1, 
                           SEL_STORE0 => SEL_STORE0, SEL_LOAD2 => SEL_LOAD2, 
                           SEL_LOAD1 => SEL_LOAD1, SEL_LOAD0 => SEL_LOAD0, 
                           DRAM_WR => DRAM_WR, WB_MUX_SEL => WB_MUX_SEL, RF_WR 
                           => RF_WR, flush(1) => flush_1_port, flush(0) => 
                           flush_0_port, PC_out(31) => PC(31), PC_out(30) => 
                           PC(30), PC_out(29) => PC(29), PC_out(28) => PC(28), 
                           PC_out(27) => PC(27), PC_out(26) => PC(26), 
                           PC_out(25) => PC(25), PC_out(24) => PC(24), 
                           PC_out(23) => PC(23), PC_out(22) => PC(22), 
                           PC_out(21) => PC(21), PC_out(20) => PC(20), 
                           PC_out(19) => PC(19), PC_out(18) => PC(18), 
                           PC_out(17) => PC(17), PC_out(16) => PC(16), 
                           PC_out(15) => PC(15), PC_out(14) => PC(14), 
                           PC_out(13) => PC(13), PC_out(12) => PC(12), 
                           PC_out(11) => PC(11), PC_out(10) => PC(10), 
                           PC_out(9) => PC(9), PC_out(8) => PC(8), PC_out(7) =>
                           PC(7), PC_out(6) => PC(6), PC_out(5) => PC(5), 
                           PC_out(4) => PC(4), PC_out(3) => PC(3), PC_out(2) =>
                           PC(2), PC_out(1) => PC(1), PC_out(0) => PC(0));
   CTRLU : CU_HW port map( Clk => Clk, Rst => Rst, IR_IN(31) => IR(31), 
                           IR_IN(30) => IR(30), IR_IN(29) => IR(29), IR_IN(28) 
                           => IR(28), IR_IN(27) => IR(27), IR_IN(26) => IR(26),
                           IR_IN(25) => IR(25), IR_IN(24) => IR(24), IR_IN(23) 
                           => IR(23), IR_IN(22) => IR(22), IR_IN(21) => IR(21),
                           IR_IN(20) => IR(20), IR_IN(19) => IR(19), IR_IN(18) 
                           => IR(18), IR_IN(17) => IR(17), IR_IN(16) => IR(16),
                           IR_IN(15) => IR(15), IR_IN(14) => IR(14), IR_IN(13) 
                           => IR(13), IR_IN(12) => IR(12), IR_IN(11) => IR(11),
                           IR_IN(10) => IR(10), IR_IN(9) => IR(9), IR_IN(8) => 
                           IR(8), IR_IN(7) => IR(7), IR_IN(6) => IR(6), 
                           IR_IN(5) => IR(5), IR_IN(4) => IR(4), IR_IN(3) => 
                           IR(3), IR_IN(2) => IR(2), IR_IN(1) => IR(1), 
                           IR_IN(0) => IR(0), flush(1) => flush_1_port, 
                           flush(0) => flush_0_port, JUMP_EN => net271204, 
                           RF_RD1_EN => net271205, RF_RD2_EN => net271206, 
                           RF_EN => net271207, CALL => net271208, RET => 
                           net271209, IMM_SEL => net271210, MUXA_SEL => 
                           net271211, MUXB_SEL => net271212, EQ_COND => 
                           net271213, ALU_OPCODE(0) => net271214, ALU_OPCODE(1)
                           => net271215, ALU_OPCODE(2) => net271216, 
                           ALU_OPCODE(3) => net271217, ALU_OPCODE(4) => 
                           net271218, SEL_STORE1 => net271219, SEL_STORE0 => 
                           net271220, SEL_LOAD2 => net271221, SEL_LOAD1 => 
                           net271222, SEL_LOAD0 => net271223, DRAM_WR => 
                           net271224, WB_MUX_SEL => net271225, RF_WR => 
                           net271226);

end SYN_struct;
