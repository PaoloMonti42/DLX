
module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_217 UIV ( .A(S), .Y(SB) );
  ND2_663 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_662 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_661 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_216 UIV ( .A(S), .Y(SB) );
  ND2_660 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_659 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_658 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_215 UIV ( .A(S), .Y(SB) );
  ND2_657 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_656 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_655 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_214 UIV ( .A(S), .Y(SB) );
  ND2_654 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_653 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_652 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_213 UIV ( .A(S), .Y(SB) );
  ND2_651 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_650 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_649 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_212 UIV ( .A(S), .Y(SB) );
  ND2_648 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_647 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_646 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_211 UIV ( .A(S), .Y(SB) );
  ND2_645 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_644 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_643 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_210 UIV ( .A(S), .Y(SB) );
  ND2_642 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_641 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_640 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_209 UIV ( .A(S), .Y(SB) );
  ND2_639 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_638 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_637 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_208 UIV ( .A(S), .Y(SB) );
  ND2_636 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_635 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_634 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_207 UIV ( .A(S), .Y(SB) );
  ND2_633 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_632 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_631 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_206 UIV ( .A(S), .Y(SB) );
  ND2_630 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_629 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_628 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_205 UIV ( .A(S), .Y(SB) );
  ND2_627 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_626 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_625 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_204 UIV ( .A(S), .Y(SB) );
  ND2_624 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_623 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_622 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_203 UIV ( .A(S), .Y(SB) );
  ND2_621 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_620 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_619 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_202 UIV ( .A(S), .Y(SB) );
  ND2_618 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_617 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_616 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_201 UIV ( .A(S), .Y(SB) );
  ND2_615 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_614 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_613 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_200 UIV ( .A(S), .Y(SB) );
  ND2_612 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_611 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_610 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_199 UIV ( .A(S), .Y(SB) );
  ND2_609 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_608 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_607 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_198 UIV ( .A(S), .Y(SB) );
  ND2_606 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_605 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_604 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_197 UIV ( .A(S), .Y(SB) );
  ND2_603 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_602 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_601 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_196 UIV ( .A(S), .Y(SB) );
  ND2_600 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_599 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_598 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_195 UIV ( .A(S), .Y(SB) );
  ND2_597 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_596 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_595 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_194 UIV ( .A(S), .Y(SB) );
  ND2_594 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_593 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_592 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_193 UIV ( .A(S), .Y(SB) );
  ND2_591 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_590 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_589 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_192 UIV ( .A(S), .Y(SB) );
  ND2_588 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_587 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_586 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_585 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_584 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_583 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_582 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_581 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_580 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_579 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_578 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_577 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_576 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module reg_N2_1 ( clk, rst, d_in, d_out );
  input [1:0] d_in;
  output [1:0] d_out;
  input clk, rst;
  wire   N2, N3;

  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in[1]), .ZN(N3) );
  AND2_X1 U4 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
endmodule


module ff_31 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_30 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_29 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_28 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_27 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_26 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_25 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_24 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_23 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_22 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_21 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_20 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_19 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_18 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_17 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_16 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_15 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_14 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_13 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_12 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_11 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_10 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_9 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_8 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_7 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_6 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_5 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_4 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_3 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_2 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module ff_1 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module MUX21_GENERIC_N32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_186 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_185 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_184 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_183 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_182 M_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_181 M_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_180 M_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_179 M_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_178 M_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_177 M_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_176 M_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_175 M_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_174 M_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_173 M_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_172 M_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_171 M_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_170 M_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_169 M_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_168 M_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_167 M_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_166 M_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_165 M_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_164 M_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_163 M_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_162 M_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_161 M_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_160 M_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_159 M_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_158 M_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_157 M_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_156 M_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_155 M_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module MUX21_GENERIC_N32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_154 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_153 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_152 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_151 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_150 M_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_149 M_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_148 M_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_147 M_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_146 M_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_145 M_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_144 M_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_143 M_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_142 M_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_141 M_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_140 M_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_139 M_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_138 M_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_137 M_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_136 M_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_135 M_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_134 M_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_133 M_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_132 M_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_131 M_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_130 M_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_129 M_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_128 M_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_127 M_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_126 M_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_125 M_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_124 M_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_123 M_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module MUX21_GENERIC_N32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_122 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_121 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_120 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_119 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_118 M_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_117 M_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_116 M_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_115 M_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_114 M_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_113 M_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_112 M_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_111 M_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_110 M_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_109 M_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_108 M_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_107 M_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_106 M_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_105 M_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_104 M_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_103 M_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_102 M_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_101 M_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_100 M_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_99 M_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_98 M_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_97 M_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_96 M_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_95 M_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_94 M_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_93 M_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_92 M_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_91 M_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module reg_N32_7 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U9 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U10 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U11 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U12 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U13 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U14 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U15 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U16 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U17 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U18 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U19 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U20 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U21 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U22 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U23 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U24 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U25 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U26 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U27 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U28 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U29 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U30 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U31 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U32 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U33 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U34 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U35 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U36 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  AND2_X1 U37 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
endmodule


module reg_N32_2 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U9 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U10 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U11 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U12 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U13 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U14 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U15 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U16 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U17 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U18 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U19 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U20 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U21 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U22 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U23 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U24 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U25 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U26 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U27 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U28 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U29 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U30 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U31 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U32 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U33 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U34 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U35 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U36 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  AND2_X1 U37 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
endmodule


module reg_N32_12 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module reg_N32_11 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module reg_N32_9 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module reg_N32_8 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module reg_N32_3 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module reg_N32_1 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_30_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_31_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_94_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_0_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_0_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_30_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_31_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_94_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_0_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_0_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n18), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n18) );
  INV_X1 U1 ( .A(n17), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n18), .B2(Ci), .ZN(n17) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_30_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30_1 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_31_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31_1 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_0_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0_1 UIV ( .A(S), .Y(SB) );
  ND2_0_1 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95_1 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_62_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_63_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_0_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n8), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U1 ( .A(n7), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_98 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_97 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_96 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_101 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_100 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_99 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_104 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_103 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_102 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_107 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_106 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_105 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_110 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_109 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_108 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_113 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_112 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_111 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_116 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_115 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_114 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_119 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_118 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_117 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_122 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_121 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_120 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_125 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_124 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_123 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_128 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_127 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_126 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_131 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_130 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_129 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_134 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_133 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_132 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_137 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_136 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_135 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_140 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_139 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_138 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_143 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_142 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_141 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_146 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_145 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_144 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_149 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_148 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_147 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_152 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_151 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_150 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_155 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_154 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_153 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_158 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_157 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_156 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_161 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_160 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_159 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_164 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_163 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_162 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_167 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_166 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_165 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_170 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_169 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_168 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_173 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_172 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_171 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_176 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_175 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_174 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_179 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_178 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_177 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_182 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_181 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_180 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_30_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30_0 UIV ( .A(S), .Y(SB) );
  ND2_185 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_184 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_183 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_31_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31_0 UIV ( .A(S), .Y(SB) );
  ND2_188 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_187 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_186 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_0_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0_0 UIV ( .A(S), .Y(SB) );
  ND2_0_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95_0 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94_0 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_62_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_0_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module ND2 ( A, B, Y );
  input A, B;
  output Y;
  wire   N0;

  GTECH_NOT I_0 ( .A(N0), .Z(Y) );
  GTECH_AND2 C7 ( .A(A), .B(B), .Z(N0) );
endmodule


module IV ( A, Y );
  input A;
  output Y;


  GTECH_NOT I_0 ( .A(A), .Z(Y) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_6_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_7_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_14_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_0_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_0_1 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31_1 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30_1 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_15_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_0_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0_1 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63_1 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62_1 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_8 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_35 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_34 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_33 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_32 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_259 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_258 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_257 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_256 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_263 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_262 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_261 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_260 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_9 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_39 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_38 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_37 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_36 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_267 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_266 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_265 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_264 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_271 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_270 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_269 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_268 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_10 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_43 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_42 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_41 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_40 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_275 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_274 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_273 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_272 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_279 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_278 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_277 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_276 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_11 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_47 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_46 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_45 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_44 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_283 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_282 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_281 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_280 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_287 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_286 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_285 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_284 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_12 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_51 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_50 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_49 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_48 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_291 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_290 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_289 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_288 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_295 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_294 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_293 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_292 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_6_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_55 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_54 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_53 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_52 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_299 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_298 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_297 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_296 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_303 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_302 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_301 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_300 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_7_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_59 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_58 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_57 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_56 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_307 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_306 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_305 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_304 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_14_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_311 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_310 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_309 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_308 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_0_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_0_0 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31_0 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30_0 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_60 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4_15_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_315 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_314 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_313 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_312 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module rca_generic_N4_0_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63_0 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62_0 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_316 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV UIV ( .A(S), .Y(SB) );
  ND2 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   N0, N1, N2, N3, N4;

  GTECH_XOR2 C7 ( .A(N0), .B(Ci), .Z(S) );
  GTECH_XOR2 C8 ( .A(A), .B(B), .Z(N0) );
  GTECH_OR2 C9 ( .A(N3), .B(N4), .Z(Co) );
  GTECH_OR2 C10 ( .A(N1), .B(N2), .Z(N3) );
  GTECH_AND2 C11 ( .A(A), .B(B), .Z(N1) );
  GTECH_AND2 C12 ( .A(B), .B(Ci), .Z(N2) );
  GTECH_AND2 C13 ( .A(A), .B(Ci), .Z(N4) );
endmodule


module carry_select_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_1 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_2 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_3 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_4 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_5 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_6_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_6_1 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module carry_select_N4_7_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_14_1 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_7_1 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module carry_select_N4_0_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_0_1 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_15_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_0_1 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module G_3 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module G_4 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n8) );
endmodule


module G_7 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module G_9 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module PG_2 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module G_5_1 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n8) );
endmodule


module G_6_1 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n6) );
endmodule


module PG_3 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_4_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n6) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_13 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module G_1 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n11;

  INV_X1 U1 ( .A(n11), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n11) );
endmodule


module PG_5 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_6 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n9;

  INV_X1 U1 ( .A(n9), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n9) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_14 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_15 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_16 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n10) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_17 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n10) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_19 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  AOI21_X1 U1 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  INV_X1 U2 ( .A(n8), .ZN(gout) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module G_8_1 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n6) );
endmodule


module PG_7 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_8 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_9 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_10 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_20 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n9;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n9), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n9) );
endmodule


module PG_18_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n8), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module PG_11 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_23 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_21_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_22_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_12 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_24_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n6) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_25_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n9;

  INV_X1 U1 ( .A(n9), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n9) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_26_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_0_1 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module G_2 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n8) );
endmodule


module PGnet_block_1 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_2 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_3 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_4 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_5 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_6 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_7 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_8 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_9 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_10 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_11 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_12 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_13 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_14 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_15 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_16 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_17 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_18 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_19 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_20 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_21 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_22 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_23 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_24 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_25 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_26 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_27 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_28 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_29 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_30_1 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_31_1 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module G_0_1 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module PGnet_block_0_1 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module carry_select_N4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_17 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_16 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_8 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_19 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_18 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_9 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_21 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_20 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_10 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_23 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_22 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_11 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_25 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_24 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_12 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module carry_select_N4_6_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_27 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_26 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_6_0 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module carry_select_N4_7_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_14_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_28 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_7_0 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module carry_select_N4_0_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4_0_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4_15_0 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4_0_0 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S)
         );
endmodule


module G_10 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module G_11 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n8) );
endmodule


module G_12 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n7) );
endmodule


module G_13 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module PG_27 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
endmodule


module PG_28 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module G_5_0 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module G_6_0 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module PG_29 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_4_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_30 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module G_14 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module PG_31 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  AOI21_X1 U1 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_32 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n9;

  INV_X1 U1 ( .A(n9), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n9) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_33 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_34 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_35 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n10) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_36 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_37 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(gout) );
  AND2_X1 U2 ( .A1(pright), .A2(pleft), .ZN(pout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n8) );
endmodule


module G_8_0 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module PG_38 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_39 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_40 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_41 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_42 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n2), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
endmodule


module PG_18_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n2), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
endmodule


module PG_43 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n7) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_44 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_21_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  AND2_X1 U1 ( .A1(pright), .A2(pleft), .ZN(pout) );
  INV_X1 U2 ( .A(n2), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
endmodule


module PG_22_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_45 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_24_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_25_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_26_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module PG_0_0 ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gright), .B2(pleft), .A(gleft), .ZN(n2) );
  AND2_X1 U3 ( .A1(pright), .A2(pleft), .ZN(pout) );
endmodule


module G_15 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
endmodule


module PGnet_block_32 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_33 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_34 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_35 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_36 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_37 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_38 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_39 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_40 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_41 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_42 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_43 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_44 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_45 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_46 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_47 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_48 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_49 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_50 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_51 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_52 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_53 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_54 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_55 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_56 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_57 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_58 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_59 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_60 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_30_0 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module PGnet_block_31_0 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module G_0_0 ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   n2;

  AOI21_X1 U1 ( .B1(pleft), .B2(gright), .A(gleft), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(gout) );
endmodule


module PGnet_block_0_0 ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(pout) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(gout) );
endmodule


module MUX21_GENERIC_N4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module rca_generic_N4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module sum_generator_Nbits32_Nblocks8_1 ( A, B, Carry, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Carry;
  output [31:0] S;
  output Cout;

  assign Cout = Carry[8];

  carry_select_N4_0_1 CS_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Carry[0]), .S(S[3:0])
         );
  carry_select_N4_7_1 CS_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Carry[1]), .S(S[7:4])
         );
  carry_select_N4_6_1 CS_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Carry[2]), .S(
        S[11:8]) );
  carry_select_N4_5 CS_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Carry[3]), .S(
        S[15:12]) );
  carry_select_N4_4 CS_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Carry[4]), .S(
        S[19:16]) );
  carry_select_N4_3 CS_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Carry[5]), .S(
        S[23:20]) );
  carry_select_N4_2 CS_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Carry[6]), .S(
        S[27:24]) );
  carry_select_N4_1 CS_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Carry[7]), .S(
        S[31:28]) );
endmodule


module carry_generator_N32_Nblocks8_1 ( A, B, Ci, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, g_cin, p_cin, \Gsignal[1][31] , \Gsignal[1][30] ,
         \Gsignal[1][29] , \Gsignal[1][28] , \Gsignal[1][27] ,
         \Gsignal[1][26] , \Gsignal[1][25] , \Gsignal[1][24] ,
         \Gsignal[1][23] , \Gsignal[1][22] , \Gsignal[1][21] ,
         \Gsignal[1][20] , \Gsignal[1][19] , \Gsignal[1][18] ,
         \Gsignal[1][17] , \Gsignal[1][16] , \Gsignal[1][15] ,
         \Gsignal[1][14] , \Gsignal[1][13] , \Gsignal[1][12] ,
         \Gsignal[1][11] , \Gsignal[1][10] , \Gsignal[1][9] , \Gsignal[1][8] ,
         \Gsignal[1][7] , \Gsignal[1][6] , \Gsignal[1][5] , \Gsignal[1][4] ,
         \Gsignal[1][3] , \Gsignal[1][2] , \Gsignal[1][1] , \Gsignal[1][0] ,
         \Gsignal[2][31] , \Gsignal[2][29] , \Gsignal[2][27] ,
         \Gsignal[2][25] , \Gsignal[2][23] , \Gsignal[2][21] ,
         \Gsignal[2][19] , \Gsignal[2][17] , \Gsignal[2][15] ,
         \Gsignal[2][13] , \Gsignal[2][11] , \Gsignal[2][9] , \Gsignal[2][7] ,
         \Gsignal[2][5] , \Gsignal[2][3] , \Gsignal[2][1] , \Gsignal[3][31] ,
         \Gsignal[3][23] , \Gsignal[3][15] , \Gsignal[3][7] , \Gsignal[4][31] ,
         \Gsignal[4][15] , \Gsignal[5][31] , \Gsignal[5][27] ,
         \Psignal[1][31] , \Psignal[1][30] , \Psignal[1][29] ,
         \Psignal[1][28] , \Psignal[1][27] , \Psignal[1][26] ,
         \Psignal[1][25] , \Psignal[1][24] , \Psignal[1][23] ,
         \Psignal[1][22] , \Psignal[1][21] , \Psignal[1][20] ,
         \Psignal[1][19] , \Psignal[1][18] , \Psignal[1][17] ,
         \Psignal[1][16] , \Psignal[1][15] , \Psignal[1][14] ,
         \Psignal[1][13] , \Psignal[1][12] , \Psignal[1][11] ,
         \Psignal[1][10] , \Psignal[1][9] , \Psignal[1][8] , \Psignal[1][7] ,
         \Psignal[1][6] , \Psignal[1][5] , \Psignal[1][4] , \Psignal[1][3] ,
         \Psignal[1][2] , \Psignal[1][1] , \Psignal[2][31] , \Psignal[2][29] ,
         \Psignal[2][27] , \Psignal[2][25] , \Psignal[2][23] ,
         \Psignal[2][21] , \Psignal[2][19] , \Psignal[2][17] ,
         \Psignal[2][15] , \Psignal[2][13] , \Psignal[2][11] , \Psignal[2][9] ,
         \Psignal[2][7] , \Psignal[2][5] , \Psignal[2][3] , \Psignal[3][31] ,
         \Psignal[3][27] , \Psignal[3][23] , \Psignal[3][19] ,
         \Psignal[3][15] , \Psignal[3][7] , \Psignal[4][31] , \Psignal[4][23] ,
         \Psignal[4][15] , \Psignal[5][31] , \Psignal[5][27] , n8, n10, n12,
         n13, n15;
  assign Cout[0] = Ci;

  PGnet_block_0_1 PGnet_Cin_0 ( .A(A[0]), .B(B[0]), .pout(p_cin), .gout(g_cin)
         );
  G_0_1 GCin_0 ( .gleft(g_cin), .gright(Ci), .pleft(p_cin), .gout(
        \Gsignal[1][0] ) );
  PGnet_block_31_1 PGnet_1 ( .A(A[1]), .B(B[1]), .pout(\Psignal[1][1] ), 
        .gout(\Gsignal[1][1] ) );
  PGnet_block_30_1 PGnet_2 ( .A(A[2]), .B(B[2]), .pout(\Psignal[1][2] ), 
        .gout(\Gsignal[1][2] ) );
  PGnet_block_29 PGnet_3 ( .A(A[3]), .B(B[3]), .pout(\Psignal[1][3] ), .gout(
        \Gsignal[1][3] ) );
  PGnet_block_28 PGnet_4 ( .A(A[4]), .B(B[4]), .pout(\Psignal[1][4] ), .gout(
        \Gsignal[1][4] ) );
  PGnet_block_27 PGnet_5 ( .A(A[5]), .B(B[5]), .pout(\Psignal[1][5] ), .gout(
        \Gsignal[1][5] ) );
  PGnet_block_26 PGnet_6 ( .A(A[6]), .B(B[6]), .pout(\Psignal[1][6] ), .gout(
        \Gsignal[1][6] ) );
  PGnet_block_25 PGnet_7 ( .A(A[7]), .B(B[7]), .pout(\Psignal[1][7] ), .gout(
        \Gsignal[1][7] ) );
  PGnet_block_24 PGnet_8 ( .A(A[8]), .B(B[8]), .pout(\Psignal[1][8] ), .gout(
        \Gsignal[1][8] ) );
  PGnet_block_23 PGnet_9 ( .A(A[9]), .B(B[9]), .pout(\Psignal[1][9] ), .gout(
        \Gsignal[1][9] ) );
  PGnet_block_22 PGnet_10 ( .A(A[10]), .B(B[10]), .pout(\Psignal[1][10] ), 
        .gout(\Gsignal[1][10] ) );
  PGnet_block_21 PGnet_11 ( .A(A[11]), .B(B[11]), .pout(\Psignal[1][11] ), 
        .gout(\Gsignal[1][11] ) );
  PGnet_block_20 PGnet_12 ( .A(A[12]), .B(B[12]), .pout(\Psignal[1][12] ), 
        .gout(\Gsignal[1][12] ) );
  PGnet_block_19 PGnet_13 ( .A(A[13]), .B(B[13]), .pout(\Psignal[1][13] ), 
        .gout(\Gsignal[1][13] ) );
  PGnet_block_18 PGnet_14 ( .A(A[14]), .B(B[14]), .pout(\Psignal[1][14] ), 
        .gout(\Gsignal[1][14] ) );
  PGnet_block_17 PGnet_15 ( .A(A[15]), .B(B[15]), .pout(\Psignal[1][15] ), 
        .gout(\Gsignal[1][15] ) );
  PGnet_block_16 PGnet_16 ( .A(A[16]), .B(B[16]), .pout(\Psignal[1][16] ), 
        .gout(\Gsignal[1][16] ) );
  PGnet_block_15 PGnet_17 ( .A(A[17]), .B(B[17]), .pout(\Psignal[1][17] ), 
        .gout(\Gsignal[1][17] ) );
  PGnet_block_14 PGnet_18 ( .A(A[18]), .B(B[18]), .pout(\Psignal[1][18] ), 
        .gout(\Gsignal[1][18] ) );
  PGnet_block_13 PGnet_19 ( .A(A[19]), .B(B[19]), .pout(\Psignal[1][19] ), 
        .gout(\Gsignal[1][19] ) );
  PGnet_block_12 PGnet_20 ( .A(A[20]), .B(B[20]), .pout(\Psignal[1][20] ), 
        .gout(\Gsignal[1][20] ) );
  PGnet_block_11 PGnet_21 ( .A(A[21]), .B(B[21]), .pout(\Psignal[1][21] ), 
        .gout(\Gsignal[1][21] ) );
  PGnet_block_10 PGnet_22 ( .A(A[22]), .B(B[22]), .pout(\Psignal[1][22] ), 
        .gout(\Gsignal[1][22] ) );
  PGnet_block_9 PGnet_23 ( .A(A[23]), .B(B[23]), .pout(\Psignal[1][23] ), 
        .gout(\Gsignal[1][23] ) );
  PGnet_block_8 PGnet_24 ( .A(A[24]), .B(B[24]), .pout(\Psignal[1][24] ), 
        .gout(\Gsignal[1][24] ) );
  PGnet_block_7 PGnet_25 ( .A(A[25]), .B(B[25]), .pout(\Psignal[1][25] ), 
        .gout(\Gsignal[1][25] ) );
  PGnet_block_6 PGnet_26 ( .A(A[26]), .B(B[26]), .pout(\Psignal[1][26] ), 
        .gout(\Gsignal[1][26] ) );
  PGnet_block_5 PGnet_27 ( .A(A[27]), .B(B[27]), .pout(\Psignal[1][27] ), 
        .gout(\Gsignal[1][27] ) );
  PGnet_block_4 PGnet_28 ( .A(A[28]), .B(B[28]), .pout(\Psignal[1][28] ), 
        .gout(\Gsignal[1][28] ) );
  PGnet_block_3 PGnet_29 ( .A(A[29]), .B(B[29]), .pout(\Psignal[1][29] ), 
        .gout(\Gsignal[1][29] ) );
  PGnet_block_2 PGnet_30 ( .A(A[30]), .B(B[30]), .pout(\Psignal[1][30] ), 
        .gout(\Gsignal[1][30] ) );
  PGnet_block_1 PGnet_31 ( .A(A[31]), .B(B[31]), .pout(\Psignal[1][31] ), 
        .gout(\Gsignal[1][31] ) );
  G_2 Gblock_1_1 ( .gleft(\Gsignal[1][1] ), .gright(\Gsignal[1][0] ), .pleft(
        \Psignal[1][1] ), .gout(\Gsignal[2][1] ) );
  PG_0_1 PGblock_1_3 ( .gleft(\Gsignal[1][3] ), .gright(\Gsignal[1][2] ), 
        .pleft(\Psignal[1][3] ), .pright(\Psignal[1][2] ), .pout(
        \Psignal[2][3] ), .gout(\Gsignal[2][3] ) );
  PG_26_1 PGblock_1_5 ( .gleft(\Gsignal[1][5] ), .gright(\Gsignal[1][4] ), 
        .pleft(\Psignal[1][5] ), .pright(\Psignal[1][4] ), .pout(
        \Psignal[2][5] ), .gout(\Gsignal[2][5] ) );
  PG_25_1 PGblock_1_7 ( .gleft(\Gsignal[1][7] ), .gright(\Gsignal[1][6] ), 
        .pleft(\Psignal[1][7] ), .pright(\Psignal[1][6] ), .pout(
        \Psignal[2][7] ), .gout(\Gsignal[2][7] ) );
  PG_24_1 PGblock_1_9 ( .gleft(\Gsignal[1][9] ), .gright(\Gsignal[1][8] ), 
        .pleft(\Psignal[1][9] ), .pright(\Psignal[1][8] ), .pout(
        \Psignal[2][9] ), .gout(\Gsignal[2][9] ) );
  PG_12 PGblock_1_11 ( .gleft(\Gsignal[1][11] ), .gright(\Gsignal[1][10] ), 
        .pleft(\Psignal[1][11] ), .pright(\Psignal[1][10] ), .pout(
        \Psignal[2][11] ), .gout(\Gsignal[2][11] ) );
  PG_22_1 PGblock_1_13 ( .gleft(\Gsignal[1][13] ), .gright(\Gsignal[1][12] ), 
        .pleft(\Psignal[1][13] ), .pright(\Psignal[1][12] ), .pout(
        \Psignal[2][13] ), .gout(\Gsignal[2][13] ) );
  PG_21_1 PGblock_1_15 ( .gleft(\Gsignal[1][15] ), .gright(\Gsignal[1][14] ), 
        .pleft(\Psignal[1][15] ), .pright(\Psignal[1][14] ), .pout(
        \Psignal[2][15] ), .gout(\Gsignal[2][15] ) );
  PG_23 PGblock_1_17 ( .gleft(\Gsignal[1][17] ), .gright(\Gsignal[1][16] ), 
        .pleft(\Psignal[1][17] ), .pright(\Psignal[1][16] ), .pout(
        \Psignal[2][17] ), .gout(\Gsignal[2][17] ) );
  PG_11 PGblock_1_19 ( .gleft(\Gsignal[1][19] ), .gright(\Gsignal[1][18] ), 
        .pleft(\Psignal[1][19] ), .pright(\Psignal[1][18] ), .pout(
        \Psignal[2][19] ), .gout(\Gsignal[2][19] ) );
  PG_18_1 PGblock_1_21 ( .gleft(\Gsignal[1][21] ), .gright(\Gsignal[1][20] ), 
        .pleft(\Psignal[1][21] ), .pright(\Psignal[1][20] ), .pout(
        \Psignal[2][21] ), .gout(\Gsignal[2][21] ) );
  PG_20 PGblock_1_23 ( .gleft(\Gsignal[1][23] ), .gright(\Gsignal[1][22] ), 
        .pleft(\Psignal[1][23] ), .pright(\Psignal[1][22] ), .pout(
        \Psignal[2][23] ), .gout(\Gsignal[2][23] ) );
  PG_10 PGblock_1_25 ( .gleft(\Gsignal[1][25] ), .gright(\Gsignal[1][24] ), 
        .pleft(\Psignal[1][25] ), .pright(\Psignal[1][24] ), .pout(
        \Psignal[2][25] ), .gout(\Gsignal[2][25] ) );
  PG_9 PGblock_1_27 ( .gleft(\Gsignal[1][27] ), .gright(\Gsignal[1][26] ), 
        .pleft(\Psignal[1][27] ), .pright(\Psignal[1][26] ), .pout(
        \Psignal[2][27] ), .gout(\Gsignal[2][27] ) );
  PG_8 PGblock_1_29 ( .gleft(\Gsignal[1][29] ), .gright(\Gsignal[1][28] ), 
        .pleft(\Psignal[1][29] ), .pright(\Psignal[1][28] ), .pout(
        \Psignal[2][29] ), .gout(\Gsignal[2][29] ) );
  PG_7 PGblock_1_31 ( .gleft(\Gsignal[1][31] ), .gright(\Gsignal[1][30] ), 
        .pleft(\Psignal[1][31] ), .pright(\Psignal[1][30] ), .pout(
        \Psignal[2][31] ), .gout(\Gsignal[2][31] ) );
  G_8_1 Gblock_2_3 ( .gleft(\Gsignal[2][3] ), .gright(\Gsignal[2][1] ), 
        .pleft(\Psignal[2][3] ), .gout(Cout[1]) );
  PG_19 PGblock_2_7 ( .gleft(\Gsignal[2][7] ), .gright(\Gsignal[2][5] ), 
        .pleft(\Psignal[2][7] ), .pright(\Psignal[2][5] ), .pout(
        \Psignal[3][7] ), .gout(\Gsignal[3][7] ) );
  PG_17 PGblock_2_11 ( .gleft(\Gsignal[2][11] ), .gright(\Gsignal[2][9] ), 
        .pleft(\Psignal[2][11] ), .pright(\Psignal[2][9] ), .pout(n8), .gout(
        n10) );
  PG_16 PGblock_2_15 ( .gleft(\Gsignal[2][15] ), .gright(\Gsignal[2][13] ), 
        .pleft(\Psignal[2][15] ), .pright(\Psignal[2][13] ), .pout(
        \Psignal[3][15] ), .gout(\Gsignal[3][15] ) );
  PG_15 PGblock_2_19 ( .gleft(\Gsignal[2][19] ), .gright(\Gsignal[2][17] ), 
        .pleft(\Psignal[2][19] ), .pright(\Psignal[2][17] ), .pout(
        \Psignal[3][19] ), .gout(n13) );
  PG_14 PGblock_2_23 ( .gleft(\Gsignal[2][23] ), .gright(\Gsignal[2][21] ), 
        .pleft(\Psignal[2][23] ), .pright(\Psignal[2][21] ), .pout(
        \Psignal[3][23] ), .gout(\Gsignal[3][23] ) );
  PG_6 PGblock_2_27 ( .gleft(\Gsignal[2][27] ), .gright(\Gsignal[2][25] ), 
        .pleft(\Psignal[2][27] ), .pright(\Psignal[2][25] ), .pout(
        \Psignal[3][27] ), .gout(n12) );
  PG_5 PGblock_2_31 ( .gleft(\Gsignal[2][31] ), .gright(\Gsignal[2][29] ), 
        .pleft(\Psignal[2][31] ), .pright(\Psignal[2][29] ), .pout(
        \Psignal[3][31] ), .gout(\Gsignal[3][31] ) );
  G_1 Gblock_3_7 ( .gleft(\Gsignal[3][7] ), .gright(Cout[1]), .pleft(
        \Psignal[3][7] ), .gout(Cout[2]) );
  PG_13 PGblock_3_15 ( .gleft(\Gsignal[3][15] ), .gright(n10), .pleft(
        \Psignal[3][15] ), .pright(n8), .pout(\Psignal[4][15] ), .gout(
        \Gsignal[4][15] ) );
  PG_4_1 PGblock_3_23 ( .gleft(\Gsignal[3][23] ), .gright(n13), .pleft(
        \Psignal[3][23] ), .pright(\Psignal[3][19] ), .pout(\Psignal[4][23] ), 
        .gout(n15) );
  PG_3 PGblock_3_31 ( .gleft(\Gsignal[3][31] ), .gright(n12), .pleft(
        \Psignal[3][31] ), .pright(\Psignal[3][27] ), .pout(\Psignal[4][31] ), 
        .gout(\Gsignal[4][31] ) );
  G_6_1 Gblock_4_11 ( .gleft(n10), .gright(Cout[2]), .pleft(n8), .gout(Cout[3]) );
  G_5_1 Gblock_4_15 ( .gleft(\Gsignal[4][15] ), .gright(Cout[2]), .pleft(
        \Psignal[4][15] ), .gout(Cout[4]) );
  PG_1 PGblock_4_27 ( .gleft(n12), .gright(n15), .pleft(\Psignal[3][27] ), 
        .pright(\Psignal[4][23] ), .pout(\Psignal[5][27] ), .gout(
        \Gsignal[5][27] ) );
  PG_2 PGblock_4_31 ( .gleft(\Gsignal[4][31] ), .gright(n15), .pleft(
        \Psignal[4][31] ), .pright(\Psignal[4][23] ), .pout(\Psignal[5][31] ), 
        .gout(\Gsignal[5][31] ) );
  G_9 Gblock_5_19 ( .gleft(n13), .gright(Cout[4]), .pleft(\Psignal[3][19] ), 
        .gout(Cout[5]) );
  G_7 Gblock_5_23 ( .gleft(n15), .gright(Cout[4]), .pleft(\Psignal[4][23] ), 
        .gout(Cout[6]) );
  G_4 Gblock_5_27 ( .gleft(\Gsignal[5][27] ), .gright(Cout[4]), .pleft(
        \Psignal[5][27] ), .gout(Cout[7]) );
  G_3 Gblock_5_31 ( .gleft(\Gsignal[5][31] ), .gright(Cout[4]), .pleft(
        \Psignal[5][31] ), .gout(Cout[8]) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U3 ( .A(Ci), .B(n13), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n13) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n13), .B2(Ci), .ZN(n12) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n16, n17;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n16), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n16) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net26715, n2, n3;
  assign net26715 = A;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(net26715), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(net26715), .A2(B), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net25115, n2, n3;
  assign net25115 = B;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(net25115), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(net25115), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n13, n14;

  XOR2_X1 U3 ( .A(Ci), .B(n14), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n14) );
  INV_X1 U1 ( .A(n13), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n14), .B2(Ci), .ZN(n13) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n16, n17;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n16), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n16) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n16, n17;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n16), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n16) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n15, n16;

  XOR2_X1 U3 ( .A(Ci), .B(n16), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n16) );
  INV_X1 U1 ( .A(n15), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n16), .B2(Ci), .ZN(n15) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U3 ( .A(Ci), .B(n10), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  INV_X1 U1 ( .A(n9), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n9) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U3 ( .A(Ci), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  INV_X1 U1 ( .A(n8), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n12), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
  INV_X1 U1 ( .A(n11), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n11) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n10), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n10) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module sum_generator_Nbits32_Nblocks8_0 ( A, B, Carry, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Carry;
  output [31:0] S;
  output Cout;

  assign Cout = Carry[8];

  carry_select_N4_0_0 CS_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Carry[0]), .S(S[3:0])
         );
  carry_select_N4_7_0 CS_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Carry[1]), .S(S[7:4])
         );
  carry_select_N4_6_0 CS_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Carry[2]), .S(
        S[11:8]) );
  carry_select_N4_12 CS_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Carry[3]), .S(
        S[15:12]) );
  carry_select_N4_11 CS_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Carry[4]), .S(
        S[19:16]) );
  carry_select_N4_10 CS_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Carry[5]), .S(
        S[23:20]) );
  carry_select_N4_9 CS_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Carry[6]), .S(
        S[27:24]) );
  carry_select_N4_8 CS_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Carry[7]), .S(
        S[31:28]) );
endmodule


module carry_generator_N32_Nblocks8_0 ( A, B, Ci, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, g_cin, p_cin, \Gsignal[1][31] , \Gsignal[1][30] ,
         \Gsignal[1][29] , \Gsignal[1][28] , \Gsignal[1][27] ,
         \Gsignal[1][26] , \Gsignal[1][25] , \Gsignal[1][24] ,
         \Gsignal[1][23] , \Gsignal[1][22] , \Gsignal[1][21] ,
         \Gsignal[1][20] , \Gsignal[1][19] , \Gsignal[1][18] ,
         \Gsignal[1][17] , \Gsignal[1][16] , \Gsignal[1][15] ,
         \Gsignal[1][14] , \Gsignal[1][13] , \Gsignal[1][12] ,
         \Gsignal[1][11] , \Gsignal[1][10] , \Gsignal[1][9] , \Gsignal[1][8] ,
         \Gsignal[1][7] , \Gsignal[1][6] , \Gsignal[1][5] , \Gsignal[1][4] ,
         \Gsignal[1][3] , \Gsignal[1][2] , \Gsignal[1][1] , \Gsignal[1][0] ,
         \Gsignal[2][31] , \Gsignal[2][29] , \Gsignal[2][27] ,
         \Gsignal[2][25] , \Gsignal[2][23] , \Gsignal[2][21] ,
         \Gsignal[2][19] , \Gsignal[2][17] , \Gsignal[2][15] ,
         \Gsignal[2][13] , \Gsignal[2][11] , \Gsignal[2][9] , \Gsignal[2][7] ,
         \Gsignal[2][5] , \Gsignal[2][3] , \Gsignal[2][1] , \Gsignal[3][31] ,
         \Gsignal[3][23] , \Gsignal[3][15] , \Gsignal[3][7] , \Gsignal[4][31] ,
         \Gsignal[4][15] , \Gsignal[5][31] , \Gsignal[5][27] ,
         \Psignal[1][31] , \Psignal[1][30] , \Psignal[1][29] ,
         \Psignal[1][28] , \Psignal[1][27] , \Psignal[1][26] ,
         \Psignal[1][25] , \Psignal[1][24] , \Psignal[1][23] ,
         \Psignal[1][22] , \Psignal[1][21] , \Psignal[1][20] ,
         \Psignal[1][19] , \Psignal[1][18] , \Psignal[1][17] ,
         \Psignal[1][16] , \Psignal[1][15] , \Psignal[1][14] ,
         \Psignal[1][13] , \Psignal[1][12] , \Psignal[1][11] ,
         \Psignal[1][10] , \Psignal[1][9] , \Psignal[1][8] , \Psignal[1][7] ,
         \Psignal[1][6] , \Psignal[1][5] , \Psignal[1][4] , \Psignal[1][3] ,
         \Psignal[1][2] , \Psignal[1][1] , \Psignal[2][31] , \Psignal[2][29] ,
         \Psignal[2][27] , \Psignal[2][25] , \Psignal[2][23] ,
         \Psignal[2][21] , \Psignal[2][19] , \Psignal[2][17] ,
         \Psignal[2][15] , \Psignal[2][13] , \Psignal[2][11] , \Psignal[2][9] ,
         \Psignal[2][7] , \Psignal[2][5] , \Psignal[2][3] , \Psignal[3][31] ,
         \Psignal[3][27] , \Psignal[3][23] , \Psignal[3][19] ,
         \Psignal[3][15] , \Psignal[3][7] , \Psignal[4][31] , \Psignal[4][23] ,
         \Psignal[4][15] , \Psignal[5][31] , \Psignal[5][27] , n8, n10, n12,
         n13, n15;
  assign Cout[0] = Ci;

  PGnet_block_0_0 PGnet_Cin_0 ( .A(A[0]), .B(B[0]), .pout(p_cin), .gout(g_cin)
         );
  G_0_0 GCin_0 ( .gleft(g_cin), .gright(Ci), .pleft(p_cin), .gout(
        \Gsignal[1][0] ) );
  PGnet_block_31_0 PGnet_1 ( .A(A[1]), .B(B[1]), .pout(\Psignal[1][1] ), 
        .gout(\Gsignal[1][1] ) );
  PGnet_block_30_0 PGnet_2 ( .A(A[2]), .B(B[2]), .pout(\Psignal[1][2] ), 
        .gout(\Gsignal[1][2] ) );
  PGnet_block_60 PGnet_3 ( .A(A[3]), .B(B[3]), .pout(\Psignal[1][3] ), .gout(
        \Gsignal[1][3] ) );
  PGnet_block_59 PGnet_4 ( .A(A[4]), .B(B[4]), .pout(\Psignal[1][4] ), .gout(
        \Gsignal[1][4] ) );
  PGnet_block_58 PGnet_5 ( .A(A[5]), .B(B[5]), .pout(\Psignal[1][5] ), .gout(
        \Gsignal[1][5] ) );
  PGnet_block_57 PGnet_6 ( .A(A[6]), .B(B[6]), .pout(\Psignal[1][6] ), .gout(
        \Gsignal[1][6] ) );
  PGnet_block_56 PGnet_7 ( .A(A[7]), .B(B[7]), .pout(\Psignal[1][7] ), .gout(
        \Gsignal[1][7] ) );
  PGnet_block_55 PGnet_8 ( .A(A[8]), .B(B[8]), .pout(\Psignal[1][8] ), .gout(
        \Gsignal[1][8] ) );
  PGnet_block_54 PGnet_9 ( .A(A[9]), .B(B[9]), .pout(\Psignal[1][9] ), .gout(
        \Gsignal[1][9] ) );
  PGnet_block_53 PGnet_10 ( .A(A[10]), .B(B[10]), .pout(\Psignal[1][10] ), 
        .gout(\Gsignal[1][10] ) );
  PGnet_block_52 PGnet_11 ( .A(A[11]), .B(B[11]), .pout(\Psignal[1][11] ), 
        .gout(\Gsignal[1][11] ) );
  PGnet_block_51 PGnet_12 ( .A(A[12]), .B(B[12]), .pout(\Psignal[1][12] ), 
        .gout(\Gsignal[1][12] ) );
  PGnet_block_50 PGnet_13 ( .A(A[13]), .B(B[13]), .pout(\Psignal[1][13] ), 
        .gout(\Gsignal[1][13] ) );
  PGnet_block_49 PGnet_14 ( .A(A[14]), .B(B[14]), .pout(\Psignal[1][14] ), 
        .gout(\Gsignal[1][14] ) );
  PGnet_block_48 PGnet_15 ( .A(A[15]), .B(B[15]), .pout(\Psignal[1][15] ), 
        .gout(\Gsignal[1][15] ) );
  PGnet_block_47 PGnet_16 ( .A(A[16]), .B(B[16]), .pout(\Psignal[1][16] ), 
        .gout(\Gsignal[1][16] ) );
  PGnet_block_46 PGnet_17 ( .A(A[17]), .B(B[17]), .pout(\Psignal[1][17] ), 
        .gout(\Gsignal[1][17] ) );
  PGnet_block_45 PGnet_18 ( .A(A[18]), .B(B[18]), .pout(\Psignal[1][18] ), 
        .gout(\Gsignal[1][18] ) );
  PGnet_block_44 PGnet_19 ( .A(A[19]), .B(B[19]), .pout(\Psignal[1][19] ), 
        .gout(\Gsignal[1][19] ) );
  PGnet_block_43 PGnet_20 ( .A(A[20]), .B(B[20]), .pout(\Psignal[1][20] ), 
        .gout(\Gsignal[1][20] ) );
  PGnet_block_42 PGnet_21 ( .A(A[21]), .B(B[21]), .pout(\Psignal[1][21] ), 
        .gout(\Gsignal[1][21] ) );
  PGnet_block_41 PGnet_22 ( .A(A[22]), .B(B[22]), .pout(\Psignal[1][22] ), 
        .gout(\Gsignal[1][22] ) );
  PGnet_block_40 PGnet_23 ( .A(A[23]), .B(B[23]), .pout(\Psignal[1][23] ), 
        .gout(\Gsignal[1][23] ) );
  PGnet_block_39 PGnet_24 ( .A(A[24]), .B(B[24]), .pout(\Psignal[1][24] ), 
        .gout(\Gsignal[1][24] ) );
  PGnet_block_38 PGnet_25 ( .A(A[25]), .B(B[25]), .pout(\Psignal[1][25] ), 
        .gout(\Gsignal[1][25] ) );
  PGnet_block_37 PGnet_26 ( .A(A[26]), .B(B[26]), .pout(\Psignal[1][26] ), 
        .gout(\Gsignal[1][26] ) );
  PGnet_block_36 PGnet_27 ( .A(A[27]), .B(B[27]), .pout(\Psignal[1][27] ), 
        .gout(\Gsignal[1][27] ) );
  PGnet_block_35 PGnet_28 ( .A(A[28]), .B(B[28]), .pout(\Psignal[1][28] ), 
        .gout(\Gsignal[1][28] ) );
  PGnet_block_34 PGnet_29 ( .A(A[29]), .B(B[29]), .pout(\Psignal[1][29] ), 
        .gout(\Gsignal[1][29] ) );
  PGnet_block_33 PGnet_30 ( .A(A[30]), .B(B[30]), .pout(\Psignal[1][30] ), 
        .gout(\Gsignal[1][30] ) );
  PGnet_block_32 PGnet_31 ( .A(A[31]), .B(B[31]), .pout(\Psignal[1][31] ), 
        .gout(\Gsignal[1][31] ) );
  G_15 Gblock_1_1 ( .gleft(\Gsignal[1][1] ), .gright(\Gsignal[1][0] ), .pleft(
        \Psignal[1][1] ), .gout(\Gsignal[2][1] ) );
  PG_0_0 PGblock_1_3 ( .gleft(\Gsignal[1][3] ), .gright(\Gsignal[1][2] ), 
        .pleft(\Psignal[1][3] ), .pright(\Psignal[1][2] ), .pout(
        \Psignal[2][3] ), .gout(\Gsignal[2][3] ) );
  PG_26_0 PGblock_1_5 ( .gleft(\Gsignal[1][5] ), .gright(\Gsignal[1][4] ), 
        .pleft(\Psignal[1][5] ), .pright(\Psignal[1][4] ), .pout(
        \Psignal[2][5] ), .gout(\Gsignal[2][5] ) );
  PG_25_0 PGblock_1_7 ( .gleft(\Gsignal[1][7] ), .gright(\Gsignal[1][6] ), 
        .pleft(\Psignal[1][7] ), .pright(\Psignal[1][6] ), .pout(
        \Psignal[2][7] ), .gout(\Gsignal[2][7] ) );
  PG_24_0 PGblock_1_9 ( .gleft(\Gsignal[1][9] ), .gright(\Gsignal[1][8] ), 
        .pleft(\Psignal[1][9] ), .pright(\Psignal[1][8] ), .pout(
        \Psignal[2][9] ), .gout(\Gsignal[2][9] ) );
  PG_45 PGblock_1_11 ( .gleft(\Gsignal[1][11] ), .gright(\Gsignal[1][10] ), 
        .pleft(\Psignal[1][11] ), .pright(\Psignal[1][10] ), .pout(
        \Psignal[2][11] ), .gout(\Gsignal[2][11] ) );
  PG_22_0 PGblock_1_13 ( .gleft(\Gsignal[1][13] ), .gright(\Gsignal[1][12] ), 
        .pleft(\Psignal[1][13] ), .pright(\Psignal[1][12] ), .pout(
        \Psignal[2][13] ), .gout(\Gsignal[2][13] ) );
  PG_21_0 PGblock_1_15 ( .gleft(\Gsignal[1][15] ), .gright(\Gsignal[1][14] ), 
        .pleft(\Psignal[1][15] ), .pright(\Psignal[1][14] ), .pout(
        \Psignal[2][15] ), .gout(\Gsignal[2][15] ) );
  PG_44 PGblock_1_17 ( .gleft(\Gsignal[1][17] ), .gright(\Gsignal[1][16] ), 
        .pleft(\Psignal[1][17] ), .pright(\Psignal[1][16] ), .pout(
        \Psignal[2][17] ), .gout(\Gsignal[2][17] ) );
  PG_43 PGblock_1_19 ( .gleft(\Gsignal[1][19] ), .gright(\Gsignal[1][18] ), 
        .pleft(\Psignal[1][19] ), .pright(\Psignal[1][18] ), .pout(
        \Psignal[2][19] ), .gout(\Gsignal[2][19] ) );
  PG_18_0 PGblock_1_21 ( .gleft(\Gsignal[1][21] ), .gright(\Gsignal[1][20] ), 
        .pleft(\Psignal[1][21] ), .pright(\Psignal[1][20] ), .pout(
        \Psignal[2][21] ), .gout(\Gsignal[2][21] ) );
  PG_42 PGblock_1_23 ( .gleft(\Gsignal[1][23] ), .gright(\Gsignal[1][22] ), 
        .pleft(\Psignal[1][23] ), .pright(\Psignal[1][22] ), .pout(
        \Psignal[2][23] ), .gout(\Gsignal[2][23] ) );
  PG_41 PGblock_1_25 ( .gleft(\Gsignal[1][25] ), .gright(\Gsignal[1][24] ), 
        .pleft(\Psignal[1][25] ), .pright(\Psignal[1][24] ), .pout(
        \Psignal[2][25] ), .gout(\Gsignal[2][25] ) );
  PG_40 PGblock_1_27 ( .gleft(\Gsignal[1][27] ), .gright(\Gsignal[1][26] ), 
        .pleft(\Psignal[1][27] ), .pright(\Psignal[1][26] ), .pout(
        \Psignal[2][27] ), .gout(\Gsignal[2][27] ) );
  PG_39 PGblock_1_29 ( .gleft(\Gsignal[1][29] ), .gright(\Gsignal[1][28] ), 
        .pleft(\Psignal[1][29] ), .pright(\Psignal[1][28] ), .pout(
        \Psignal[2][29] ), .gout(\Gsignal[2][29] ) );
  PG_38 PGblock_1_31 ( .gleft(\Gsignal[1][31] ), .gright(\Gsignal[1][30] ), 
        .pleft(\Psignal[1][31] ), .pright(\Psignal[1][30] ), .pout(
        \Psignal[2][31] ), .gout(\Gsignal[2][31] ) );
  G_8_0 Gblock_2_3 ( .gleft(\Gsignal[2][3] ), .gright(\Gsignal[2][1] ), 
        .pleft(\Psignal[2][3] ), .gout(Cout[1]) );
  PG_37 PGblock_2_7 ( .gleft(\Gsignal[2][7] ), .gright(\Gsignal[2][5] ), 
        .pleft(\Psignal[2][7] ), .pright(\Psignal[2][5] ), .pout(
        \Psignal[3][7] ), .gout(\Gsignal[3][7] ) );
  PG_36 PGblock_2_11 ( .gleft(\Gsignal[2][11] ), .gright(\Gsignal[2][9] ), 
        .pleft(\Psignal[2][11] ), .pright(\Psignal[2][9] ), .pout(n8), .gout(
        n10) );
  PG_35 PGblock_2_15 ( .gleft(\Gsignal[2][15] ), .gright(\Gsignal[2][13] ), 
        .pleft(\Psignal[2][15] ), .pright(\Psignal[2][13] ), .pout(
        \Psignal[3][15] ), .gout(\Gsignal[3][15] ) );
  PG_34 PGblock_2_19 ( .gleft(\Gsignal[2][19] ), .gright(\Gsignal[2][17] ), 
        .pleft(\Psignal[2][19] ), .pright(\Psignal[2][17] ), .pout(
        \Psignal[3][19] ), .gout(n13) );
  PG_33 PGblock_2_23 ( .gleft(\Gsignal[2][23] ), .gright(\Gsignal[2][21] ), 
        .pleft(\Psignal[2][23] ), .pright(\Psignal[2][21] ), .pout(
        \Psignal[3][23] ), .gout(\Gsignal[3][23] ) );
  PG_32 PGblock_2_27 ( .gleft(\Gsignal[2][27] ), .gright(\Gsignal[2][25] ), 
        .pleft(\Psignal[2][27] ), .pright(\Psignal[2][25] ), .pout(
        \Psignal[3][27] ), .gout(n12) );
  PG_31 PGblock_2_31 ( .gleft(\Gsignal[2][31] ), .gright(\Gsignal[2][29] ), 
        .pleft(\Psignal[2][31] ), .pright(\Psignal[2][29] ), .pout(
        \Psignal[3][31] ), .gout(\Gsignal[3][31] ) );
  G_14 Gblock_3_7 ( .gleft(\Gsignal[3][7] ), .gright(Cout[1]), .pleft(
        \Psignal[3][7] ), .gout(Cout[2]) );
  PG_30 PGblock_3_15 ( .gleft(\Gsignal[3][15] ), .gright(n10), .pleft(
        \Psignal[3][15] ), .pright(n8), .pout(\Psignal[4][15] ), .gout(
        \Gsignal[4][15] ) );
  PG_4_0 PGblock_3_23 ( .gleft(\Gsignal[3][23] ), .gright(n13), .pleft(
        \Psignal[3][23] ), .pright(\Psignal[3][19] ), .pout(\Psignal[4][23] ), 
        .gout(n15) );
  PG_29 PGblock_3_31 ( .gleft(\Gsignal[3][31] ), .gright(n12), .pleft(
        \Psignal[3][31] ), .pright(\Psignal[3][27] ), .pout(\Psignal[4][31] ), 
        .gout(\Gsignal[4][31] ) );
  G_6_0 Gblock_4_11 ( .gleft(n10), .gright(Cout[2]), .pleft(n8), .gout(Cout[3]) );
  G_5_0 Gblock_4_15 ( .gleft(\Gsignal[4][15] ), .gright(Cout[2]), .pleft(
        \Psignal[4][15] ), .gout(Cout[4]) );
  PG_28 PGblock_4_27 ( .gleft(n12), .gright(n15), .pleft(\Psignal[3][27] ), 
        .pright(\Psignal[4][23] ), .pout(\Psignal[5][27] ), .gout(
        \Gsignal[5][27] ) );
  PG_27 PGblock_4_31 ( .gleft(\Gsignal[4][31] ), .gright(n15), .pleft(
        \Psignal[4][31] ), .pright(\Psignal[4][23] ), .pout(\Psignal[5][31] ), 
        .gout(\Gsignal[5][31] ) );
  G_13 Gblock_5_19 ( .gleft(n13), .gright(Cout[4]), .pleft(\Psignal[3][19] ), 
        .gout(Cout[5]) );
  G_12 Gblock_5_23 ( .gleft(n15), .gright(Cout[4]), .pleft(\Psignal[4][23] ), 
        .gout(Cout[6]) );
  G_11 Gblock_5_27 ( .gleft(\Gsignal[5][27] ), .gright(Cout[4]), .pleft(
        \Psignal[5][27] ), .gout(Cout[7]) );
  G_10 Gblock_5_31 ( .gleft(\Gsignal[5][31] ), .gright(Cout[4]), .pleft(
        \Psignal[5][31] ), .gout(Cout[8]) );
endmodule


module xor_gate_1 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_2 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_3 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_4 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_5 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_6 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_7 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_8 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_9 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_10 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_11 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_12 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_13 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_14 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_15 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_16 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_17 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_18 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_19 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_20 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_21 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_22 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_23 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_24 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_25 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_26 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_27 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_28 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_29 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_30 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_31 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module xor_gate_0 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module carry_select_N4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum_carry0;
  wire   [3:0] sum_carry1;

  rca_generic_N4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_carry0) );
  rca_generic_N4 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_carry1) );
  MUX21_GENERIC_N4 MUX ( .A(sum_carry1), .B(sum_carry0), .SEL(Ci), .Y(S) );
endmodule


module PG ( gleft, gright, pleft, pright, pout, gout );
  input gleft, gright, pleft, pright;
  output pout, gout;
  wire   N0;

  GTECH_OR2 C7 ( .A(gleft), .B(N0), .Z(gout) );
  GTECH_AND2 C8 ( .A(gright), .B(pleft), .Z(N0) );
  GTECH_AND2 C9 ( .A(pleft), .B(pright), .Z(pout) );
endmodule


module G ( gleft, gright, pleft, gout );
  input gleft, gright, pleft;
  output gout;
  wire   N0;

  GTECH_OR2 C6 ( .A(gleft), .B(N0), .Z(gout) );
  GTECH_AND2 C7 ( .A(gright), .B(pleft), .Z(N0) );
endmodule


module PGnet_block ( A, B, pout, gout );
  input A, B;
  output pout, gout;


  GTECH_AND2 C7 ( .A(A), .B(B), .Z(gout) );
  GTECH_XOR2 C8 ( .A(A), .B(B), .Z(pout) );
endmodule


module shift_thirdLevel ( sel, A, Y );
  input [2:0] sel;
  input [38:0] A;
  output [31:0] Y;
  wire   n40, n41, n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167;

  AND2_X1 U1 ( .A1(sel[2]), .A2(n148), .ZN(n149) );
  INV_X1 U2 ( .A(n157), .ZN(n156) );
  INV_X1 U3 ( .A(n149), .ZN(n154) );
  INV_X1 U4 ( .A(n161), .ZN(n158) );
  INV_X1 U5 ( .A(n153), .ZN(n152) );
  INV_X1 U6 ( .A(n149), .ZN(n155) );
  OAI22_X1 U7 ( .A1(n165), .A2(n126), .B1(sel[0]), .B2(n123), .ZN(Y[15]) );
  OAI22_X1 U8 ( .A1(n166), .A2(n129), .B1(sel[0]), .B2(n126), .ZN(Y[14]) );
  OAI22_X1 U9 ( .A1(n166), .A2(n132), .B1(sel[0]), .B2(n129), .ZN(Y[13]) );
  OAI22_X1 U10 ( .A1(n166), .A2(n135), .B1(sel[0]), .B2(n132), .ZN(Y[12]) );
  OAI22_X1 U11 ( .A1(n166), .A2(n138), .B1(sel[0]), .B2(n135), .ZN(Y[11]) );
  INV_X1 U12 ( .A(n151), .ZN(n150) );
  OAI22_X1 U13 ( .A1(sel[0]), .A2(n40), .B1(n41), .B2(n159), .ZN(Y[9]) );
  OAI22_X1 U14 ( .A1(n161), .A2(n83), .B1(n158), .B2(n74), .ZN(Y[29]) );
  OAI22_X1 U15 ( .A1(n162), .A2(n86), .B1(n158), .B2(n83), .ZN(Y[28]) );
  OAI22_X1 U16 ( .A1(n162), .A2(n89), .B1(n158), .B2(n86), .ZN(Y[27]) );
  OAI22_X1 U17 ( .A1(n162), .A2(n91), .B1(n158), .B2(n89), .ZN(Y[26]) );
  OAI22_X1 U18 ( .A1(n162), .A2(n93), .B1(n158), .B2(n91), .ZN(Y[25]) );
  OAI22_X1 U19 ( .A1(n163), .A2(n96), .B1(n158), .B2(n93), .ZN(Y[24]) );
  OAI22_X1 U20 ( .A1(n163), .A2(n99), .B1(n158), .B2(n96), .ZN(Y[23]) );
  OAI22_X1 U21 ( .A1(n163), .A2(n102), .B1(n158), .B2(n99), .ZN(Y[22]) );
  OAI22_X1 U22 ( .A1(n164), .A2(n105), .B1(n158), .B2(n102), .ZN(Y[21]) );
  OAI22_X1 U23 ( .A1(n164), .A2(n108), .B1(n158), .B2(n105), .ZN(Y[20]) );
  OAI22_X1 U24 ( .A1(n164), .A2(n114), .B1(n158), .B2(n108), .ZN(Y[19]) );
  OAI22_X1 U25 ( .A1(n165), .A2(n117), .B1(n158), .B2(n114), .ZN(Y[18]) );
  OAI22_X1 U26 ( .A1(n165), .A2(n120), .B1(n158), .B2(n117), .ZN(Y[17]) );
  OAI22_X1 U27 ( .A1(n165), .A2(n123), .B1(n158), .B2(n120), .ZN(Y[16]) );
  OAI22_X1 U28 ( .A1(n159), .A2(n43), .B1(n158), .B2(n41), .ZN(Y[8]) );
  OAI22_X1 U29 ( .A1(sel[0]), .A2(n138), .B1(n159), .B2(n40), .ZN(Y[10]) );
  OAI221_X1 U30 ( .B1(A[13]), .B2(n154), .C1(A[11]), .C2(n44), .A(n142), .ZN(
        n138) );
  AOI22_X1 U31 ( .A1(n47), .A2(n50), .B1(n150), .B2(n137), .ZN(n142) );
  OAI221_X1 U32 ( .B1(A[20]), .B2(n155), .C1(A[18]), .C2(n156), .A(n121), .ZN(
        n117) );
  AOI22_X1 U33 ( .A1(n152), .A2(n122), .B1(n150), .B2(n116), .ZN(n121) );
  OAI221_X1 U34 ( .B1(A[19]), .B2(n154), .C1(A[17]), .C2(n156), .A(n124), .ZN(
        n120) );
  AOI22_X1 U35 ( .A1(n152), .A2(n125), .B1(n150), .B2(n119), .ZN(n124) );
  OAI221_X1 U36 ( .B1(A[18]), .B2(n155), .C1(A[16]), .C2(n156), .A(n127), .ZN(
        n123) );
  AOI22_X1 U37 ( .A1(n152), .A2(n128), .B1(n150), .B2(n122), .ZN(n127) );
  OAI221_X1 U38 ( .B1(A[16]), .B2(n154), .C1(A[14]), .C2(n156), .A(n133), .ZN(
        n129) );
  AOI22_X1 U39 ( .A1(n152), .A2(n134), .B1(n150), .B2(n128), .ZN(n133) );
  OAI221_X1 U40 ( .B1(A[15]), .B2(n155), .C1(A[13]), .C2(n156), .A(n136), .ZN(
        n132) );
  AOI22_X1 U41 ( .A1(n152), .A2(n137), .B1(n150), .B2(n131), .ZN(n136) );
  OAI221_X1 U42 ( .B1(A[14]), .B2(n154), .C1(A[12]), .C2(n156), .A(n139), .ZN(
        n135) );
  AOI22_X1 U43 ( .A1(n152), .A2(n140), .B1(n150), .B2(n134), .ZN(n139) );
  OAI221_X1 U44 ( .B1(A[12]), .B2(n154), .C1(A[10]), .C2(n156), .A(n141), .ZN(
        n40) );
  AOI22_X1 U45 ( .A1(n152), .A2(n54), .B1(n150), .B2(n140), .ZN(n141) );
  OAI221_X1 U46 ( .B1(A[8]), .B2(n44), .C1(A[10]), .C2(n154), .A(n52), .ZN(n43) );
  AOI22_X1 U47 ( .A1(n152), .A2(n53), .B1(n49), .B2(n54), .ZN(n52) );
  OAI221_X1 U48 ( .B1(A[32]), .B2(n154), .C1(A[30]), .C2(n156), .A(n84), .ZN(
        n74) );
  AOI22_X1 U49 ( .A1(n152), .A2(n72), .B1(n49), .B2(n85), .ZN(n84) );
  INV_X1 U50 ( .A(A[36]), .ZN(n85) );
  OAI221_X1 U51 ( .B1(A[31]), .B2(n155), .C1(A[29]), .C2(n44), .A(n87), .ZN(
        n83) );
  AOI22_X1 U52 ( .A1(n152), .A2(n79), .B1(n49), .B2(n88), .ZN(n87) );
  INV_X1 U53 ( .A(A[35]), .ZN(n88) );
  OAI221_X1 U54 ( .B1(A[30]), .B2(n155), .C1(A[28]), .C2(n156), .A(n90), .ZN(
        n86) );
  AOI22_X1 U55 ( .A1(n47), .A2(n73), .B1(n49), .B2(n72), .ZN(n90) );
  OAI221_X1 U56 ( .B1(A[29]), .B2(n155), .C1(A[27]), .C2(n44), .A(n92), .ZN(
        n89) );
  AOI22_X1 U57 ( .A1(n47), .A2(n77), .B1(n49), .B2(n79), .ZN(n92) );
  OAI221_X1 U58 ( .B1(A[28]), .B2(n155), .C1(A[26]), .C2(n156), .A(n94), .ZN(
        n91) );
  AOI22_X1 U59 ( .A1(n47), .A2(n95), .B1(n49), .B2(n73), .ZN(n94) );
  OAI221_X1 U60 ( .B1(A[27]), .B2(n155), .C1(A[25]), .C2(n44), .A(n97), .ZN(
        n93) );
  AOI22_X1 U61 ( .A1(n47), .A2(n98), .B1(n49), .B2(n77), .ZN(n97) );
  OAI221_X1 U62 ( .B1(A[26]), .B2(n155), .C1(A[24]), .C2(n156), .A(n100), .ZN(
        n96) );
  AOI22_X1 U63 ( .A1(n47), .A2(n101), .B1(n49), .B2(n95), .ZN(n100) );
  OAI221_X1 U64 ( .B1(A[25]), .B2(n155), .C1(A[23]), .C2(n44), .A(n103), .ZN(
        n99) );
  AOI22_X1 U65 ( .A1(n47), .A2(n104), .B1(n150), .B2(n98), .ZN(n103) );
  OAI221_X1 U66 ( .B1(A[24]), .B2(n155), .C1(A[22]), .C2(n156), .A(n106), .ZN(
        n102) );
  AOI22_X1 U67 ( .A1(n47), .A2(n107), .B1(n150), .B2(n101), .ZN(n106) );
  OAI221_X1 U68 ( .B1(A[23]), .B2(n155), .C1(A[21]), .C2(n156), .A(n109), .ZN(
        n105) );
  AOI22_X1 U69 ( .A1(n152), .A2(n110), .B1(n150), .B2(n104), .ZN(n109) );
  OAI221_X1 U70 ( .B1(A[22]), .B2(n155), .C1(A[20]), .C2(n156), .A(n115), .ZN(
        n108) );
  AOI22_X1 U71 ( .A1(n152), .A2(n116), .B1(n150), .B2(n107), .ZN(n115) );
  OAI221_X1 U72 ( .B1(A[21]), .B2(n155), .C1(A[19]), .C2(n156), .A(n118), .ZN(
        n114) );
  AOI22_X1 U73 ( .A1(n152), .A2(n119), .B1(n150), .B2(n110), .ZN(n118) );
  OAI221_X1 U74 ( .B1(A[17]), .B2(n155), .C1(A[15]), .C2(n156), .A(n130), .ZN(
        n126) );
  AOI22_X1 U75 ( .A1(n152), .A2(n131), .B1(n150), .B2(n125), .ZN(n130) );
  OAI221_X1 U76 ( .B1(A[9]), .B2(n44), .C1(A[11]), .C2(n154), .A(n46), .ZN(n41) );
  AOI22_X1 U77 ( .A1(n152), .A2(n48), .B1(n150), .B2(n50), .ZN(n46) );
  OAI22_X1 U78 ( .A1(n163), .A2(n74), .B1(n158), .B2(n69), .ZN(Y[30]) );
  OAI22_X1 U79 ( .A1(n160), .A2(n51), .B1(n158), .B2(n43), .ZN(Y[7]) );
  OAI22_X1 U80 ( .A1(n160), .A2(n55), .B1(n158), .B2(n51), .ZN(Y[6]) );
  OAI22_X1 U81 ( .A1(n160), .A2(n58), .B1(n158), .B2(n55), .ZN(Y[5]) );
  OAI22_X1 U82 ( .A1(n160), .A2(n61), .B1(n158), .B2(n58), .ZN(Y[4]) );
  OAI22_X1 U83 ( .A1(n161), .A2(n66), .B1(sel[0]), .B2(n61), .ZN(Y[3]) );
  OAI22_X1 U84 ( .A1(n161), .A2(n80), .B1(sel[0]), .B2(n66), .ZN(Y[2]) );
  OAI22_X1 U85 ( .A1(n164), .A2(n111), .B1(n158), .B2(n80), .ZN(Y[1]) );
  BUF_X1 U86 ( .A(n167), .Z(n160) );
  BUF_X1 U87 ( .A(n167), .Z(n161) );
  BUF_X1 U88 ( .A(n165), .Z(n162) );
  INV_X1 U89 ( .A(A[31]), .ZN(n77) );
  INV_X1 U90 ( .A(A[32]), .ZN(n73) );
  BUF_X1 U91 ( .A(n167), .Z(n159) );
  BUF_X1 U92 ( .A(n166), .Z(n163) );
  BUF_X1 U93 ( .A(n167), .Z(n165) );
  BUF_X1 U94 ( .A(n167), .Z(n166) );
  BUF_X1 U95 ( .A(n167), .Z(n164) );
  INV_X1 U96 ( .A(A[30]), .ZN(n95) );
  INV_X1 U97 ( .A(A[29]), .ZN(n98) );
  INV_X1 U98 ( .A(A[28]), .ZN(n101) );
  INV_X1 U99 ( .A(A[27]), .ZN(n104) );
  INV_X1 U100 ( .A(A[26]), .ZN(n107) );
  INV_X1 U101 ( .A(A[25]), .ZN(n110) );
  INV_X1 U102 ( .A(A[24]), .ZN(n116) );
  INV_X1 U103 ( .A(A[23]), .ZN(n119) );
  INV_X1 U104 ( .A(A[22]), .ZN(n122) );
  INV_X1 U105 ( .A(A[21]), .ZN(n125) );
  INV_X1 U106 ( .A(A[20]), .ZN(n128) );
  INV_X1 U107 ( .A(A[19]), .ZN(n131) );
  INV_X1 U108 ( .A(A[18]), .ZN(n134) );
  INV_X1 U109 ( .A(A[17]), .ZN(n137) );
  INV_X1 U110 ( .A(A[16]), .ZN(n140) );
  INV_X1 U111 ( .A(A[15]), .ZN(n50) );
  INV_X1 U112 ( .A(A[14]), .ZN(n54) );
  INV_X1 U113 ( .A(A[13]), .ZN(n48) );
  INV_X1 U114 ( .A(A[12]), .ZN(n53) );
  OAI221_X1 U115 ( .B1(A[1]), .B2(n44), .C1(A[3]), .C2(n154), .A(n146), .ZN(
        n111) );
  INV_X1 U116 ( .A(n147), .ZN(n146) );
  OAI22_X1 U117 ( .A1(n153), .A2(A[5]), .B1(n151), .B2(A[7]), .ZN(n147) );
  OAI221_X1 U118 ( .B1(A[3]), .B2(n44), .C1(A[5]), .C2(n154), .A(n81), .ZN(n66) );
  INV_X1 U119 ( .A(n82), .ZN(n81) );
  OAI22_X1 U120 ( .A1(n153), .A2(A[7]), .B1(n151), .B2(A[9]), .ZN(n82) );
  OAI221_X1 U121 ( .B1(A[2]), .B2(n44), .C1(A[4]), .C2(n154), .A(n112), .ZN(
        n80) );
  INV_X1 U122 ( .A(n113), .ZN(n112) );
  OAI22_X1 U123 ( .A1(n153), .A2(A[6]), .B1(n151), .B2(A[8]), .ZN(n113) );
  OAI221_X1 U124 ( .B1(A[9]), .B2(n154), .C1(A[7]), .C2(n44), .A(n56), .ZN(n51) );
  AOI22_X1 U125 ( .A1(n47), .A2(n57), .B1(n49), .B2(n48), .ZN(n56) );
  INV_X1 U126 ( .A(A[11]), .ZN(n57) );
  OAI221_X1 U127 ( .B1(A[8]), .B2(n154), .C1(A[6]), .C2(n44), .A(n59), .ZN(n55) );
  AOI22_X1 U128 ( .A1(n152), .A2(n60), .B1(n150), .B2(n53), .ZN(n59) );
  INV_X1 U129 ( .A(A[10]), .ZN(n60) );
  OAI221_X1 U130 ( .B1(A[7]), .B2(n154), .C1(A[5]), .C2(n44), .A(n62), .ZN(n58) );
  INV_X1 U131 ( .A(n63), .ZN(n62) );
  OAI22_X1 U132 ( .A1(n153), .A2(A[9]), .B1(n151), .B2(A[11]), .ZN(n63) );
  OAI221_X1 U133 ( .B1(A[6]), .B2(n154), .C1(A[4]), .C2(n44), .A(n67), .ZN(n61) );
  INV_X1 U134 ( .A(n68), .ZN(n67) );
  OAI22_X1 U135 ( .A1(n153), .A2(A[8]), .B1(n151), .B2(A[10]), .ZN(n68) );
  OAI221_X1 U136 ( .B1(A[35]), .B2(n153), .C1(A[37]), .C2(n151), .A(n75), .ZN(
        n69) );
  AOI22_X1 U137 ( .A1(n157), .A2(n77), .B1(n149), .B2(n79), .ZN(n75) );
  OAI22_X1 U138 ( .A1(n161), .A2(n69), .B1(n158), .B2(n70), .ZN(Y[31]) );
  AOI221_X1 U139 ( .B1(A[36]), .B2(n47), .C1(A[38]), .C2(n49), .A(n71), .ZN(
        n70) );
  OAI22_X1 U140 ( .A1(n154), .A2(n72), .B1(n44), .B2(n73), .ZN(n71) );
  OAI22_X1 U141 ( .A1(sel[0]), .A2(n111), .B1(n143), .B2(n159), .ZN(Y[0]) );
  AOI221_X1 U142 ( .B1(A[0]), .B2(n157), .C1(A[2]), .C2(n149), .A(n144), .ZN(
        n143) );
  INV_X1 U143 ( .A(n145), .ZN(n144) );
  NOR2_X1 U144 ( .A1(sel[1]), .A2(sel[2]), .ZN(n49) );
  NOR2_X1 U145 ( .A1(n148), .A2(sel[2]), .ZN(n47) );
  AOI22_X1 U146 ( .A1(n49), .A2(A[6]), .B1(n47), .B2(A[4]), .ZN(n145) );
  NAND2_X1 U147 ( .A1(sel[2]), .A2(sel[1]), .ZN(n44) );
  INV_X1 U148 ( .A(A[33]), .ZN(n79) );
  INV_X1 U149 ( .A(A[34]), .ZN(n72) );
  INV_X1 U150 ( .A(sel[1]), .ZN(n148) );
  INV_X1 U151 ( .A(sel[0]), .ZN(n167) );
  INV_X1 U152 ( .A(n49), .ZN(n151) );
  INV_X1 U153 ( .A(n47), .ZN(n153) );
  INV_X1 U154 ( .A(n44), .ZN(n157) );
endmodule


module shift_secondLevel ( sel, mask00, mask08, mask16, Y );
  input [1:0] sel;
  input [38:0] mask00;
  input [38:0] mask08;
  input [38:0] mask16;
  output [38:0] Y;
  wire   n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101;

  BUF_X1 U2 ( .A(n90), .Z(n93) );
  BUF_X1 U3 ( .A(n91), .Z(n94) );
  BUF_X1 U4 ( .A(n90), .Z(n92) );
  BUF_X1 U5 ( .A(n84), .Z(n87) );
  BUF_X1 U6 ( .A(n85), .Z(n88) );
  BUF_X1 U7 ( .A(n84), .Z(n86) );
  BUF_X1 U8 ( .A(n96), .Z(n99) );
  BUF_X1 U9 ( .A(n97), .Z(n100) );
  BUF_X1 U10 ( .A(n96), .Z(n98) );
  BUF_X1 U11 ( .A(n91), .Z(n95) );
  BUF_X1 U12 ( .A(n85), .Z(n89) );
  BUF_X1 U13 ( .A(n97), .Z(n101) );
  INV_X1 U14 ( .A(n71), .ZN(Y[1]) );
  INV_X1 U15 ( .A(n52), .ZN(Y[37]) );
  AOI222_X1 U16 ( .A1(mask00[37]), .A2(n100), .B1(mask16[37]), .B2(n94), .C1(
        mask08[37]), .C2(n88), .ZN(n52) );
  INV_X1 U17 ( .A(n51), .ZN(Y[38]) );
  INV_X1 U18 ( .A(n82), .ZN(Y[0]) );
  INV_X1 U19 ( .A(n41), .ZN(Y[9]) );
  AOI222_X1 U20 ( .A1(mask00[9]), .A2(n101), .B1(mask16[9]), .B2(n95), .C1(
        mask08[9]), .C2(n89), .ZN(n41) );
  INV_X1 U21 ( .A(n45), .ZN(Y[8]) );
  AOI222_X1 U22 ( .A1(mask00[8]), .A2(n101), .B1(mask16[8]), .B2(n95), .C1(
        mask08[8]), .C2(n89), .ZN(n45) );
  INV_X1 U23 ( .A(n80), .ZN(Y[11]) );
  AOI222_X1 U24 ( .A1(mask00[11]), .A2(n98), .B1(mask16[11]), .B2(n92), .C1(
        mask08[11]), .C2(n86), .ZN(n80) );
  INV_X1 U25 ( .A(n81), .ZN(Y[10]) );
  AOI222_X1 U26 ( .A1(mask00[10]), .A2(n98), .B1(mask16[10]), .B2(n92), .C1(
        mask08[10]), .C2(n86), .ZN(n81) );
  INV_X1 U27 ( .A(n59), .ZN(Y[30]) );
  AOI222_X1 U28 ( .A1(mask00[30]), .A2(n99), .B1(mask16[30]), .B2(n93), .C1(
        mask08[30]), .C2(n87), .ZN(n59) );
  INV_X1 U29 ( .A(n61), .ZN(Y[29]) );
  AOI222_X1 U30 ( .A1(mask00[29]), .A2(n99), .B1(mask16[29]), .B2(n93), .C1(
        mask08[29]), .C2(n87), .ZN(n61) );
  INV_X1 U31 ( .A(n62), .ZN(Y[28]) );
  AOI222_X1 U32 ( .A1(mask00[28]), .A2(n99), .B1(mask16[28]), .B2(n93), .C1(
        mask08[28]), .C2(n87), .ZN(n62) );
  INV_X1 U33 ( .A(n63), .ZN(Y[27]) );
  AOI222_X1 U34 ( .A1(mask00[27]), .A2(n99), .B1(mask16[27]), .B2(n93), .C1(
        mask08[27]), .C2(n87), .ZN(n63) );
  INV_X1 U35 ( .A(n64), .ZN(Y[26]) );
  AOI222_X1 U36 ( .A1(mask00[26]), .A2(n99), .B1(mask16[26]), .B2(n93), .C1(
        mask08[26]), .C2(n87), .ZN(n64) );
  INV_X1 U37 ( .A(n65), .ZN(Y[25]) );
  AOI222_X1 U38 ( .A1(mask00[25]), .A2(n99), .B1(mask16[25]), .B2(n93), .C1(
        mask08[25]), .C2(n87), .ZN(n65) );
  INV_X1 U39 ( .A(n66), .ZN(Y[24]) );
  AOI222_X1 U40 ( .A1(mask00[24]), .A2(n99), .B1(mask16[24]), .B2(n93), .C1(
        mask08[24]), .C2(n87), .ZN(n66) );
  INV_X1 U41 ( .A(n67), .ZN(Y[23]) );
  AOI222_X1 U42 ( .A1(mask00[23]), .A2(n99), .B1(mask16[23]), .B2(n93), .C1(
        mask08[23]), .C2(n87), .ZN(n67) );
  INV_X1 U43 ( .A(n68), .ZN(Y[22]) );
  AOI222_X1 U44 ( .A1(mask00[22]), .A2(n99), .B1(mask16[22]), .B2(n93), .C1(
        mask08[22]), .C2(n87), .ZN(n68) );
  INV_X1 U45 ( .A(n69), .ZN(Y[21]) );
  AOI222_X1 U46 ( .A1(mask00[21]), .A2(n99), .B1(mask16[21]), .B2(n93), .C1(
        mask08[21]), .C2(n87), .ZN(n69) );
  INV_X1 U47 ( .A(n70), .ZN(Y[20]) );
  AOI222_X1 U48 ( .A1(mask00[20]), .A2(n99), .B1(mask16[20]), .B2(n93), .C1(
        mask08[20]), .C2(n87), .ZN(n70) );
  INV_X1 U49 ( .A(n72), .ZN(Y[19]) );
  AOI222_X1 U50 ( .A1(mask00[19]), .A2(n98), .B1(mask16[19]), .B2(n92), .C1(
        mask08[19]), .C2(n86), .ZN(n72) );
  INV_X1 U51 ( .A(n73), .ZN(Y[18]) );
  AOI222_X1 U52 ( .A1(mask00[18]), .A2(n98), .B1(mask16[18]), .B2(n92), .C1(
        mask08[18]), .C2(n86), .ZN(n73) );
  INV_X1 U53 ( .A(n74), .ZN(Y[17]) );
  AOI222_X1 U54 ( .A1(mask00[17]), .A2(n98), .B1(mask16[17]), .B2(n92), .C1(
        mask08[17]), .C2(n86), .ZN(n74) );
  INV_X1 U55 ( .A(n75), .ZN(Y[16]) );
  AOI222_X1 U56 ( .A1(mask00[16]), .A2(n98), .B1(mask16[16]), .B2(n92), .C1(
        mask08[16]), .C2(n86), .ZN(n75) );
  INV_X1 U57 ( .A(n76), .ZN(Y[15]) );
  AOI222_X1 U58 ( .A1(mask00[15]), .A2(n98), .B1(mask16[15]), .B2(n92), .C1(
        mask08[15]), .C2(n86), .ZN(n76) );
  INV_X1 U59 ( .A(n77), .ZN(Y[14]) );
  AOI222_X1 U60 ( .A1(mask00[14]), .A2(n98), .B1(mask16[14]), .B2(n92), .C1(
        mask08[14]), .C2(n86), .ZN(n77) );
  INV_X1 U61 ( .A(n78), .ZN(Y[13]) );
  AOI222_X1 U62 ( .A1(mask00[13]), .A2(n98), .B1(mask16[13]), .B2(n92), .C1(
        mask08[13]), .C2(n86), .ZN(n78) );
  INV_X1 U63 ( .A(n79), .ZN(Y[12]) );
  AOI222_X1 U64 ( .A1(mask00[12]), .A2(n98), .B1(mask16[12]), .B2(n92), .C1(
        mask08[12]), .C2(n86), .ZN(n79) );
  INV_X1 U65 ( .A(n56), .ZN(Y[33]) );
  AOI222_X1 U66 ( .A1(mask00[33]), .A2(n100), .B1(mask16[33]), .B2(n94), .C1(
        mask08[33]), .C2(n88), .ZN(n56) );
  INV_X1 U67 ( .A(n55), .ZN(Y[34]) );
  AOI222_X1 U68 ( .A1(mask00[34]), .A2(n100), .B1(mask16[34]), .B2(n94), .C1(
        mask08[34]), .C2(n88), .ZN(n55) );
  INV_X1 U69 ( .A(n54), .ZN(Y[35]) );
  AOI222_X1 U70 ( .A1(mask00[35]), .A2(n100), .B1(mask16[35]), .B2(n94), .C1(
        mask08[35]), .C2(n88), .ZN(n54) );
  INV_X1 U71 ( .A(n57), .ZN(Y[32]) );
  AOI222_X1 U72 ( .A1(mask00[32]), .A2(n100), .B1(mask16[32]), .B2(n94), .C1(
        mask08[32]), .C2(n88), .ZN(n57) );
  INV_X1 U73 ( .A(n58), .ZN(Y[31]) );
  AOI222_X1 U74 ( .A1(mask00[31]), .A2(n100), .B1(mask16[31]), .B2(n94), .C1(
        mask08[31]), .C2(n88), .ZN(n58) );
  INV_X1 U75 ( .A(n53), .ZN(Y[36]) );
  AOI222_X1 U76 ( .A1(mask00[36]), .A2(n100), .B1(mask16[36]), .B2(n94), .C1(
        mask08[36]), .C2(n88), .ZN(n53) );
  BUF_X1 U77 ( .A(n42), .Z(n96) );
  BUF_X1 U78 ( .A(n43), .Z(n90) );
  BUF_X1 U79 ( .A(n44), .Z(n84) );
  BUF_X1 U80 ( .A(n42), .Z(n97) );
  BUF_X1 U81 ( .A(n43), .Z(n91) );
  BUF_X1 U82 ( .A(n44), .Z(n85) );
  AOI222_X1 U83 ( .A1(mask00[38]), .A2(n100), .B1(mask16[38]), .B2(n94), .C1(
        mask08[38]), .C2(n88), .ZN(n51) );
  AOI222_X1 U84 ( .A1(mask00[1]), .A2(n98), .B1(mask16[1]), .B2(n92), .C1(
        mask08[1]), .C2(n86), .ZN(n71) );
  AOI222_X1 U85 ( .A1(mask00[0]), .A2(n98), .B1(mask16[0]), .B2(n92), .C1(
        mask08[0]), .C2(n86), .ZN(n82) );
  INV_X1 U86 ( .A(n47), .ZN(Y[6]) );
  AOI222_X1 U87 ( .A1(mask00[6]), .A2(n100), .B1(mask16[6]), .B2(n94), .C1(
        mask08[6]), .C2(n88), .ZN(n47) );
  INV_X1 U88 ( .A(n46), .ZN(Y[7]) );
  AOI222_X1 U89 ( .A1(mask00[7]), .A2(n101), .B1(mask16[7]), .B2(n95), .C1(
        mask08[7]), .C2(n89), .ZN(n46) );
  NOR2_X1 U90 ( .A1(sel[0]), .A2(sel[1]), .ZN(n42) );
  NOR2_X1 U91 ( .A1(n83), .A2(sel[0]), .ZN(n43) );
  INV_X1 U92 ( .A(n49), .ZN(Y[4]) );
  AOI222_X1 U93 ( .A1(mask00[4]), .A2(n100), .B1(mask16[4]), .B2(n94), .C1(
        mask08[4]), .C2(n88), .ZN(n49) );
  INV_X1 U94 ( .A(n48), .ZN(Y[5]) );
  AOI222_X1 U95 ( .A1(mask00[5]), .A2(n100), .B1(mask16[5]), .B2(n94), .C1(
        mask08[5]), .C2(n88), .ZN(n48) );
  INV_X1 U96 ( .A(n60), .ZN(Y[2]) );
  AOI222_X1 U97 ( .A1(mask00[2]), .A2(n99), .B1(mask16[2]), .B2(n93), .C1(
        mask08[2]), .C2(n87), .ZN(n60) );
  INV_X1 U98 ( .A(n50), .ZN(Y[3]) );
  AOI222_X1 U99 ( .A1(mask00[3]), .A2(n100), .B1(mask16[3]), .B2(n94), .C1(
        mask08[3]), .C2(n88), .ZN(n50) );
  INV_X1 U100 ( .A(sel[1]), .ZN(n83) );
  AND2_X1 U101 ( .A1(sel[0]), .A2(n83), .ZN(n44) );
endmodule


module shift_firstLevel ( A, sel, mask00, mask08, mask16 );
  input [31:0] A;
  input [1:0] sel;
  output [38:0] mask00;
  output [38:0] mask08;
  output [38:0] mask16;
  wire   n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n98, n116, n117,
         \mask16[22] , n119, n120, n121;
  assign mask08[30] = mask16[38];
  assign mask08[29] = mask16[37];
  assign mask08[28] = mask16[36];
  assign mask08[27] = mask16[35];
  assign mask08[26] = mask16[34];
  assign mask08[25] = mask16[33];
  assign mask08[24] = mask16[32];
  assign mask08[14] = mask16[6];
  assign mask08[13] = mask16[5];
  assign mask08[12] = mask16[4];
  assign mask08[11] = mask16[3];
  assign mask08[10] = mask16[2];
  assign mask08[9] = mask16[1];
  assign mask08[8] = mask16[0];
  assign mask16[18] = \mask16[22] ;
  assign mask16[17] = \mask16[22] ;
  assign mask16[21] = \mask16[22] ;
  assign mask16[20] = \mask16[22] ;
  assign mask16[19] = \mask16[22] ;
  assign mask16[16] = \mask16[22] ;
  assign mask16[22] = \mask16[22] ;

  NAND3_X1 U161 ( .A1(sel[1]), .A2(n108), .A3(A[31]), .ZN(n61) );
  INV_X1 U2 ( .A(n116), .ZN(n98) );
  INV_X1 U3 ( .A(\mask16[22] ), .ZN(n117) );
  BUF_X1 U4 ( .A(n59), .Z(n121) );
  BUF_X1 U5 ( .A(n59), .Z(n120) );
  BUF_X1 U6 ( .A(n59), .Z(n119) );
  INV_X1 U7 ( .A(mask16[7]), .ZN(n94) );
  INV_X1 U8 ( .A(mask08[6]), .ZN(n111) );
  INV_X1 U9 ( .A(mask08[1]), .ZN(n96) );
  INV_X1 U10 ( .A(mask08[5]), .ZN(n112) );
  INV_X1 U11 ( .A(mask08[4]), .ZN(n113) );
  INV_X1 U12 ( .A(mask08[3]), .ZN(n114) );
  INV_X1 U13 ( .A(mask08[2]), .ZN(n115) );
  OAI21_X1 U14 ( .B1(n120), .B2(n60), .A(n117), .ZN(mask16[38]) );
  OAI21_X1 U15 ( .B1(n120), .B2(n63), .A(n117), .ZN(mask16[36]) );
  OAI21_X1 U16 ( .B1(n120), .B2(n64), .A(n117), .ZN(mask16[35]) );
  OAI21_X1 U17 ( .B1(n120), .B2(n65), .A(n117), .ZN(mask16[34]) );
  OAI21_X1 U18 ( .B1(n120), .B2(n66), .A(n117), .ZN(mask16[33]) );
  OAI21_X1 U19 ( .B1(n120), .B2(n67), .A(n117), .ZN(mask16[32]) );
  OAI21_X1 U20 ( .B1(n120), .B2(n62), .A(n117), .ZN(mask16[37]) );
  NOR2_X1 U21 ( .A1(n86), .A2(n116), .ZN(mask16[7]) );
  NOR2_X1 U22 ( .A1(n60), .A2(n116), .ZN(mask08[7]) );
  NOR2_X1 U23 ( .A1(n62), .A2(n116), .ZN(mask08[6]) );
  NOR2_X1 U24 ( .A1(n67), .A2(n116), .ZN(mask08[1]) );
  NOR2_X1 U25 ( .A1(n65), .A2(n116), .ZN(mask08[3]) );
  NOR2_X1 U26 ( .A1(n66), .A2(n116), .ZN(mask08[2]) );
  NOR2_X1 U27 ( .A1(n63), .A2(n116), .ZN(mask08[5]) );
  NOR2_X1 U28 ( .A1(n64), .A2(n116), .ZN(mask08[4]) );
  INV_X1 U29 ( .A(n61), .ZN(\mask16[22] ) );
  INV_X1 U30 ( .A(n53), .ZN(mask16[9]) );
  NAND2_X1 U31 ( .A1(n96), .A2(n75), .ZN(mask00[9]) );
  INV_X1 U32 ( .A(n54), .ZN(mask16[8]) );
  NAND2_X1 U33 ( .A1(n95), .A2(n76), .ZN(mask00[8]) );
  INV_X1 U34 ( .A(n83), .ZN(mask16[11]) );
  NAND2_X1 U35 ( .A1(n114), .A2(n73), .ZN(mask00[11]) );
  INV_X1 U36 ( .A(n84), .ZN(mask16[10]) );
  NAND2_X1 U37 ( .A1(n115), .A2(n74), .ZN(mask00[10]) );
  OAI21_X1 U38 ( .B1(n121), .B2(n93), .A(n94), .ZN(mask00[23]) );
  OAI21_X1 U39 ( .B1(n87), .B2(n119), .A(n117), .ZN(mask08[37]) );
  INV_X1 U40 ( .A(n97), .ZN(n59) );
  NAND2_X1 U41 ( .A1(n61), .A2(n69), .ZN(mask16[30]) );
  OAI21_X1 U42 ( .B1(n86), .B2(n119), .A(n80), .ZN(mask00[30]) );
  NAND2_X1 U43 ( .A1(n61), .A2(n71), .ZN(mask16[29]) );
  OAI21_X1 U44 ( .B1(n87), .B2(n119), .A(n81), .ZN(mask00[29]) );
  NAND2_X1 U45 ( .A1(n61), .A2(n72), .ZN(mask16[28]) );
  OAI21_X1 U46 ( .B1(n88), .B2(n119), .A(n82), .ZN(mask00[28]) );
  NAND2_X1 U47 ( .A1(n61), .A2(n73), .ZN(mask16[27]) );
  OAI21_X1 U48 ( .B1(n89), .B2(n119), .A(n83), .ZN(mask00[27]) );
  NAND2_X1 U49 ( .A1(n61), .A2(n74), .ZN(mask16[26]) );
  OAI21_X1 U50 ( .B1(n90), .B2(n119), .A(n84), .ZN(mask00[26]) );
  NAND2_X1 U51 ( .A1(n61), .A2(n75), .ZN(mask16[25]) );
  OAI21_X1 U52 ( .B1(n121), .B2(n91), .A(n53), .ZN(mask00[25]) );
  NAND2_X1 U53 ( .A1(n117), .A2(n76), .ZN(mask16[24]) );
  OAI21_X1 U54 ( .B1(n121), .B2(n92), .A(n54), .ZN(mask00[24]) );
  NAND2_X1 U55 ( .A1(n79), .A2(n68), .ZN(mask08[23]) );
  NAND2_X1 U56 ( .A1(n61), .A2(n77), .ZN(mask16[23]) );
  NAND2_X1 U57 ( .A1(n80), .A2(n69), .ZN(mask08[22]) );
  OAI21_X1 U58 ( .B1(n121), .B2(n60), .A(n55), .ZN(mask00[22]) );
  NAND2_X1 U59 ( .A1(n81), .A2(n71), .ZN(mask08[21]) );
  OAI21_X1 U60 ( .B1(n121), .B2(n62), .A(n56), .ZN(mask00[21]) );
  NAND2_X1 U61 ( .A1(n82), .A2(n72), .ZN(mask08[20]) );
  OAI21_X1 U62 ( .B1(n121), .B2(n63), .A(n57), .ZN(mask00[20]) );
  NAND2_X1 U63 ( .A1(n83), .A2(n73), .ZN(mask08[19]) );
  OAI21_X1 U64 ( .B1(n121), .B2(n64), .A(n58), .ZN(mask00[19]) );
  NAND2_X1 U65 ( .A1(n84), .A2(n74), .ZN(mask08[18]) );
  OAI21_X1 U66 ( .B1(n121), .B2(n65), .A(n70), .ZN(mask00[18]) );
  NAND2_X1 U67 ( .A1(n53), .A2(n75), .ZN(mask08[17]) );
  OAI21_X1 U68 ( .B1(n121), .B2(n66), .A(n78), .ZN(mask00[17]) );
  NAND2_X1 U69 ( .A1(n54), .A2(n76), .ZN(mask08[16]) );
  OAI21_X1 U70 ( .B1(n120), .B2(n67), .A(n85), .ZN(mask00[16]) );
  INV_X1 U71 ( .A(n79), .ZN(mask16[15]) );
  NAND2_X1 U72 ( .A1(n94), .A2(n77), .ZN(mask08[15]) );
  INV_X1 U73 ( .A(n80), .ZN(mask16[14]) );
  NAND2_X1 U74 ( .A1(n111), .A2(n69), .ZN(mask00[14]) );
  INV_X1 U75 ( .A(n81), .ZN(mask16[13]) );
  NAND2_X1 U76 ( .A1(n112), .A2(n71), .ZN(mask00[13]) );
  INV_X1 U77 ( .A(n82), .ZN(mask16[12]) );
  NAND2_X1 U78 ( .A1(n113), .A2(n72), .ZN(mask00[12]) );
  OAI21_X1 U79 ( .B1(n120), .B2(n91), .A(n61), .ZN(mask08[33]) );
  OAI21_X1 U80 ( .B1(n90), .B2(n119), .A(n117), .ZN(mask08[34]) );
  OAI21_X1 U81 ( .B1(n89), .B2(n119), .A(n117), .ZN(mask08[35]) );
  OAI21_X1 U82 ( .B1(n121), .B2(n104), .A(n61), .ZN(mask00[35]) );
  OAI21_X1 U83 ( .B1(n120), .B2(n92), .A(n117), .ZN(mask08[32]) );
  OAI21_X1 U84 ( .B1(n107), .B2(n119), .A(n117), .ZN(mask00[32]) );
  NAND2_X1 U85 ( .A1(n61), .A2(n68), .ZN(mask16[31]) );
  OAI21_X1 U86 ( .B1(n120), .B2(n93), .A(n61), .ZN(mask08[31]) );
  OAI21_X1 U87 ( .B1(n88), .B2(n119), .A(n117), .ZN(mask08[36]) );
  OAI21_X1 U88 ( .B1(n121), .B2(n103), .A(n117), .ZN(mask00[36]) );
  INV_X1 U89 ( .A(n55), .ZN(mask16[6]) );
  INV_X1 U90 ( .A(n56), .ZN(mask16[5]) );
  INV_X1 U91 ( .A(n57), .ZN(mask16[4]) );
  INV_X1 U92 ( .A(n58), .ZN(mask16[3]) );
  INV_X1 U93 ( .A(n78), .ZN(mask16[1]) );
  INV_X1 U94 ( .A(n85), .ZN(mask16[0]) );
  INV_X1 U95 ( .A(n70), .ZN(mask16[2]) );
  NAND2_X1 U96 ( .A1(n110), .A2(n68), .ZN(mask00[15]) );
  INV_X1 U97 ( .A(mask08[7]), .ZN(n110) );
  NOR2_X1 U98 ( .A1(sel[0]), .A2(sel[1]), .ZN(n97) );
  OAI21_X1 U99 ( .B1(n86), .B2(n119), .A(n117), .ZN(mask08[38]) );
  OAI21_X1 U100 ( .B1(n120), .B2(n101), .A(n61), .ZN(mask00[38]) );
  INV_X1 U101 ( .A(A[31]), .ZN(n101) );
  AND2_X1 U102 ( .A1(n99), .A2(A[1]), .ZN(mask00[1]) );
  INV_X1 U103 ( .A(n95), .ZN(mask08[0]) );
  AND2_X1 U104 ( .A1(n99), .A2(A[0]), .ZN(mask00[0]) );
  INV_X1 U105 ( .A(sel[0]), .ZN(n108) );
  AOI21_X1 U106 ( .B1(sel[0]), .B2(sel[1]), .A(n97), .ZN(n99) );
  NAND2_X1 U107 ( .A1(A[8]), .A2(n97), .ZN(n68) );
  NAND2_X1 U108 ( .A1(A[7]), .A2(n97), .ZN(n69) );
  NAND2_X1 U109 ( .A1(A[2]), .A2(n97), .ZN(n75) );
  NAND2_X1 U110 ( .A1(A[1]), .A2(n97), .ZN(n76) );
  NAND2_X1 U111 ( .A1(A[6]), .A2(n97), .ZN(n71) );
  NAND2_X1 U112 ( .A1(A[5]), .A2(n97), .ZN(n72) );
  NAND2_X1 U113 ( .A1(A[4]), .A2(n97), .ZN(n73) );
  NAND2_X1 U114 ( .A1(A[3]), .A2(n97), .ZN(n74) );
  AND2_X1 U115 ( .A1(n99), .A2(A[6]), .ZN(mask00[6]) );
  NAND2_X1 U116 ( .A1(A[0]), .A2(n97), .ZN(n77) );
  OAI21_X1 U117 ( .B1(n116), .B2(n100), .A(n77), .ZN(mask00[7]) );
  INV_X1 U118 ( .A(A[7]), .ZN(n100) );
  NAND2_X1 U119 ( .A1(A[31]), .A2(n98), .ZN(n79) );
  NAND2_X1 U120 ( .A1(A[30]), .A2(n98), .ZN(n80) );
  NAND2_X1 U121 ( .A1(A[25]), .A2(n98), .ZN(n53) );
  NAND2_X1 U122 ( .A1(A[24]), .A2(n98), .ZN(n54) );
  NAND2_X1 U123 ( .A1(A[29]), .A2(n98), .ZN(n81) );
  NAND2_X1 U124 ( .A1(A[28]), .A2(n98), .ZN(n82) );
  NAND2_X1 U125 ( .A1(A[27]), .A2(n98), .ZN(n83) );
  NAND2_X1 U126 ( .A1(A[26]), .A2(n98), .ZN(n84) );
  OAI21_X1 U127 ( .B1(n109), .B2(n119), .A(n79), .ZN(mask00[31]) );
  INV_X1 U128 ( .A(A[24]), .ZN(n109) );
  OAI21_X1 U129 ( .B1(n121), .B2(n105), .A(n61), .ZN(mask00[34]) );
  INV_X1 U130 ( .A(A[27]), .ZN(n105) );
  OAI21_X1 U131 ( .B1(n121), .B2(n106), .A(n61), .ZN(mask00[33]) );
  INV_X1 U132 ( .A(A[26]), .ZN(n106) );
  OAI21_X1 U133 ( .B1(n120), .B2(n102), .A(n61), .ZN(mask00[37]) );
  INV_X1 U134 ( .A(A[30]), .ZN(n102) );
  NAND2_X1 U135 ( .A1(A[21]), .A2(n98), .ZN(n56) );
  NAND2_X1 U136 ( .A1(A[20]), .A2(n98), .ZN(n57) );
  NAND2_X1 U137 ( .A1(A[19]), .A2(n98), .ZN(n58) );
  NAND2_X1 U138 ( .A1(A[22]), .A2(n98), .ZN(n55) );
  AND2_X1 U139 ( .A1(n99), .A2(A[4]), .ZN(mask00[4]) );
  AND2_X1 U140 ( .A1(n99), .A2(A[5]), .ZN(mask00[5]) );
  INV_X1 U141 ( .A(A[15]), .ZN(n60) );
  INV_X1 U142 ( .A(A[14]), .ZN(n62) );
  INV_X1 U143 ( .A(A[9]), .ZN(n67) );
  INV_X1 U144 ( .A(A[11]), .ZN(n65) );
  INV_X1 U145 ( .A(A[10]), .ZN(n66) );
  INV_X1 U146 ( .A(A[13]), .ZN(n63) );
  INV_X1 U147 ( .A(A[12]), .ZN(n64) );
  INV_X1 U148 ( .A(A[23]), .ZN(n86) );
  NAND2_X1 U149 ( .A1(A[18]), .A2(n99), .ZN(n70) );
  NAND2_X1 U150 ( .A1(A[17]), .A2(n99), .ZN(n78) );
  NAND2_X1 U151 ( .A1(A[16]), .A2(n99), .ZN(n85) );
  NAND2_X1 U152 ( .A1(A[8]), .A2(n99), .ZN(n95) );
  AND2_X1 U153 ( .A1(n99), .A2(A[2]), .ZN(mask00[2]) );
  AND2_X1 U154 ( .A1(n99), .A2(A[3]), .ZN(mask00[3]) );
  INV_X1 U155 ( .A(A[18]), .ZN(n91) );
  INV_X1 U156 ( .A(A[17]), .ZN(n92) );
  INV_X1 U157 ( .A(A[16]), .ZN(n93) );
  INV_X1 U158 ( .A(A[22]), .ZN(n87) );
  INV_X1 U159 ( .A(A[21]), .ZN(n88) );
  INV_X1 U160 ( .A(A[20]), .ZN(n89) );
  INV_X1 U162 ( .A(A[19]), .ZN(n90) );
  INV_X1 U163 ( .A(A[29]), .ZN(n103) );
  INV_X1 U164 ( .A(A[28]), .ZN(n104) );
  INV_X1 U165 ( .A(A[25]), .ZN(n107) );
  INV_X1 U166 ( .A(n99), .ZN(n116) );
endmodule


module cla_adder_N32_1 ( A, B, Ci, Cout, Sum );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Ci;
  output Cout;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50;
  wire   [8:0] Carry;
  assign n3 = A[5];
  assign n4 = B[6];
  assign n5 = A[2];
  assign n6 = A[12];
  assign n7 = A[0];
  assign n8 = B[10];
  assign n9 = B[26];
  assign n10 = B[5];
  assign n11 = B[22];
  assign n12 = B[3];
  assign n13 = A[1];
  assign n14 = A[6];
  assign n15 = A[18];
  assign n16 = A[7];
  assign n17 = B[7];
  assign n18 = B[11];
  assign n19 = A[19];
  assign n20 = A[3];
  assign n21 = B[9];
  assign n22 = A[29];
  assign n23 = B[12];
  assign n24 = A[10];
  assign n25 = B[18];
  assign n26 = B[14];
  assign n27 = A[11];
  assign n28 = A[22];
  assign n29 = B[19];
  assign n30 = A[17];
  assign n31 = B[15];
  assign n32 = A[9];
  assign n33 = B[17];
  assign n34 = A[25];
  assign n35 = A[26];
  assign n36 = B[29];
  assign n37 = A[21];
  assign n38 = B[13];
  assign n39 = A[13];
  assign n40 = A[14];
  assign n41 = A[15];
  assign n42 = B[24];
  assign n43 = B[27];
  assign n44 = B[28];
  assign n45 = A[27];
  assign n46 = B[21];
  assign n47 = A[28];
  assign n48 = A[24];
  assign n49 = B[23];
  assign n50 = A[23];

  carry_generator_N32_Nblocks8_1 CG ( .A({A[31:30], n22, n47, n45, n35, n34, 
        n48, n50, n28, n37, A[20], n19, n15, n30, A[16], n41, n40, n39, n6, 
        n27, n24, n32, A[8], n16, n14, n3, A[4], n20, n5, n13, n7}), .B({
        B[31:30], n36, n44, n43, n9, B[25], n42, n49, n11, n46, B[20], n29, 
        n25, n33, B[16], n31, n26, n38, n23, n18, n8, n21, B[8], n17, n4, n10, 
        B[4], n12, B[2:0]}), .Ci(Ci), .Cout(Carry) );
  sum_generator_Nbits32_Nblocks8_1 SG ( .A({A[31:30], n22, n47, n45, n35, n34, 
        n48, n50, n28, n37, A[20], n19, n15, n30, A[16], n41, n40, n39, n6, 
        n27, n24, n32, A[8], n16, n14, n3, A[4], n20, n5, n13, n7}), .B({
        B[31:30], n36, n44, n43, n9, B[25], n42, n49, n11, n46, B[20], n29, 
        n25, n33, B[16], n31, n26, n38, n23, n18, n8, n21, B[8], n17, n4, n10, 
        B[4], n12, B[2:0]}), .Carry(Carry), .S(Sum), .Cout(Cout) );
endmodule


module CSA_Nbits32_1 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_96 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_95 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_94 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_93 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_92 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_91 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_90 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_89 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_88 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_87 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_86 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(Cout[11]) );
  FA_85 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(Cout[12]) );
  FA_84 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(Cout[13]) );
  FA_83 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(Cout[14]) );
  FA_82 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(Cout[15]) );
  FA_81 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(Cout[16]) );
  FA_80 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(Cout[17]) );
  FA_79 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(Cout[18]) );
  FA_78 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(Cout[19]) );
  FA_77 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(Cout[20]) );
  FA_76 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(Cout[21]) );
  FA_75 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(Cout[22]) );
  FA_74 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(Cout[23]) );
  FA_73 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(Cout[24]) );
  FA_72 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(Cout[25]) );
  FA_71 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(Cout[26]) );
  FA_70 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(Cout[27]) );
  FA_69 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(Cout[28]) );
  FA_68 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(Cout[29]) );
  FA_67 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(Cout[30]) );
  FA_66 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(Cout[31]) );
  FA_65 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module CSA_Nbits32_2 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_128 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_127 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_126 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_125 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_124 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_123 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_122 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_121 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_120 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_119 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_118 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(
        Cout[11]) );
  FA_117 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(
        Cout[12]) );
  FA_116 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(
        Cout[13]) );
  FA_115 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(
        Cout[14]) );
  FA_114 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(
        Cout[15]) );
  FA_113 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(
        Cout[16]) );
  FA_112 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(
        Cout[17]) );
  FA_111 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(
        Cout[18]) );
  FA_110 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(
        Cout[19]) );
  FA_109 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(
        Cout[20]) );
  FA_108 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(
        Cout[21]) );
  FA_107 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(
        Cout[22]) );
  FA_106 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(
        Cout[23]) );
  FA_105 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(
        Cout[24]) );
  FA_104 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(
        Cout[25]) );
  FA_103 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(
        Cout[26]) );
  FA_102 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(
        Cout[27]) );
  FA_101 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(
        Cout[28]) );
  FA_100 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(
        Cout[29]) );
  FA_99 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(Cout[30]) );
  FA_98 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(Cout[31]) );
  FA_97 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module CSA_Nbits32_3 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_160 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_159 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_158 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_157 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_156 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_155 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_154 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_153 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_152 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_151 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_150 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(
        Cout[11]) );
  FA_149 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(
        Cout[12]) );
  FA_148 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(
        Cout[13]) );
  FA_147 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(
        Cout[14]) );
  FA_146 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(
        Cout[15]) );
  FA_145 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(
        Cout[16]) );
  FA_144 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(
        Cout[17]) );
  FA_143 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(
        Cout[18]) );
  FA_142 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(
        Cout[19]) );
  FA_141 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(
        Cout[20]) );
  FA_140 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(
        Cout[21]) );
  FA_139 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(
        Cout[22]) );
  FA_138 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(
        Cout[23]) );
  FA_137 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(
        Cout[24]) );
  FA_136 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(
        Cout[25]) );
  FA_135 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(
        Cout[26]) );
  FA_134 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(
        Cout[27]) );
  FA_133 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(
        Cout[28]) );
  FA_132 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(
        Cout[29]) );
  FA_131 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(
        Cout[30]) );
  FA_130 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(
        Cout[31]) );
  FA_129 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module CSA_Nbits32_4 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_192 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_191 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_190 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_189 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_188 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_187 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_186 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_185 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_184 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_183 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_182 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(
        Cout[11]) );
  FA_181 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(
        Cout[12]) );
  FA_180 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(
        Cout[13]) );
  FA_179 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(
        Cout[14]) );
  FA_178 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(
        Cout[15]) );
  FA_177 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(
        Cout[16]) );
  FA_176 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(
        Cout[17]) );
  FA_175 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(
        Cout[18]) );
  FA_174 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(
        Cout[19]) );
  FA_173 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(
        Cout[20]) );
  FA_172 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(
        Cout[21]) );
  FA_171 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(
        Cout[22]) );
  FA_170 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(
        Cout[23]) );
  FA_169 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(
        Cout[24]) );
  FA_168 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(
        Cout[25]) );
  FA_167 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(
        Cout[26]) );
  FA_166 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(
        Cout[27]) );
  FA_165 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(
        Cout[28]) );
  FA_164 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(
        Cout[29]) );
  FA_163 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(
        Cout[30]) );
  FA_162 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(
        Cout[31]) );
  FA_161 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module CSA_Nbits32_5 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_224 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_223 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_222 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_221 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_220 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_219 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_218 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_217 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_216 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_215 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_214 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(
        Cout[11]) );
  FA_213 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(
        Cout[12]) );
  FA_212 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(
        Cout[13]) );
  FA_211 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(
        Cout[14]) );
  FA_210 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(
        Cout[15]) );
  FA_209 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(
        Cout[16]) );
  FA_208 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(
        Cout[17]) );
  FA_207 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(
        Cout[18]) );
  FA_206 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(
        Cout[19]) );
  FA_205 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(
        Cout[20]) );
  FA_204 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(
        Cout[21]) );
  FA_203 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(
        Cout[22]) );
  FA_202 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(
        Cout[23]) );
  FA_201 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(
        Cout[24]) );
  FA_200 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(
        Cout[25]) );
  FA_199 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(
        Cout[26]) );
  FA_198 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(
        Cout[27]) );
  FA_197 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(
        Cout[28]) );
  FA_196 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(
        Cout[29]) );
  FA_195 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(
        Cout[30]) );
  FA_194 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(
        Cout[31]) );
  FA_193 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module CSA_Nbits32_0 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] S;
  output [31:0] Cout;

  assign Cout[0] = 1'b0;

  FA_64 FullAdd_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(S[0]), .Co(Cout[1]) );
  FA_255 FullAdd_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(S[1]), .Co(Cout[2]) );
  FA_254 FullAdd_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(S[2]), .Co(Cout[3]) );
  FA_253 FullAdd_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(S[3]), .Co(Cout[4]) );
  FA_252 FullAdd_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(S[4]), .Co(Cout[5]) );
  FA_251 FullAdd_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(S[5]), .Co(Cout[6]) );
  FA_250 FullAdd_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(S[6]), .Co(Cout[7]) );
  FA_249 FullAdd_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(S[7]), .Co(Cout[8]) );
  FA_248 FullAdd_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(S[8]), .Co(Cout[9]) );
  FA_247 FullAdd_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(S[9]), .Co(Cout[10]) );
  FA_246 FullAdd_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(S[10]), .Co(
        Cout[11]) );
  FA_245 FullAdd_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(S[11]), .Co(
        Cout[12]) );
  FA_244 FullAdd_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(S[12]), .Co(
        Cout[13]) );
  FA_243 FullAdd_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(S[13]), .Co(
        Cout[14]) );
  FA_242 FullAdd_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(S[14]), .Co(
        Cout[15]) );
  FA_241 FullAdd_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(S[15]), .Co(
        Cout[16]) );
  FA_240 FullAdd_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(S[16]), .Co(
        Cout[17]) );
  FA_239 FullAdd_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(S[17]), .Co(
        Cout[18]) );
  FA_238 FullAdd_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(S[18]), .Co(
        Cout[19]) );
  FA_237 FullAdd_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(S[19]), .Co(
        Cout[20]) );
  FA_236 FullAdd_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(S[20]), .Co(
        Cout[21]) );
  FA_235 FullAdd_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(S[21]), .Co(
        Cout[22]) );
  FA_234 FullAdd_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(S[22]), .Co(
        Cout[23]) );
  FA_233 FullAdd_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(S[23]), .Co(
        Cout[24]) );
  FA_232 FullAdd_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(S[24]), .Co(
        Cout[25]) );
  FA_231 FullAdd_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(S[25]), .Co(
        Cout[26]) );
  FA_230 FullAdd_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(S[26]), .Co(
        Cout[27]) );
  FA_229 FullAdd_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(S[27]), .Co(
        Cout[28]) );
  FA_228 FullAdd_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(S[28]), .Co(
        Cout[29]) );
  FA_227 FullAdd_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(S[29]), .Co(
        Cout[30]) );
  FA_226 FullAdd_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(S[30]), .Co(
        Cout[31]) );
  FA_225 LastFA ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(S[31]) );
endmodule


module mux_N32_1 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270;

  BUF_X1 U1 ( .A(n10), .Z(n257) );
  BUF_X1 U2 ( .A(n10), .Z(n256) );
  BUF_X1 U3 ( .A(n10), .Z(n258) );
  BUF_X1 U4 ( .A(n6), .Z(n269) );
  BUF_X1 U5 ( .A(n6), .Z(n268) );
  BUF_X1 U6 ( .A(n9), .Z(n260) );
  BUF_X1 U7 ( .A(n9), .Z(n259) );
  BUF_X1 U8 ( .A(n7), .Z(n266) );
  BUF_X1 U9 ( .A(n7), .Z(n265) );
  BUF_X1 U10 ( .A(n8), .Z(n263) );
  BUF_X1 U11 ( .A(n8), .Z(n262) );
  BUF_X1 U12 ( .A(n9), .Z(n261) );
  BUF_X1 U13 ( .A(n7), .Z(n267) );
  BUF_X1 U14 ( .A(n8), .Z(n264) );
  BUF_X1 U15 ( .A(n6), .Z(n270) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  NAND2_X1 U22 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U23 ( .A1(A[28]), .A2(n260), .B1(B[28]), .B2(n257), .ZN(n31) );
  AOI222_X1 U24 ( .A1(D[28]), .A2(n269), .B1(E[28]), .B2(n266), .C1(C[28]), 
        .C2(n263), .ZN(n32) );
  NAND2_X1 U25 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U26 ( .A1(A[14]), .A2(n259), .B1(B[14]), .B2(n256), .ZN(n61) );
  AOI222_X1 U27 ( .A1(D[14]), .A2(n268), .B1(E[14]), .B2(n265), .C1(C[14]), 
        .C2(n262), .ZN(n62) );
  NAND2_X1 U28 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U29 ( .A1(A[24]), .A2(n260), .B1(B[24]), .B2(n257), .ZN(n39) );
  AOI222_X1 U30 ( .A1(D[24]), .A2(n269), .B1(E[24]), .B2(n266), .C1(C[24]), 
        .C2(n263), .ZN(n40) );
  NAND2_X1 U31 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U32 ( .A1(A[18]), .A2(n259), .B1(B[18]), .B2(n256), .ZN(n53) );
  AOI222_X1 U33 ( .A1(D[18]), .A2(n268), .B1(E[18]), .B2(n265), .C1(C[18]), 
        .C2(n262), .ZN(n54) );
  NAND2_X1 U34 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U35 ( .A1(A[15]), .A2(n259), .B1(B[15]), .B2(n256), .ZN(n59) );
  AOI222_X1 U36 ( .A1(D[15]), .A2(n268), .B1(E[15]), .B2(n265), .C1(C[15]), 
        .C2(n262), .ZN(n60) );
  NAND2_X1 U37 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U38 ( .A1(A[22]), .A2(n260), .B1(B[22]), .B2(n257), .ZN(n43) );
  AOI222_X1 U39 ( .A1(D[22]), .A2(n269), .B1(E[22]), .B2(n266), .C1(C[22]), 
        .C2(n263), .ZN(n44) );
  NAND2_X1 U40 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U41 ( .A1(A[16]), .A2(n259), .B1(B[16]), .B2(n256), .ZN(n57) );
  AOI222_X1 U42 ( .A1(D[16]), .A2(n268), .B1(E[16]), .B2(n265), .C1(C[16]), 
        .C2(n262), .ZN(n58) );
  NAND2_X1 U43 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U44 ( .A1(A[20]), .A2(n260), .B1(B[20]), .B2(n257), .ZN(n47) );
  AOI222_X1 U45 ( .A1(D[20]), .A2(n269), .B1(E[20]), .B2(n266), .C1(C[20]), 
        .C2(n263), .ZN(n48) );
  NAND2_X1 U46 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U47 ( .A1(A[27]), .A2(n260), .B1(B[27]), .B2(n257), .ZN(n33) );
  AOI222_X1 U48 ( .A1(D[27]), .A2(n269), .B1(E[27]), .B2(n266), .C1(C[27]), 
        .C2(n263), .ZN(n34) );
  NAND2_X1 U49 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U50 ( .A1(A[23]), .A2(n260), .B1(B[23]), .B2(n257), .ZN(n41) );
  AOI222_X1 U51 ( .A1(D[23]), .A2(n269), .B1(E[23]), .B2(n266), .C1(C[23]), 
        .C2(n263), .ZN(n42) );
  NAND2_X1 U52 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U53 ( .A1(A[17]), .A2(n259), .B1(B[17]), .B2(n256), .ZN(n55) );
  AOI222_X1 U54 ( .A1(D[17]), .A2(n268), .B1(E[17]), .B2(n265), .C1(C[17]), 
        .C2(n262), .ZN(n56) );
  NAND2_X1 U55 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U56 ( .A1(A[21]), .A2(n260), .B1(B[21]), .B2(n257), .ZN(n45) );
  AOI222_X1 U57 ( .A1(D[21]), .A2(n269), .B1(E[21]), .B2(n266), .C1(C[21]), 
        .C2(n263), .ZN(n46) );
  NAND2_X1 U58 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U59 ( .A1(A[19]), .A2(n259), .B1(B[19]), .B2(n256), .ZN(n51) );
  AOI222_X1 U60 ( .A1(D[19]), .A2(n268), .B1(E[19]), .B2(n265), .C1(C[19]), 
        .C2(n262), .ZN(n52) );
  AND2_X1 U61 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U62 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U63 ( .A1(A[25]), .A2(n260), .B1(B[25]), .B2(n257), .ZN(n37) );
  AOI222_X1 U64 ( .A1(D[25]), .A2(n269), .B1(E[25]), .B2(n266), .C1(C[25]), 
        .C2(n263), .ZN(n38) );
  NAND2_X1 U65 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U66 ( .A1(A[29]), .A2(n260), .B1(B[29]), .B2(n257), .ZN(n29) );
  AOI222_X1 U67 ( .A1(D[29]), .A2(n269), .B1(E[29]), .B2(n266), .C1(C[29]), 
        .C2(n263), .ZN(n30) );
  INV_X1 U68 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U69 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U70 ( .A1(A[26]), .A2(n260), .B1(B[26]), .B2(n257), .ZN(n35) );
  AOI222_X1 U71 ( .A1(D[26]), .A2(n269), .B1(E[26]), .B2(n266), .C1(C[26]), 
        .C2(n263), .ZN(n36) );
  NAND2_X1 U72 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U73 ( .A1(A[6]), .A2(n261), .B1(B[6]), .B2(n258), .ZN(n15) );
  AOI222_X1 U74 ( .A1(D[6]), .A2(n270), .B1(E[6]), .B2(n267), .C1(C[6]), .C2(
        n264), .ZN(n16) );
  NAND2_X1 U75 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U76 ( .A1(A[3]), .A2(n261), .B1(B[3]), .B2(n258), .ZN(n21) );
  AOI222_X1 U77 ( .A1(D[3]), .A2(n270), .B1(E[3]), .B2(n267), .C1(C[3]), .C2(
        n264), .ZN(n22) );
  NAND2_X1 U78 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U79 ( .A1(A[7]), .A2(n261), .B1(B[7]), .B2(n258), .ZN(n13) );
  AOI222_X1 U80 ( .A1(D[7]), .A2(n270), .B1(E[7]), .B2(n267), .C1(C[7]), .C2(
        n264), .ZN(n14) );
  NAND2_X1 U81 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U82 ( .A1(A[4]), .A2(n261), .B1(B[4]), .B2(n258), .ZN(n19) );
  AOI222_X1 U83 ( .A1(D[4]), .A2(n270), .B1(E[4]), .B2(n267), .C1(C[4]), .C2(
        n264), .ZN(n20) );
  NAND2_X1 U84 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U85 ( .A1(A[8]), .A2(n261), .B1(B[8]), .B2(n258), .ZN(n11) );
  AOI222_X1 U86 ( .A1(D[8]), .A2(n270), .B1(E[8]), .B2(n267), .C1(C[8]), .C2(
        n264), .ZN(n12) );
  NAND2_X1 U87 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U88 ( .A1(A[9]), .A2(n261), .B1(B[9]), .B2(n258), .ZN(n4) );
  AOI222_X1 U89 ( .A1(D[9]), .A2(n270), .B1(E[9]), .B2(n267), .C1(C[9]), .C2(
        n264), .ZN(n5) );
  NAND2_X1 U90 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U91 ( .A1(A[5]), .A2(n261), .B1(B[5]), .B2(n258), .ZN(n17) );
  AOI222_X1 U92 ( .A1(D[5]), .A2(n270), .B1(E[5]), .B2(n267), .C1(C[5]), .C2(
        n264), .ZN(n18) );
  NAND2_X1 U93 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U94 ( .A1(A[31]), .A2(n261), .B1(B[31]), .B2(n258), .ZN(n23) );
  AOI222_X1 U95 ( .A1(D[31]), .A2(n270), .B1(E[31]), .B2(n267), .C1(C[31]), 
        .C2(n264), .ZN(n24) );
  NAND2_X1 U96 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U97 ( .A1(A[2]), .A2(n260), .B1(B[2]), .B2(n257), .ZN(n27) );
  AOI222_X1 U98 ( .A1(D[2]), .A2(n269), .B1(E[2]), .B2(n266), .C1(C[2]), .C2(
        n263), .ZN(n28) );
  NAND2_X1 U99 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U100 ( .A1(A[10]), .A2(n259), .B1(B[10]), .B2(n256), .ZN(n69) );
  AOI222_X1 U101 ( .A1(D[10]), .A2(n268), .B1(E[10]), .B2(n265), .C1(C[10]), 
        .C2(n262), .ZN(n70) );
  NAND2_X1 U102 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U103 ( .A1(A[11]), .A2(n259), .B1(B[11]), .B2(n256), .ZN(n67) );
  AOI222_X1 U104 ( .A1(D[11]), .A2(n268), .B1(E[11]), .B2(n265), .C1(C[11]), 
        .C2(n262), .ZN(n68) );
  NAND2_X1 U105 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U106 ( .A1(A[0]), .A2(n259), .B1(B[0]), .B2(n256), .ZN(n71) );
  AOI222_X1 U107 ( .A1(D[0]), .A2(n268), .B1(E[0]), .B2(n265), .C1(C[0]), .C2(
        n262), .ZN(n72) );
  NAND2_X1 U108 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U109 ( .A1(A[12]), .A2(n259), .B1(B[12]), .B2(n256), .ZN(n65) );
  AOI222_X1 U110 ( .A1(D[12]), .A2(n268), .B1(E[12]), .B2(n265), .C1(C[12]), 
        .C2(n262), .ZN(n66) );
  NAND2_X1 U111 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U112 ( .A1(A[13]), .A2(n259), .B1(B[13]), .B2(n256), .ZN(n63) );
  AOI222_X1 U113 ( .A1(D[13]), .A2(n268), .B1(E[13]), .B2(n265), .C1(C[13]), 
        .C2(n262), .ZN(n64) );
  NAND2_X1 U114 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U115 ( .A1(A[1]), .A2(n259), .B1(B[1]), .B2(n256), .ZN(n49) );
  AOI222_X1 U116 ( .A1(D[1]), .A2(n268), .B1(E[1]), .B2(n265), .C1(C[1]), .C2(
        n262), .ZN(n50) );
  NAND2_X1 U117 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U118 ( .A1(A[30]), .A2(n260), .B1(B[30]), .B2(n257), .ZN(n25) );
  AOI222_X1 U119 ( .A1(D[30]), .A2(n269), .B1(E[30]), .B2(n266), .C1(C[30]), 
        .C2(n263), .ZN(n26) );
  INV_X1 U120 ( .A(Sel[1]), .ZN(n75) );
endmodule


module mux_N32_2 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282;

  BUF_X1 U1 ( .A(n10), .Z(n269) );
  BUF_X1 U2 ( .A(n10), .Z(n268) );
  BUF_X1 U3 ( .A(n10), .Z(n270) );
  BUF_X1 U4 ( .A(n6), .Z(n281) );
  BUF_X1 U5 ( .A(n6), .Z(n280) );
  BUF_X1 U6 ( .A(n9), .Z(n272) );
  BUF_X1 U7 ( .A(n9), .Z(n271) );
  BUF_X1 U8 ( .A(n7), .Z(n278) );
  BUF_X1 U9 ( .A(n7), .Z(n277) );
  BUF_X1 U10 ( .A(n8), .Z(n275) );
  BUF_X1 U11 ( .A(n8), .Z(n274) );
  BUF_X1 U12 ( .A(n9), .Z(n273) );
  BUF_X1 U13 ( .A(n7), .Z(n279) );
  BUF_X1 U14 ( .A(n8), .Z(n276) );
  BUF_X1 U15 ( .A(n6), .Z(n282) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  INV_X1 U22 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U23 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U24 ( .A1(A[26]), .A2(n272), .B1(B[26]), .B2(n269), .ZN(n35) );
  AOI222_X1 U25 ( .A1(D[26]), .A2(n281), .B1(E[26]), .B2(n278), .C1(C[26]), 
        .C2(n275), .ZN(n36) );
  NAND2_X1 U26 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U27 ( .A1(A[22]), .A2(n272), .B1(B[22]), .B2(n269), .ZN(n43) );
  AOI222_X1 U28 ( .A1(D[22]), .A2(n281), .B1(E[22]), .B2(n278), .C1(C[22]), 
        .C2(n275), .ZN(n44) );
  NAND2_X1 U29 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U30 ( .A1(A[28]), .A2(n272), .B1(B[28]), .B2(n269), .ZN(n31) );
  AOI222_X1 U31 ( .A1(D[28]), .A2(n281), .B1(E[28]), .B2(n278), .C1(C[28]), 
        .C2(n275), .ZN(n32) );
  NAND2_X1 U32 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U33 ( .A1(A[29]), .A2(n272), .B1(B[29]), .B2(n269), .ZN(n29) );
  AOI222_X1 U34 ( .A1(D[29]), .A2(n281), .B1(E[29]), .B2(n278), .C1(C[29]), 
        .C2(n275), .ZN(n30) );
  NAND2_X1 U35 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U36 ( .A1(A[30]), .A2(n272), .B1(B[30]), .B2(n269), .ZN(n25) );
  AOI222_X1 U37 ( .A1(D[30]), .A2(n281), .B1(E[30]), .B2(n278), .C1(C[30]), 
        .C2(n275), .ZN(n26) );
  NAND2_X1 U38 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U39 ( .A1(A[31]), .A2(n273), .B1(B[31]), .B2(n270), .ZN(n23) );
  AOI222_X1 U40 ( .A1(D[31]), .A2(n282), .B1(E[31]), .B2(n279), .C1(C[31]), 
        .C2(n276), .ZN(n24) );
  NAND2_X1 U41 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U42 ( .A1(A[16]), .A2(n271), .B1(B[16]), .B2(n268), .ZN(n57) );
  AOI222_X1 U43 ( .A1(D[16]), .A2(n280), .B1(E[16]), .B2(n277), .C1(C[16]), 
        .C2(n274), .ZN(n58) );
  NAND2_X1 U44 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U45 ( .A1(A[20]), .A2(n272), .B1(B[20]), .B2(n269), .ZN(n47) );
  AOI222_X1 U46 ( .A1(D[20]), .A2(n281), .B1(E[20]), .B2(n278), .C1(C[20]), 
        .C2(n275), .ZN(n48) );
  NAND2_X1 U47 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U48 ( .A1(A[14]), .A2(n271), .B1(B[14]), .B2(n268), .ZN(n61) );
  AOI222_X1 U49 ( .A1(D[14]), .A2(n280), .B1(E[14]), .B2(n277), .C1(C[14]), 
        .C2(n274), .ZN(n62) );
  NAND2_X1 U50 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U51 ( .A1(A[18]), .A2(n271), .B1(B[18]), .B2(n268), .ZN(n53) );
  AOI222_X1 U52 ( .A1(D[18]), .A2(n280), .B1(E[18]), .B2(n277), .C1(C[18]), 
        .C2(n274), .ZN(n54) );
  NAND2_X1 U53 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U54 ( .A1(A[25]), .A2(n272), .B1(B[25]), .B2(n269), .ZN(n37) );
  AOI222_X1 U55 ( .A1(D[25]), .A2(n281), .B1(E[25]), .B2(n278), .C1(C[25]), 
        .C2(n275), .ZN(n38) );
  NAND2_X1 U56 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U57 ( .A1(A[21]), .A2(n272), .B1(B[21]), .B2(n269), .ZN(n45) );
  AOI222_X1 U58 ( .A1(D[21]), .A2(n281), .B1(E[21]), .B2(n278), .C1(C[21]), 
        .C2(n275), .ZN(n46) );
  AND2_X1 U59 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U60 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U61 ( .A1(A[15]), .A2(n271), .B1(B[15]), .B2(n268), .ZN(n59) );
  AOI222_X1 U62 ( .A1(D[15]), .A2(n280), .B1(E[15]), .B2(n277), .C1(C[15]), 
        .C2(n274), .ZN(n60) );
  NAND2_X1 U63 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U64 ( .A1(A[19]), .A2(n271), .B1(B[19]), .B2(n268), .ZN(n51) );
  AOI222_X1 U65 ( .A1(D[19]), .A2(n280), .B1(E[19]), .B2(n277), .C1(C[19]), 
        .C2(n274), .ZN(n52) );
  NAND2_X1 U66 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U67 ( .A1(A[17]), .A2(n271), .B1(B[17]), .B2(n268), .ZN(n55) );
  AOI222_X1 U68 ( .A1(D[17]), .A2(n280), .B1(E[17]), .B2(n277), .C1(C[17]), 
        .C2(n274), .ZN(n56) );
  NAND2_X1 U69 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U70 ( .A1(A[12]), .A2(n271), .B1(B[12]), .B2(n268), .ZN(n65) );
  AOI222_X1 U71 ( .A1(D[12]), .A2(n280), .B1(E[12]), .B2(n277), .C1(C[12]), 
        .C2(n274), .ZN(n66) );
  NAND2_X1 U72 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U73 ( .A1(A[13]), .A2(n271), .B1(B[13]), .B2(n268), .ZN(n63) );
  AOI222_X1 U74 ( .A1(D[13]), .A2(n280), .B1(E[13]), .B2(n277), .C1(C[13]), 
        .C2(n274), .ZN(n64) );
  NAND2_X1 U75 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U76 ( .A1(A[23]), .A2(n272), .B1(B[23]), .B2(n269), .ZN(n41) );
  AOI222_X1 U77 ( .A1(D[23]), .A2(n281), .B1(E[23]), .B2(n278), .C1(C[23]), 
        .C2(n275), .ZN(n42) );
  NAND2_X1 U78 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U79 ( .A1(A[27]), .A2(n272), .B1(B[27]), .B2(n269), .ZN(n33) );
  AOI222_X1 U80 ( .A1(D[27]), .A2(n281), .B1(E[27]), .B2(n278), .C1(C[27]), 
        .C2(n275), .ZN(n34) );
  NAND2_X1 U81 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U82 ( .A1(A[24]), .A2(n272), .B1(B[24]), .B2(n269), .ZN(n39) );
  AOI222_X1 U83 ( .A1(D[24]), .A2(n281), .B1(E[24]), .B2(n278), .C1(C[24]), 
        .C2(n275), .ZN(n40) );
  INV_X1 U84 ( .A(Sel[1]), .ZN(n75) );
  NAND2_X1 U85 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U86 ( .A1(A[6]), .A2(n273), .B1(B[6]), .B2(n270), .ZN(n15) );
  AOI222_X1 U87 ( .A1(D[6]), .A2(n282), .B1(E[6]), .B2(n279), .C1(C[6]), .C2(
        n276), .ZN(n16) );
  NAND2_X1 U88 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U89 ( .A1(A[3]), .A2(n273), .B1(B[3]), .B2(n270), .ZN(n21) );
  AOI222_X1 U90 ( .A1(D[3]), .A2(n282), .B1(E[3]), .B2(n279), .C1(C[3]), .C2(
        n276), .ZN(n22) );
  NAND2_X1 U91 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U92 ( .A1(A[7]), .A2(n273), .B1(B[7]), .B2(n270), .ZN(n13) );
  AOI222_X1 U93 ( .A1(D[7]), .A2(n282), .B1(E[7]), .B2(n279), .C1(C[7]), .C2(
        n276), .ZN(n14) );
  NAND2_X1 U94 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U95 ( .A1(A[4]), .A2(n273), .B1(B[4]), .B2(n270), .ZN(n19) );
  AOI222_X1 U96 ( .A1(D[4]), .A2(n282), .B1(E[4]), .B2(n279), .C1(C[4]), .C2(
        n276), .ZN(n20) );
  NAND2_X1 U97 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U98 ( .A1(A[8]), .A2(n273), .B1(B[8]), .B2(n270), .ZN(n11) );
  AOI222_X1 U99 ( .A1(D[8]), .A2(n282), .B1(E[8]), .B2(n279), .C1(C[8]), .C2(
        n276), .ZN(n12) );
  NAND2_X1 U100 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U101 ( .A1(A[9]), .A2(n273), .B1(B[9]), .B2(n270), .ZN(n4) );
  AOI222_X1 U102 ( .A1(D[9]), .A2(n282), .B1(E[9]), .B2(n279), .C1(C[9]), .C2(
        n276), .ZN(n5) );
  NAND2_X1 U103 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U104 ( .A1(A[5]), .A2(n273), .B1(B[5]), .B2(n270), .ZN(n17) );
  AOI222_X1 U105 ( .A1(D[5]), .A2(n282), .B1(E[5]), .B2(n279), .C1(C[5]), .C2(
        n276), .ZN(n18) );
  NAND2_X1 U106 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U107 ( .A1(A[2]), .A2(n272), .B1(B[2]), .B2(n269), .ZN(n27) );
  AOI222_X1 U108 ( .A1(D[2]), .A2(n281), .B1(E[2]), .B2(n278), .C1(C[2]), .C2(
        n275), .ZN(n28) );
  NAND2_X1 U109 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U110 ( .A1(A[10]), .A2(n271), .B1(B[10]), .B2(n268), .ZN(n69) );
  AOI222_X1 U111 ( .A1(D[10]), .A2(n280), .B1(E[10]), .B2(n277), .C1(C[10]), 
        .C2(n274), .ZN(n70) );
  NAND2_X1 U112 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U113 ( .A1(A[11]), .A2(n271), .B1(B[11]), .B2(n268), .ZN(n67) );
  AOI222_X1 U114 ( .A1(D[11]), .A2(n280), .B1(E[11]), .B2(n277), .C1(C[11]), 
        .C2(n274), .ZN(n68) );
  NAND2_X1 U115 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U116 ( .A1(A[0]), .A2(n271), .B1(B[0]), .B2(n268), .ZN(n71) );
  AOI222_X1 U117 ( .A1(D[0]), .A2(n280), .B1(E[0]), .B2(n277), .C1(C[0]), .C2(
        n274), .ZN(n72) );
  NAND2_X1 U118 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U119 ( .A1(A[1]), .A2(n271), .B1(B[1]), .B2(n268), .ZN(n49) );
  AOI222_X1 U120 ( .A1(D[1]), .A2(n280), .B1(E[1]), .B2(n277), .C1(C[1]), .C2(
        n274), .ZN(n50) );
endmodule


module mux_N32_3 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279;

  BUF_X1 U1 ( .A(n10), .Z(n265) );
  BUF_X1 U2 ( .A(n10), .Z(n266) );
  BUF_X1 U3 ( .A(n10), .Z(n267) );
  BUF_X1 U4 ( .A(n6), .Z(n277) );
  BUF_X1 U5 ( .A(n6), .Z(n278) );
  BUF_X1 U6 ( .A(n9), .Z(n268) );
  BUF_X1 U7 ( .A(n9), .Z(n269) );
  BUF_X1 U8 ( .A(n7), .Z(n274) );
  BUF_X1 U9 ( .A(n7), .Z(n275) );
  BUF_X1 U10 ( .A(n8), .Z(n271) );
  BUF_X1 U11 ( .A(n8), .Z(n272) );
  BUF_X1 U12 ( .A(n9), .Z(n270) );
  BUF_X1 U13 ( .A(n7), .Z(n276) );
  BUF_X1 U14 ( .A(n8), .Z(n273) );
  BUF_X1 U15 ( .A(n6), .Z(n279) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  INV_X1 U22 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U23 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U24 ( .A1(A[24]), .A2(n269), .B1(B[24]), .B2(n266), .ZN(n39) );
  AOI222_X1 U25 ( .A1(D[24]), .A2(n278), .B1(E[24]), .B2(n275), .C1(C[24]), 
        .C2(n272), .ZN(n40) );
  NAND2_X1 U26 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U27 ( .A1(A[20]), .A2(n269), .B1(B[20]), .B2(n266), .ZN(n47) );
  AOI222_X1 U28 ( .A1(D[20]), .A2(n278), .B1(E[20]), .B2(n275), .C1(C[20]), 
        .C2(n272), .ZN(n48) );
  NAND2_X1 U29 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U30 ( .A1(A[14]), .A2(n268), .B1(B[14]), .B2(n265), .ZN(n61) );
  AOI222_X1 U31 ( .A1(D[14]), .A2(n277), .B1(E[14]), .B2(n274), .C1(C[14]), 
        .C2(n271), .ZN(n62) );
  NAND2_X1 U32 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U33 ( .A1(A[18]), .A2(n268), .B1(B[18]), .B2(n265), .ZN(n53) );
  AOI222_X1 U34 ( .A1(D[18]), .A2(n277), .B1(E[18]), .B2(n274), .C1(C[18]), 
        .C2(n271), .ZN(n54) );
  NAND2_X1 U35 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U36 ( .A1(A[12]), .A2(n268), .B1(B[12]), .B2(n265), .ZN(n65) );
  AOI222_X1 U37 ( .A1(D[12]), .A2(n277), .B1(E[12]), .B2(n274), .C1(C[12]), 
        .C2(n271), .ZN(n66) );
  NAND2_X1 U38 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U39 ( .A1(A[16]), .A2(n268), .B1(B[16]), .B2(n265), .ZN(n57) );
  AOI222_X1 U40 ( .A1(D[16]), .A2(n277), .B1(E[16]), .B2(n274), .C1(C[16]), 
        .C2(n271), .ZN(n58) );
  NAND2_X1 U41 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U42 ( .A1(A[23]), .A2(n269), .B1(B[23]), .B2(n266), .ZN(n41) );
  AOI222_X1 U43 ( .A1(D[23]), .A2(n278), .B1(E[23]), .B2(n275), .C1(C[23]), 
        .C2(n272), .ZN(n42) );
  NAND2_X1 U44 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U45 ( .A1(A[19]), .A2(n268), .B1(B[19]), .B2(n265), .ZN(n51) );
  AOI222_X1 U46 ( .A1(D[19]), .A2(n277), .B1(E[19]), .B2(n274), .C1(C[19]), 
        .C2(n271), .ZN(n52) );
  AND2_X1 U47 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U48 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U49 ( .A1(A[13]), .A2(n268), .B1(B[13]), .B2(n265), .ZN(n63) );
  AOI222_X1 U50 ( .A1(D[13]), .A2(n277), .B1(E[13]), .B2(n274), .C1(C[13]), 
        .C2(n271), .ZN(n64) );
  NAND2_X1 U51 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U52 ( .A1(A[17]), .A2(n268), .B1(B[17]), .B2(n265), .ZN(n55) );
  AOI222_X1 U53 ( .A1(D[17]), .A2(n277), .B1(E[17]), .B2(n274), .C1(C[17]), 
        .C2(n271), .ZN(n56) );
  NAND2_X1 U54 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U55 ( .A1(A[15]), .A2(n268), .B1(B[15]), .B2(n265), .ZN(n59) );
  AOI222_X1 U56 ( .A1(D[15]), .A2(n277), .B1(E[15]), .B2(n274), .C1(C[15]), 
        .C2(n271), .ZN(n60) );
  NAND2_X1 U57 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U58 ( .A1(A[10]), .A2(n268), .B1(B[10]), .B2(n265), .ZN(n69) );
  AOI222_X1 U59 ( .A1(D[10]), .A2(n277), .B1(E[10]), .B2(n274), .C1(C[10]), 
        .C2(n271), .ZN(n70) );
  NAND2_X1 U60 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U61 ( .A1(A[11]), .A2(n268), .B1(B[11]), .B2(n265), .ZN(n67) );
  AOI222_X1 U62 ( .A1(D[11]), .A2(n277), .B1(E[11]), .B2(n274), .C1(C[11]), 
        .C2(n271), .ZN(n68) );
  NAND2_X1 U63 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U64 ( .A1(A[21]), .A2(n269), .B1(B[21]), .B2(n266), .ZN(n45) );
  AOI222_X1 U65 ( .A1(D[21]), .A2(n278), .B1(E[21]), .B2(n275), .C1(C[21]), 
        .C2(n272), .ZN(n46) );
  NAND2_X1 U66 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U67 ( .A1(A[25]), .A2(n269), .B1(B[25]), .B2(n266), .ZN(n37) );
  AOI222_X1 U68 ( .A1(D[25]), .A2(n278), .B1(E[25]), .B2(n275), .C1(C[25]), 
        .C2(n272), .ZN(n38) );
  NAND2_X1 U69 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U70 ( .A1(A[26]), .A2(n269), .B1(B[26]), .B2(n266), .ZN(n35) );
  AOI222_X1 U71 ( .A1(D[26]), .A2(n278), .B1(E[26]), .B2(n275), .C1(C[26]), 
        .C2(n272), .ZN(n36) );
  NAND2_X1 U72 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U73 ( .A1(A[27]), .A2(n269), .B1(B[27]), .B2(n266), .ZN(n33) );
  AOI222_X1 U74 ( .A1(D[27]), .A2(n278), .B1(E[27]), .B2(n275), .C1(C[27]), 
        .C2(n272), .ZN(n34) );
  NAND2_X1 U75 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U76 ( .A1(A[28]), .A2(n269), .B1(B[28]), .B2(n266), .ZN(n31) );
  AOI222_X1 U77 ( .A1(D[28]), .A2(n278), .B1(E[28]), .B2(n275), .C1(C[28]), 
        .C2(n272), .ZN(n32) );
  NAND2_X1 U78 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U79 ( .A1(A[29]), .A2(n269), .B1(B[29]), .B2(n266), .ZN(n29) );
  AOI222_X1 U80 ( .A1(D[29]), .A2(n278), .B1(E[29]), .B2(n275), .C1(C[29]), 
        .C2(n272), .ZN(n30) );
  NAND2_X1 U81 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U82 ( .A1(A[30]), .A2(n269), .B1(B[30]), .B2(n266), .ZN(n25) );
  AOI222_X1 U83 ( .A1(D[30]), .A2(n278), .B1(E[30]), .B2(n275), .C1(C[30]), 
        .C2(n272), .ZN(n26) );
  NAND2_X1 U84 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U85 ( .A1(A[31]), .A2(n270), .B1(B[31]), .B2(n267), .ZN(n23) );
  AOI222_X1 U86 ( .A1(D[31]), .A2(n279), .B1(E[31]), .B2(n276), .C1(C[31]), 
        .C2(n273), .ZN(n24) );
  NAND2_X1 U87 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U88 ( .A1(A[22]), .A2(n269), .B1(B[22]), .B2(n266), .ZN(n43) );
  AOI222_X1 U89 ( .A1(D[22]), .A2(n278), .B1(E[22]), .B2(n275), .C1(C[22]), 
        .C2(n272), .ZN(n44) );
  NAND2_X1 U90 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U91 ( .A1(A[9]), .A2(n270), .B1(B[9]), .B2(n267), .ZN(n4) );
  AOI222_X1 U92 ( .A1(D[9]), .A2(n279), .B1(E[9]), .B2(n276), .C1(C[9]), .C2(
        n273), .ZN(n5) );
  NAND2_X1 U93 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U94 ( .A1(A[5]), .A2(n270), .B1(B[5]), .B2(n267), .ZN(n17) );
  AOI222_X1 U95 ( .A1(D[5]), .A2(n279), .B1(E[5]), .B2(n276), .C1(C[5]), .C2(
        n273), .ZN(n18) );
  NAND2_X1 U96 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U97 ( .A1(A[6]), .A2(n270), .B1(B[6]), .B2(n267), .ZN(n15) );
  AOI222_X1 U98 ( .A1(D[6]), .A2(n279), .B1(E[6]), .B2(n276), .C1(C[6]), .C2(
        n273), .ZN(n16) );
  NAND2_X1 U99 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U100 ( .A1(A[3]), .A2(n270), .B1(B[3]), .B2(n267), .ZN(n21) );
  AOI222_X1 U101 ( .A1(D[3]), .A2(n279), .B1(E[3]), .B2(n276), .C1(C[3]), .C2(
        n273), .ZN(n22) );
  NAND2_X1 U102 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U103 ( .A1(A[7]), .A2(n270), .B1(B[7]), .B2(n267), .ZN(n13) );
  AOI222_X1 U104 ( .A1(D[7]), .A2(n279), .B1(E[7]), .B2(n276), .C1(C[7]), .C2(
        n273), .ZN(n14) );
  NAND2_X1 U105 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U106 ( .A1(A[4]), .A2(n270), .B1(B[4]), .B2(n267), .ZN(n19) );
  AOI222_X1 U107 ( .A1(D[4]), .A2(n279), .B1(E[4]), .B2(n276), .C1(C[4]), .C2(
        n273), .ZN(n20) );
  NAND2_X1 U108 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U109 ( .A1(A[8]), .A2(n270), .B1(B[8]), .B2(n267), .ZN(n11) );
  AOI222_X1 U110 ( .A1(D[8]), .A2(n279), .B1(E[8]), .B2(n276), .C1(C[8]), .C2(
        n273), .ZN(n12) );
  NAND2_X1 U111 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U112 ( .A1(A[1]), .A2(n268), .B1(B[1]), .B2(n265), .ZN(n49) );
  AOI222_X1 U113 ( .A1(D[1]), .A2(n277), .B1(E[1]), .B2(n274), .C1(C[1]), .C2(
        n271), .ZN(n50) );
  NAND2_X1 U114 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U115 ( .A1(A[2]), .A2(n269), .B1(B[2]), .B2(n266), .ZN(n27) );
  AOI222_X1 U116 ( .A1(D[2]), .A2(n278), .B1(E[2]), .B2(n275), .C1(C[2]), .C2(
        n272), .ZN(n28) );
  NAND2_X1 U117 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U118 ( .A1(A[0]), .A2(n268), .B1(B[0]), .B2(n265), .ZN(n71) );
  AOI222_X1 U119 ( .A1(D[0]), .A2(n277), .B1(E[0]), .B2(n274), .C1(C[0]), .C2(
        n271), .ZN(n72) );
  INV_X1 U120 ( .A(Sel[1]), .ZN(n75) );
endmodule


module mux_N32_4 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294;

  BUF_X1 U1 ( .A(n10), .Z(n280) );
  BUF_X1 U2 ( .A(n10), .Z(n281) );
  BUF_X1 U3 ( .A(n10), .Z(n282) );
  BUF_X1 U4 ( .A(n6), .Z(n292) );
  BUF_X1 U5 ( .A(n6), .Z(n293) );
  BUF_X1 U6 ( .A(n9), .Z(n283) );
  BUF_X1 U7 ( .A(n9), .Z(n284) );
  BUF_X1 U8 ( .A(n7), .Z(n289) );
  BUF_X1 U9 ( .A(n7), .Z(n290) );
  BUF_X1 U10 ( .A(n8), .Z(n286) );
  BUF_X1 U11 ( .A(n8), .Z(n287) );
  BUF_X1 U12 ( .A(n9), .Z(n285) );
  BUF_X1 U13 ( .A(n7), .Z(n291) );
  BUF_X1 U14 ( .A(n8), .Z(n288) );
  BUF_X1 U15 ( .A(n6), .Z(n294) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  INV_X1 U22 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U23 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U24 ( .A1(A[22]), .A2(n284), .B1(B[22]), .B2(n281), .ZN(n43) );
  AOI222_X1 U25 ( .A1(D[22]), .A2(n293), .B1(E[22]), .B2(n290), .C1(C[22]), 
        .C2(n287), .ZN(n44) );
  NAND2_X1 U26 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U27 ( .A1(A[8]), .A2(n285), .B1(B[8]), .B2(n282), .ZN(n11) );
  AOI222_X1 U28 ( .A1(D[8]), .A2(n294), .B1(E[8]), .B2(n291), .C1(C[8]), .C2(
        n288), .ZN(n12) );
  NAND2_X1 U29 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U30 ( .A1(A[18]), .A2(n283), .B1(B[18]), .B2(n280), .ZN(n53) );
  AOI222_X1 U31 ( .A1(D[18]), .A2(n292), .B1(E[18]), .B2(n289), .C1(C[18]), 
        .C2(n286), .ZN(n54) );
  NAND2_X1 U32 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U33 ( .A1(A[25]), .A2(n284), .B1(B[25]), .B2(n281), .ZN(n37) );
  AOI222_X1 U34 ( .A1(D[25]), .A2(n293), .B1(E[25]), .B2(n290), .C1(C[25]), 
        .C2(n287), .ZN(n38) );
  NAND2_X1 U35 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U36 ( .A1(A[26]), .A2(n284), .B1(B[26]), .B2(n281), .ZN(n35) );
  AOI222_X1 U37 ( .A1(D[26]), .A2(n293), .B1(E[26]), .B2(n290), .C1(C[26]), 
        .C2(n287), .ZN(n36) );
  NAND2_X1 U38 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U39 ( .A1(A[27]), .A2(n284), .B1(B[27]), .B2(n281), .ZN(n33) );
  AOI222_X1 U40 ( .A1(D[27]), .A2(n293), .B1(E[27]), .B2(n290), .C1(C[27]), 
        .C2(n287), .ZN(n34) );
  NAND2_X1 U41 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U42 ( .A1(A[28]), .A2(n284), .B1(B[28]), .B2(n281), .ZN(n31) );
  AOI222_X1 U43 ( .A1(D[28]), .A2(n293), .B1(E[28]), .B2(n290), .C1(C[28]), 
        .C2(n287), .ZN(n32) );
  NAND2_X1 U44 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U45 ( .A1(A[24]), .A2(n284), .B1(B[24]), .B2(n281), .ZN(n39) );
  AOI222_X1 U46 ( .A1(D[24]), .A2(n293), .B1(E[24]), .B2(n290), .C1(C[24]), 
        .C2(n287), .ZN(n40) );
  NAND2_X1 U47 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U48 ( .A1(A[29]), .A2(n284), .B1(B[29]), .B2(n281), .ZN(n29) );
  AOI222_X1 U49 ( .A1(D[29]), .A2(n293), .B1(E[29]), .B2(n290), .C1(C[29]), 
        .C2(n287), .ZN(n30) );
  NAND2_X1 U50 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U51 ( .A1(A[30]), .A2(n284), .B1(B[30]), .B2(n281), .ZN(n25) );
  AOI222_X1 U52 ( .A1(D[30]), .A2(n293), .B1(E[30]), .B2(n290), .C1(C[30]), 
        .C2(n287), .ZN(n26) );
  NAND2_X1 U53 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U54 ( .A1(A[31]), .A2(n285), .B1(B[31]), .B2(n282), .ZN(n23) );
  AOI222_X1 U55 ( .A1(D[31]), .A2(n294), .B1(E[31]), .B2(n291), .C1(C[31]), 
        .C2(n288), .ZN(n24) );
  NAND2_X1 U56 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U57 ( .A1(A[12]), .A2(n283), .B1(B[12]), .B2(n280), .ZN(n65) );
  AOI222_X1 U58 ( .A1(D[12]), .A2(n292), .B1(E[12]), .B2(n289), .C1(C[12]), 
        .C2(n286), .ZN(n66) );
  NAND2_X1 U59 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U60 ( .A1(A[9]), .A2(n285), .B1(B[9]), .B2(n282), .ZN(n4) );
  AOI222_X1 U61 ( .A1(D[9]), .A2(n294), .B1(E[9]), .B2(n291), .C1(C[9]), .C2(
        n288), .ZN(n5) );
  NAND2_X1 U62 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U63 ( .A1(A[16]), .A2(n283), .B1(B[16]), .B2(n280), .ZN(n57) );
  AOI222_X1 U64 ( .A1(D[16]), .A2(n292), .B1(E[16]), .B2(n289), .C1(C[16]), 
        .C2(n286), .ZN(n58) );
  NAND2_X1 U65 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U66 ( .A1(A[10]), .A2(n283), .B1(B[10]), .B2(n280), .ZN(n69) );
  AOI222_X1 U67 ( .A1(D[10]), .A2(n292), .B1(E[10]), .B2(n289), .C1(C[10]), 
        .C2(n286), .ZN(n70) );
  NAND2_X1 U68 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U69 ( .A1(A[14]), .A2(n283), .B1(B[14]), .B2(n280), .ZN(n61) );
  AOI222_X1 U70 ( .A1(D[14]), .A2(n292), .B1(E[14]), .B2(n289), .C1(C[14]), 
        .C2(n286), .ZN(n62) );
  NAND2_X1 U71 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U72 ( .A1(A[21]), .A2(n284), .B1(B[21]), .B2(n281), .ZN(n45) );
  AOI222_X1 U73 ( .A1(D[21]), .A2(n293), .B1(E[21]), .B2(n290), .C1(C[21]), 
        .C2(n287), .ZN(n46) );
  NAND2_X1 U74 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U75 ( .A1(A[17]), .A2(n283), .B1(B[17]), .B2(n280), .ZN(n55) );
  AOI222_X1 U76 ( .A1(D[17]), .A2(n292), .B1(E[17]), .B2(n289), .C1(C[17]), 
        .C2(n286), .ZN(n56) );
  AND2_X1 U77 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U78 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U79 ( .A1(A[11]), .A2(n283), .B1(B[11]), .B2(n280), .ZN(n67) );
  AOI222_X1 U80 ( .A1(D[11]), .A2(n292), .B1(E[11]), .B2(n289), .C1(C[11]), 
        .C2(n286), .ZN(n68) );
  NAND2_X1 U81 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U82 ( .A1(A[15]), .A2(n283), .B1(B[15]), .B2(n280), .ZN(n59) );
  AOI222_X1 U83 ( .A1(D[15]), .A2(n292), .B1(E[15]), .B2(n289), .C1(C[15]), 
        .C2(n286), .ZN(n60) );
  NAND2_X1 U84 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U85 ( .A1(A[13]), .A2(n283), .B1(B[13]), .B2(n280), .ZN(n63) );
  AOI222_X1 U86 ( .A1(D[13]), .A2(n292), .B1(E[13]), .B2(n289), .C1(C[13]), 
        .C2(n286), .ZN(n64) );
  NAND2_X1 U87 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U88 ( .A1(A[20]), .A2(n284), .B1(B[20]), .B2(n281), .ZN(n47) );
  AOI222_X1 U89 ( .A1(D[20]), .A2(n293), .B1(E[20]), .B2(n290), .C1(C[20]), 
        .C2(n287), .ZN(n48) );
  NAND2_X1 U90 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U91 ( .A1(A[19]), .A2(n283), .B1(B[19]), .B2(n280), .ZN(n51) );
  AOI222_X1 U92 ( .A1(D[19]), .A2(n292), .B1(E[19]), .B2(n289), .C1(C[19]), 
        .C2(n286), .ZN(n52) );
  INV_X1 U93 ( .A(Sel[1]), .ZN(n75) );
  NAND2_X1 U94 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U95 ( .A1(A[5]), .A2(n285), .B1(B[5]), .B2(n282), .ZN(n17) );
  AOI222_X1 U96 ( .A1(D[5]), .A2(n294), .B1(E[5]), .B2(n291), .C1(C[5]), .C2(
        n288), .ZN(n18) );
  NAND2_X1 U97 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U98 ( .A1(A[6]), .A2(n285), .B1(B[6]), .B2(n282), .ZN(n15) );
  AOI222_X1 U99 ( .A1(D[6]), .A2(n294), .B1(E[6]), .B2(n291), .C1(C[6]), .C2(
        n288), .ZN(n16) );
  NAND2_X1 U100 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U101 ( .A1(A[3]), .A2(n285), .B1(B[3]), .B2(n282), .ZN(n21) );
  AOI222_X1 U102 ( .A1(D[3]), .A2(n294), .B1(E[3]), .B2(n291), .C1(C[3]), .C2(
        n288), .ZN(n22) );
  NAND2_X1 U103 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U104 ( .A1(A[7]), .A2(n285), .B1(B[7]), .B2(n282), .ZN(n13) );
  AOI222_X1 U105 ( .A1(D[7]), .A2(n294), .B1(E[7]), .B2(n291), .C1(C[7]), .C2(
        n288), .ZN(n14) );
  NAND2_X1 U106 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U107 ( .A1(A[4]), .A2(n285), .B1(B[4]), .B2(n282), .ZN(n19) );
  AOI222_X1 U108 ( .A1(D[4]), .A2(n294), .B1(E[4]), .B2(n291), .C1(C[4]), .C2(
        n288), .ZN(n20) );
  NAND2_X1 U109 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U110 ( .A1(A[1]), .A2(n283), .B1(B[1]), .B2(n280), .ZN(n49) );
  AOI222_X1 U111 ( .A1(D[1]), .A2(n292), .B1(E[1]), .B2(n289), .C1(C[1]), .C2(
        n286), .ZN(n50) );
  NAND2_X1 U112 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U113 ( .A1(A[2]), .A2(n284), .B1(B[2]), .B2(n281), .ZN(n27) );
  AOI222_X1 U114 ( .A1(D[2]), .A2(n293), .B1(E[2]), .B2(n290), .C1(C[2]), .C2(
        n287), .ZN(n28) );
  NAND2_X1 U115 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U116 ( .A1(A[23]), .A2(n284), .B1(B[23]), .B2(n281), .ZN(n41) );
  AOI222_X1 U117 ( .A1(D[23]), .A2(n293), .B1(E[23]), .B2(n290), .C1(C[23]), 
        .C2(n287), .ZN(n42) );
  NAND2_X1 U118 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U119 ( .A1(A[0]), .A2(n283), .B1(B[0]), .B2(n280), .ZN(n71) );
  AOI222_X1 U120 ( .A1(D[0]), .A2(n292), .B1(E[0]), .B2(n289), .C1(C[0]), .C2(
        n286), .ZN(n72) );
endmodule


module mux_N32_5 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288;

  BUF_X1 U1 ( .A(n10), .Z(n274) );
  BUF_X1 U2 ( .A(n10), .Z(n275) );
  BUF_X1 U3 ( .A(n10), .Z(n276) );
  BUF_X1 U4 ( .A(n6), .Z(n286) );
  BUF_X1 U5 ( .A(n6), .Z(n287) );
  BUF_X1 U6 ( .A(n9), .Z(n277) );
  BUF_X1 U7 ( .A(n9), .Z(n278) );
  BUF_X1 U8 ( .A(n7), .Z(n283) );
  BUF_X1 U9 ( .A(n7), .Z(n284) );
  BUF_X1 U10 ( .A(n8), .Z(n280) );
  BUF_X1 U11 ( .A(n8), .Z(n281) );
  BUF_X1 U12 ( .A(n9), .Z(n279) );
  BUF_X1 U13 ( .A(n7), .Z(n285) );
  BUF_X1 U14 ( .A(n8), .Z(n282) );
  BUF_X1 U15 ( .A(n6), .Z(n288) );
  AND2_X1 U16 ( .A1(n74), .A2(n73), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n73), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n73), .ZN(n8) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n74) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  INV_X1 U22 ( .A(Sel[2]), .ZN(n73) );
  NAND2_X1 U23 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U24 ( .A1(A[20]), .A2(n278), .B1(B[20]), .B2(n275), .ZN(n47) );
  AOI222_X1 U25 ( .A1(D[20]), .A2(n287), .B1(C[20]), .B2(n284), .C1(E[20]), 
        .C2(n281), .ZN(n48) );
  NAND2_X1 U26 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U27 ( .A1(A[16]), .A2(n277), .B1(B[16]), .B2(n274), .ZN(n57) );
  AOI222_X1 U28 ( .A1(D[16]), .A2(n286), .B1(C[16]), .B2(n283), .C1(E[16]), 
        .C2(n280), .ZN(n58) );
  NAND2_X1 U29 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U30 ( .A1(A[10]), .A2(n277), .B1(B[10]), .B2(n274), .ZN(n69) );
  AOI222_X1 U31 ( .A1(D[10]), .A2(n286), .B1(C[10]), .B2(n283), .C1(E[10]), 
        .C2(n280), .ZN(n70) );
  NAND2_X1 U32 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U33 ( .A1(A[14]), .A2(n277), .B1(B[14]), .B2(n274), .ZN(n61) );
  AOI222_X1 U34 ( .A1(D[14]), .A2(n286), .B1(C[14]), .B2(n283), .C1(E[14]), 
        .C2(n280), .ZN(n62) );
  NAND2_X1 U35 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U36 ( .A1(A[8]), .A2(n279), .B1(B[8]), .B2(n276), .ZN(n11) );
  AOI222_X1 U37 ( .A1(D[8]), .A2(n288), .B1(C[8]), .B2(n285), .C1(E[8]), .C2(
        n282), .ZN(n12) );
  NAND2_X1 U38 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U39 ( .A1(A[12]), .A2(n277), .B1(B[12]), .B2(n274), .ZN(n65) );
  AOI222_X1 U40 ( .A1(D[12]), .A2(n286), .B1(C[12]), .B2(n283), .C1(E[12]), 
        .C2(n280), .ZN(n66) );
  NAND2_X1 U41 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U42 ( .A1(A[19]), .A2(n277), .B1(B[19]), .B2(n274), .ZN(n51) );
  AOI222_X1 U43 ( .A1(D[19]), .A2(n286), .B1(C[19]), .B2(n283), .C1(E[19]), 
        .C2(n280), .ZN(n52) );
  NAND2_X1 U44 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U45 ( .A1(A[15]), .A2(n277), .B1(B[15]), .B2(n274), .ZN(n59) );
  AOI222_X1 U46 ( .A1(D[15]), .A2(n286), .B1(C[15]), .B2(n283), .C1(E[15]), 
        .C2(n280), .ZN(n60) );
  AND2_X1 U47 ( .A1(Sel[2]), .A2(n74), .ZN(n7) );
  NAND2_X1 U48 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U49 ( .A1(A[9]), .A2(n279), .B1(B[9]), .B2(n276), .ZN(n4) );
  AOI222_X1 U50 ( .A1(D[9]), .A2(n288), .B1(C[9]), .B2(n285), .C1(E[9]), .C2(
        n282), .ZN(n5) );
  NAND2_X1 U51 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U52 ( .A1(A[13]), .A2(n277), .B1(B[13]), .B2(n274), .ZN(n63) );
  AOI222_X1 U53 ( .A1(D[13]), .A2(n286), .B1(C[13]), .B2(n283), .C1(E[13]), 
        .C2(n280), .ZN(n64) );
  NAND2_X1 U54 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U55 ( .A1(A[7]), .A2(n279), .B1(B[7]), .B2(n276), .ZN(n13) );
  AOI222_X1 U56 ( .A1(D[7]), .A2(n288), .B1(C[7]), .B2(n285), .C1(E[7]), .C2(
        n282), .ZN(n14) );
  NAND2_X1 U57 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U58 ( .A1(A[17]), .A2(n277), .B1(B[17]), .B2(n274), .ZN(n55) );
  AOI222_X1 U59 ( .A1(D[17]), .A2(n286), .B1(C[17]), .B2(n283), .C1(E[17]), 
        .C2(n280), .ZN(n56) );
  NAND2_X1 U60 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U61 ( .A1(A[11]), .A2(n277), .B1(B[11]), .B2(n274), .ZN(n67) );
  AOI222_X1 U62 ( .A1(D[11]), .A2(n286), .B1(C[11]), .B2(n283), .C1(E[11]), 
        .C2(n280), .ZN(n68) );
  NAND2_X1 U63 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U64 ( .A1(A[6]), .A2(n279), .B1(B[6]), .B2(n276), .ZN(n15) );
  AOI222_X1 U65 ( .A1(D[6]), .A2(n288), .B1(C[6]), .B2(n285), .C1(E[6]), .C2(
        n282), .ZN(n16) );
  NAND2_X1 U66 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U67 ( .A1(A[18]), .A2(n277), .B1(B[18]), .B2(n274), .ZN(n53) );
  AOI222_X1 U68 ( .A1(D[18]), .A2(n286), .B1(C[18]), .B2(n283), .C1(E[18]), 
        .C2(n280), .ZN(n54) );
  NAND2_X1 U69 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U70 ( .A1(A[21]), .A2(n278), .B1(B[21]), .B2(n275), .ZN(n45) );
  AOI222_X1 U71 ( .A1(D[21]), .A2(n287), .B1(C[21]), .B2(n284), .C1(E[21]), 
        .C2(n281), .ZN(n46) );
  NAND2_X1 U72 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U73 ( .A1(A[5]), .A2(n279), .B1(B[5]), .B2(n276), .ZN(n17) );
  AOI222_X1 U74 ( .A1(D[5]), .A2(n288), .B1(C[5]), .B2(n285), .C1(E[5]), .C2(
        n282), .ZN(n18) );
  NAND2_X1 U75 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U76 ( .A1(A[3]), .A2(n279), .B1(B[3]), .B2(n276), .ZN(n21) );
  AOI222_X1 U77 ( .A1(D[3]), .A2(n288), .B1(C[3]), .B2(n285), .C1(E[3]), .C2(
        n282), .ZN(n22) );
  NAND2_X1 U78 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U79 ( .A1(A[4]), .A2(n279), .B1(B[4]), .B2(n276), .ZN(n19) );
  AOI222_X1 U80 ( .A1(D[4]), .A2(n288), .B1(C[4]), .B2(n285), .C1(E[4]), .C2(
        n282), .ZN(n20) );
  NAND2_X1 U81 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U82 ( .A1(A[31]), .A2(n279), .B1(B[31]), .B2(n276), .ZN(n23) );
  AOI222_X1 U83 ( .A1(D[31]), .A2(n288), .B1(C[31]), .B2(n285), .C1(E[31]), 
        .C2(n282), .ZN(n24) );
  NAND2_X1 U84 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U85 ( .A1(A[1]), .A2(n277), .B1(B[1]), .B2(n274), .ZN(n49) );
  AOI222_X1 U86 ( .A1(D[1]), .A2(n286), .B1(C[1]), .B2(n283), .C1(E[1]), .C2(
        n280), .ZN(n50) );
  NAND2_X1 U87 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U88 ( .A1(A[25]), .A2(n278), .B1(B[25]), .B2(n275), .ZN(n37) );
  AOI222_X1 U89 ( .A1(D[25]), .A2(n287), .B1(C[25]), .B2(n284), .C1(E[25]), 
        .C2(n281), .ZN(n38) );
  NAND2_X1 U90 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U91 ( .A1(A[2]), .A2(n278), .B1(B[2]), .B2(n275), .ZN(n27) );
  AOI222_X1 U92 ( .A1(D[2]), .A2(n287), .B1(C[2]), .B2(n284), .C1(E[2]), .C2(
        n281), .ZN(n28) );
  NAND2_X1 U93 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U94 ( .A1(A[26]), .A2(n278), .B1(B[26]), .B2(n275), .ZN(n35) );
  AOI222_X1 U95 ( .A1(D[26]), .A2(n287), .B1(C[26]), .B2(n284), .C1(E[26]), 
        .C2(n281), .ZN(n36) );
  NAND2_X1 U96 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U97 ( .A1(A[22]), .A2(n278), .B1(B[22]), .B2(n275), .ZN(n43) );
  AOI222_X1 U98 ( .A1(D[22]), .A2(n287), .B1(C[22]), .B2(n284), .C1(E[22]), 
        .C2(n281), .ZN(n44) );
  NAND2_X1 U99 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U100 ( .A1(A[27]), .A2(n278), .B1(B[27]), .B2(n275), .ZN(n33) );
  AOI222_X1 U101 ( .A1(D[27]), .A2(n287), .B1(C[27]), .B2(n284), .C1(E[27]), 
        .C2(n281), .ZN(n34) );
  NAND2_X1 U102 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U103 ( .A1(A[23]), .A2(n278), .B1(B[23]), .B2(n275), .ZN(n41) );
  AOI222_X1 U104 ( .A1(D[23]), .A2(n287), .B1(C[23]), .B2(n284), .C1(E[23]), 
        .C2(n281), .ZN(n42) );
  NAND2_X1 U105 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U106 ( .A1(A[0]), .A2(n277), .B1(B[0]), .B2(n274), .ZN(n71) );
  AOI222_X1 U107 ( .A1(D[0]), .A2(n286), .B1(C[0]), .B2(n283), .C1(E[0]), .C2(
        n280), .ZN(n72) );
  NAND2_X1 U108 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U109 ( .A1(A[28]), .A2(n278), .B1(B[28]), .B2(n275), .ZN(n31) );
  AOI222_X1 U110 ( .A1(D[28]), .A2(n287), .B1(C[28]), .B2(n284), .C1(E[28]), 
        .C2(n281), .ZN(n32) );
  NAND2_X1 U111 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U112 ( .A1(A[24]), .A2(n278), .B1(B[24]), .B2(n275), .ZN(n39) );
  AOI222_X1 U113 ( .A1(D[24]), .A2(n287), .B1(C[24]), .B2(n284), .C1(E[24]), 
        .C2(n281), .ZN(n40) );
  NAND2_X1 U114 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U115 ( .A1(A[29]), .A2(n278), .B1(B[29]), .B2(n275), .ZN(n29) );
  AOI222_X1 U116 ( .A1(D[29]), .A2(n287), .B1(C[29]), .B2(n284), .C1(E[29]), 
        .C2(n281), .ZN(n30) );
  NAND2_X1 U117 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U118 ( .A1(A[30]), .A2(n278), .B1(B[30]), .B2(n275), .ZN(n25) );
  AOI222_X1 U119 ( .A1(D[30]), .A2(n287), .B1(C[30]), .B2(n284), .C1(E[30]), 
        .C2(n281), .ZN(n26) );
  INV_X1 U120 ( .A(Sel[1]), .ZN(n75) );
endmodule


module mux_N32_6 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291;

  BUF_X1 U1 ( .A(n10), .Z(n277) );
  BUF_X1 U2 ( .A(n10), .Z(n278) );
  BUF_X1 U3 ( .A(n10), .Z(n279) );
  BUF_X1 U4 ( .A(n6), .Z(n289) );
  BUF_X1 U5 ( .A(n6), .Z(n290) );
  BUF_X1 U6 ( .A(n9), .Z(n280) );
  BUF_X1 U7 ( .A(n9), .Z(n281) );
  BUF_X1 U8 ( .A(n7), .Z(n286) );
  BUF_X1 U9 ( .A(n7), .Z(n287) );
  BUF_X1 U10 ( .A(n8), .Z(n283) );
  BUF_X1 U11 ( .A(n8), .Z(n284) );
  BUF_X1 U12 ( .A(n9), .Z(n282) );
  BUF_X1 U13 ( .A(n7), .Z(n288) );
  BUF_X1 U14 ( .A(n8), .Z(n285) );
  BUF_X1 U15 ( .A(n6), .Z(n291) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  NAND2_X1 U22 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U23 ( .A1(A[24]), .A2(n281), .B1(B[24]), .B2(n278), .ZN(n39) );
  AOI222_X1 U24 ( .A1(D[24]), .A2(n290), .B1(E[24]), .B2(n287), .C1(C[24]), 
        .C2(n284), .ZN(n40) );
  NAND2_X1 U25 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U26 ( .A1(A[25]), .A2(n281), .B1(B[25]), .B2(n278), .ZN(n37) );
  AOI222_X1 U27 ( .A1(D[25]), .A2(n290), .B1(E[25]), .B2(n287), .C1(C[25]), 
        .C2(n284), .ZN(n38) );
  NAND2_X1 U28 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U29 ( .A1(A[28]), .A2(n281), .B1(B[28]), .B2(n278), .ZN(n31) );
  AOI222_X1 U30 ( .A1(D[28]), .A2(n290), .B1(E[28]), .B2(n287), .C1(C[28]), 
        .C2(n284), .ZN(n32) );
  NAND2_X1 U31 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U32 ( .A1(A[29]), .A2(n281), .B1(B[29]), .B2(n278), .ZN(n29) );
  AOI222_X1 U33 ( .A1(D[29]), .A2(n290), .B1(E[29]), .B2(n287), .C1(C[29]), 
        .C2(n284), .ZN(n30) );
  NAND2_X1 U34 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U35 ( .A1(A[30]), .A2(n281), .B1(B[30]), .B2(n278), .ZN(n25) );
  AOI222_X1 U36 ( .A1(D[30]), .A2(n290), .B1(E[30]), .B2(n287), .C1(C[30]), 
        .C2(n284), .ZN(n26) );
  NAND2_X1 U37 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U38 ( .A1(A[31]), .A2(n282), .B1(B[31]), .B2(n279), .ZN(n23) );
  AOI222_X1 U39 ( .A1(D[31]), .A2(n291), .B1(E[31]), .B2(n288), .C1(C[31]), 
        .C2(n285), .ZN(n24) );
  INV_X1 U40 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U41 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U42 ( .A1(A[18]), .A2(n280), .B1(B[18]), .B2(n277), .ZN(n53) );
  AOI222_X1 U43 ( .A1(D[18]), .A2(n289), .B1(E[18]), .B2(n286), .C1(C[18]), 
        .C2(n283), .ZN(n54) );
  NAND2_X1 U44 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U45 ( .A1(A[4]), .A2(n282), .B1(B[4]), .B2(n279), .ZN(n19) );
  AOI222_X1 U46 ( .A1(D[4]), .A2(n291), .B1(E[4]), .B2(n288), .C1(C[4]), .C2(
        n285), .ZN(n20) );
  NAND2_X1 U47 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U48 ( .A1(A[14]), .A2(n280), .B1(B[14]), .B2(n277), .ZN(n61) );
  AOI222_X1 U49 ( .A1(D[14]), .A2(n289), .B1(E[14]), .B2(n286), .C1(C[14]), 
        .C2(n283), .ZN(n62) );
  NAND2_X1 U50 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U51 ( .A1(A[21]), .A2(n281), .B1(B[21]), .B2(n278), .ZN(n45) );
  AOI222_X1 U52 ( .A1(D[21]), .A2(n290), .B1(E[21]), .B2(n287), .C1(C[21]), 
        .C2(n284), .ZN(n46) );
  NAND2_X1 U53 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U54 ( .A1(A[22]), .A2(n281), .B1(B[22]), .B2(n278), .ZN(n43) );
  AOI222_X1 U55 ( .A1(D[22]), .A2(n290), .B1(E[22]), .B2(n287), .C1(C[22]), 
        .C2(n284), .ZN(n44) );
  NAND2_X1 U56 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U57 ( .A1(A[8]), .A2(n282), .B1(B[8]), .B2(n279), .ZN(n11) );
  AOI222_X1 U58 ( .A1(D[8]), .A2(n291), .B1(E[8]), .B2(n288), .C1(C[8]), .C2(
        n285), .ZN(n12) );
  NAND2_X1 U59 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U60 ( .A1(A[5]), .A2(n282), .B1(B[5]), .B2(n279), .ZN(n17) );
  AOI222_X1 U61 ( .A1(D[5]), .A2(n291), .B1(E[5]), .B2(n288), .C1(C[5]), .C2(
        n285), .ZN(n18) );
  NAND2_X1 U62 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U63 ( .A1(A[20]), .A2(n281), .B1(B[20]), .B2(n278), .ZN(n47) );
  AOI222_X1 U64 ( .A1(D[20]), .A2(n290), .B1(E[20]), .B2(n287), .C1(C[20]), 
        .C2(n284), .ZN(n48) );
  NAND2_X1 U65 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U66 ( .A1(A[26]), .A2(n281), .B1(B[26]), .B2(n278), .ZN(n35) );
  AOI222_X1 U67 ( .A1(D[26]), .A2(n290), .B1(E[26]), .B2(n287), .C1(C[26]), 
        .C2(n284), .ZN(n36) );
  NAND2_X1 U68 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U69 ( .A1(A[27]), .A2(n281), .B1(B[27]), .B2(n278), .ZN(n33) );
  AOI222_X1 U70 ( .A1(D[27]), .A2(n290), .B1(E[27]), .B2(n287), .C1(C[27]), 
        .C2(n284), .ZN(n34) );
  NAND2_X1 U71 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U72 ( .A1(A[23]), .A2(n281), .B1(B[23]), .B2(n278), .ZN(n41) );
  AOI222_X1 U73 ( .A1(D[23]), .A2(n290), .B1(E[23]), .B2(n287), .C1(C[23]), 
        .C2(n284), .ZN(n42) );
  NAND2_X1 U74 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U75 ( .A1(A[6]), .A2(n282), .B1(B[6]), .B2(n279), .ZN(n15) );
  AOI222_X1 U76 ( .A1(D[6]), .A2(n291), .B1(E[6]), .B2(n288), .C1(C[6]), .C2(
        n285), .ZN(n16) );
  NAND2_X1 U77 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U78 ( .A1(A[10]), .A2(n280), .B1(B[10]), .B2(n277), .ZN(n69) );
  AOI222_X1 U79 ( .A1(D[10]), .A2(n289), .B1(E[10]), .B2(n286), .C1(C[10]), 
        .C2(n283), .ZN(n70) );
  NAND2_X1 U80 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U81 ( .A1(A[17]), .A2(n280), .B1(B[17]), .B2(n277), .ZN(n55) );
  AOI222_X1 U82 ( .A1(D[17]), .A2(n289), .B1(E[17]), .B2(n286), .C1(C[17]), 
        .C2(n283), .ZN(n56) );
  NAND2_X1 U83 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U84 ( .A1(A[13]), .A2(n280), .B1(B[13]), .B2(n277), .ZN(n63) );
  AOI222_X1 U85 ( .A1(D[13]), .A2(n289), .B1(E[13]), .B2(n286), .C1(C[13]), 
        .C2(n283), .ZN(n64) );
  AND2_X1 U86 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U87 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U88 ( .A1(A[7]), .A2(n282), .B1(B[7]), .B2(n279), .ZN(n13) );
  AOI222_X1 U89 ( .A1(D[7]), .A2(n291), .B1(E[7]), .B2(n288), .C1(C[7]), .C2(
        n285), .ZN(n14) );
  NAND2_X1 U90 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U91 ( .A1(A[9]), .A2(n282), .B1(B[9]), .B2(n279), .ZN(n4) );
  AOI222_X1 U92 ( .A1(D[9]), .A2(n291), .B1(E[9]), .B2(n288), .C1(C[9]), .C2(
        n285), .ZN(n5) );
  NAND2_X1 U93 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U94 ( .A1(A[12]), .A2(n280), .B1(B[12]), .B2(n277), .ZN(n65) );
  AOI222_X1 U95 ( .A1(D[12]), .A2(n289), .B1(E[12]), .B2(n286), .C1(C[12]), 
        .C2(n283), .ZN(n66) );
  NAND2_X1 U96 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U97 ( .A1(A[16]), .A2(n280), .B1(B[16]), .B2(n277), .ZN(n57) );
  AOI222_X1 U98 ( .A1(D[16]), .A2(n289), .B1(E[16]), .B2(n286), .C1(C[16]), 
        .C2(n283), .ZN(n58) );
  NAND2_X1 U99 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U100 ( .A1(A[15]), .A2(n280), .B1(B[15]), .B2(n277), .ZN(n59) );
  AOI222_X1 U101 ( .A1(D[15]), .A2(n289), .B1(E[15]), .B2(n286), .C1(C[15]), 
        .C2(n283), .ZN(n60) );
  NAND2_X1 U102 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U103 ( .A1(A[11]), .A2(n280), .B1(B[11]), .B2(n277), .ZN(n67) );
  AOI222_X1 U104 ( .A1(D[11]), .A2(n289), .B1(E[11]), .B2(n286), .C1(C[11]), 
        .C2(n283), .ZN(n68) );
  NAND2_X1 U105 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U106 ( .A1(A[3]), .A2(n282), .B1(B[3]), .B2(n279), .ZN(n21) );
  AOI222_X1 U107 ( .A1(D[3]), .A2(n291), .B1(E[3]), .B2(n288), .C1(C[3]), .C2(
        n285), .ZN(n22) );
  NAND2_X1 U108 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U109 ( .A1(A[0]), .A2(n280), .B1(B[0]), .B2(n277), .ZN(n71) );
  AOI222_X1 U110 ( .A1(D[0]), .A2(n289), .B1(E[0]), .B2(n286), .C1(C[0]), .C2(
        n283), .ZN(n72) );
  NAND2_X1 U111 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U112 ( .A1(A[1]), .A2(n280), .B1(B[1]), .B2(n277), .ZN(n49) );
  AOI222_X1 U113 ( .A1(D[1]), .A2(n289), .B1(E[1]), .B2(n286), .C1(C[1]), .C2(
        n283), .ZN(n50) );
  NAND2_X1 U114 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U115 ( .A1(A[2]), .A2(n281), .B1(B[2]), .B2(n278), .ZN(n27) );
  AOI222_X1 U116 ( .A1(D[2]), .A2(n290), .B1(E[2]), .B2(n287), .C1(C[2]), .C2(
        n284), .ZN(n28) );
  NAND2_X1 U117 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U118 ( .A1(A[19]), .A2(n280), .B1(B[19]), .B2(n277), .ZN(n51) );
  AOI222_X1 U119 ( .A1(D[19]), .A2(n289), .B1(E[19]), .B2(n286), .C1(C[19]), 
        .C2(n283), .ZN(n52) );
  INV_X1 U120 ( .A(Sel[1]), .ZN(n75) );
endmodule


module mux_N32_7 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339;

  BUF_X1 U1 ( .A(n10), .Z(n325) );
  BUF_X1 U2 ( .A(n10), .Z(n326) );
  BUF_X1 U3 ( .A(n10), .Z(n327) );
  BUF_X1 U4 ( .A(n6), .Z(n337) );
  BUF_X1 U5 ( .A(n6), .Z(n338) );
  BUF_X1 U6 ( .A(n9), .Z(n328) );
  BUF_X1 U7 ( .A(n9), .Z(n329) );
  BUF_X1 U8 ( .A(n7), .Z(n334) );
  BUF_X1 U9 ( .A(n7), .Z(n335) );
  BUF_X1 U10 ( .A(n8), .Z(n331) );
  BUF_X1 U11 ( .A(n8), .Z(n332) );
  BUF_X1 U12 ( .A(n9), .Z(n330) );
  BUF_X1 U13 ( .A(n7), .Z(n336) );
  BUF_X1 U14 ( .A(n8), .Z(n333) );
  BUF_X1 U15 ( .A(n6), .Z(n339) );
  AND2_X1 U16 ( .A1(n73), .A2(n74), .ZN(n10) );
  AOI222_X1 U17 ( .A1(n75), .A2(Sel[0]), .B1(n76), .B2(Sel[2]), .C1(n74), .C2(
        Sel[1]), .ZN(n9) );
  NOR3_X1 U18 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n74), .ZN(n7) );
  NOR3_X1 U19 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n76), .B(Sel[1]), .ZN(n73) );
  INV_X1 U21 ( .A(Sel[0]), .ZN(n76) );
  INV_X1 U22 ( .A(Sel[2]), .ZN(n74) );
  NAND2_X1 U23 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U24 ( .A1(A[16]), .A2(n328), .B1(B[16]), .B2(n325), .ZN(n57) );
  AOI222_X1 U25 ( .A1(D[16]), .A2(n337), .B1(E[16]), .B2(n334), .C1(C[16]), 
        .C2(n331), .ZN(n58) );
  NAND2_X1 U26 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U27 ( .A1(A[2]), .A2(n329), .B1(B[2]), .B2(n326), .ZN(n27) );
  AOI222_X1 U28 ( .A1(D[2]), .A2(n338), .B1(E[2]), .B2(n335), .C1(C[2]), .C2(
        n332), .ZN(n28) );
  NAND2_X1 U29 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U30 ( .A1(A[12]), .A2(n328), .B1(B[12]), .B2(n325), .ZN(n65) );
  AOI222_X1 U31 ( .A1(D[12]), .A2(n337), .B1(E[12]), .B2(n334), .C1(C[12]), 
        .C2(n331), .ZN(n66) );
  NAND2_X1 U32 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U33 ( .A1(A[6]), .A2(n330), .B1(B[6]), .B2(n327), .ZN(n15) );
  AOI222_X1 U34 ( .A1(D[6]), .A2(n339), .B1(E[6]), .B2(n336), .C1(C[6]), .C2(
        n333), .ZN(n16) );
  NAND2_X1 U35 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U36 ( .A1(A[3]), .A2(n330), .B1(B[3]), .B2(n327), .ZN(n21) );
  AOI222_X1 U37 ( .A1(D[3]), .A2(n339), .B1(E[3]), .B2(n336), .C1(C[3]), .C2(
        n333), .ZN(n22) );
  NAND2_X1 U38 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U39 ( .A1(A[10]), .A2(n328), .B1(B[10]), .B2(n325), .ZN(n69) );
  AOI222_X1 U40 ( .A1(D[10]), .A2(n337), .B1(E[10]), .B2(n334), .C1(C[10]), 
        .C2(n331), .ZN(n70) );
  NAND2_X1 U41 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U42 ( .A1(A[4]), .A2(n330), .B1(B[4]), .B2(n327), .ZN(n19) );
  AOI222_X1 U43 ( .A1(D[4]), .A2(n339), .B1(E[4]), .B2(n336), .C1(C[4]), .C2(
        n333), .ZN(n20) );
  NAND2_X1 U44 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U45 ( .A1(A[8]), .A2(n330), .B1(B[8]), .B2(n327), .ZN(n11) );
  AOI222_X1 U46 ( .A1(D[8]), .A2(n339), .B1(E[8]), .B2(n336), .C1(C[8]), .C2(
        n333), .ZN(n12) );
  NAND2_X1 U47 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U48 ( .A1(A[15]), .A2(n328), .B1(B[15]), .B2(n325), .ZN(n59) );
  AOI222_X1 U49 ( .A1(D[15]), .A2(n337), .B1(E[15]), .B2(n334), .C1(C[15]), 
        .C2(n331), .ZN(n60) );
  NAND2_X1 U50 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U51 ( .A1(A[11]), .A2(n328), .B1(B[11]), .B2(n325), .ZN(n67) );
  AOI222_X1 U52 ( .A1(D[11]), .A2(n337), .B1(E[11]), .B2(n334), .C1(C[11]), 
        .C2(n331), .ZN(n68) );
  AND2_X1 U53 ( .A1(Sel[2]), .A2(n73), .ZN(n8) );
  NAND2_X1 U54 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U55 ( .A1(A[25]), .A2(n329), .B1(B[25]), .B2(n326), .ZN(n37) );
  AOI222_X1 U56 ( .A1(D[25]), .A2(n338), .B1(E[25]), .B2(n335), .C1(C[25]), 
        .C2(n332), .ZN(n38) );
  NAND2_X1 U57 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U58 ( .A1(A[26]), .A2(n329), .B1(B[26]), .B2(n326), .ZN(n35) );
  AOI222_X1 U59 ( .A1(D[26]), .A2(n338), .B1(E[26]), .B2(n335), .C1(C[26]), 
        .C2(n332), .ZN(n36) );
  NAND2_X1 U60 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U61 ( .A1(A[22]), .A2(n329), .B1(B[22]), .B2(n326), .ZN(n43) );
  AOI222_X1 U62 ( .A1(D[22]), .A2(n338), .B1(E[22]), .B2(n335), .C1(C[22]), 
        .C2(n332), .ZN(n44) );
  NAND2_X1 U63 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U64 ( .A1(A[27]), .A2(n329), .B1(B[27]), .B2(n326), .ZN(n33) );
  AOI222_X1 U65 ( .A1(D[27]), .A2(n338), .B1(E[27]), .B2(n335), .C1(C[27]), 
        .C2(n332), .ZN(n34) );
  NAND2_X1 U66 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U67 ( .A1(A[19]), .A2(n328), .B1(B[19]), .B2(n325), .ZN(n51) );
  AOI222_X1 U68 ( .A1(D[19]), .A2(n337), .B1(E[19]), .B2(n334), .C1(C[19]), 
        .C2(n331), .ZN(n52) );
  NAND2_X1 U69 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U70 ( .A1(A[28]), .A2(n329), .B1(B[28]), .B2(n326), .ZN(n31) );
  AOI222_X1 U71 ( .A1(D[28]), .A2(n338), .B1(E[28]), .B2(n335), .C1(C[28]), 
        .C2(n332), .ZN(n32) );
  NAND2_X1 U72 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U73 ( .A1(A[29]), .A2(n329), .B1(B[29]), .B2(n326), .ZN(n29) );
  AOI222_X1 U74 ( .A1(D[29]), .A2(n338), .B1(E[29]), .B2(n335), .C1(C[29]), 
        .C2(n332), .ZN(n30) );
  NAND2_X1 U75 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U76 ( .A1(A[5]), .A2(n330), .B1(B[5]), .B2(n327), .ZN(n17) );
  AOI222_X1 U77 ( .A1(D[5]), .A2(n339), .B1(E[5]), .B2(n336), .C1(C[5]), .C2(
        n333), .ZN(n18) );
  NAND2_X1 U78 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U79 ( .A1(A[9]), .A2(n330), .B1(B[9]), .B2(n327), .ZN(n4) );
  AOI222_X1 U80 ( .A1(D[9]), .A2(n339), .B1(E[9]), .B2(n336), .C1(C[9]), .C2(
        n333), .ZN(n5) );
  NAND2_X1 U81 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U82 ( .A1(A[7]), .A2(n330), .B1(B[7]), .B2(n327), .ZN(n13) );
  AOI222_X1 U83 ( .A1(D[7]), .A2(n339), .B1(E[7]), .B2(n336), .C1(C[7]), .C2(
        n333), .ZN(n14) );
  NAND2_X1 U84 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U85 ( .A1(A[13]), .A2(n328), .B1(B[13]), .B2(n325), .ZN(n63) );
  AOI222_X1 U86 ( .A1(D[13]), .A2(n337), .B1(E[13]), .B2(n334), .C1(C[13]), 
        .C2(n331), .ZN(n64) );
  NAND2_X1 U87 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U88 ( .A1(A[17]), .A2(n328), .B1(B[17]), .B2(n325), .ZN(n55) );
  AOI222_X1 U89 ( .A1(D[17]), .A2(n337), .B1(E[17]), .B2(n334), .C1(C[17]), 
        .C2(n331), .ZN(n56) );
  NAND2_X1 U90 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U91 ( .A1(A[14]), .A2(n328), .B1(B[14]), .B2(n325), .ZN(n61) );
  AOI222_X1 U92 ( .A1(D[14]), .A2(n337), .B1(E[14]), .B2(n334), .C1(C[14]), 
        .C2(n331), .ZN(n62) );
  NAND2_X1 U93 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U94 ( .A1(A[23]), .A2(n329), .B1(B[23]), .B2(n326), .ZN(n41) );
  AOI222_X1 U95 ( .A1(D[23]), .A2(n338), .B1(E[23]), .B2(n335), .C1(C[23]), 
        .C2(n332), .ZN(n42) );
  NAND2_X1 U96 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U97 ( .A1(A[24]), .A2(n329), .B1(B[24]), .B2(n326), .ZN(n39) );
  AOI222_X1 U98 ( .A1(D[24]), .A2(n338), .B1(E[24]), .B2(n335), .C1(C[24]), 
        .C2(n332), .ZN(n40) );
  NAND2_X1 U99 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U100 ( .A1(A[20]), .A2(n329), .B1(B[20]), .B2(n326), .ZN(n47) );
  AOI222_X1 U101 ( .A1(D[20]), .A2(n338), .B1(E[20]), .B2(n335), .C1(C[20]), 
        .C2(n332), .ZN(n48) );
  NAND2_X1 U102 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U103 ( .A1(A[21]), .A2(n329), .B1(B[21]), .B2(n326), .ZN(n45) );
  AOI222_X1 U104 ( .A1(D[21]), .A2(n338), .B1(E[21]), .B2(n335), .C1(C[21]), 
        .C2(n332), .ZN(n46) );
  NAND2_X1 U105 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U106 ( .A1(A[18]), .A2(n328), .B1(B[18]), .B2(n325), .ZN(n53) );
  AOI222_X1 U107 ( .A1(D[18]), .A2(n337), .B1(E[18]), .B2(n334), .C1(C[18]), 
        .C2(n331), .ZN(n54) );
  NAND2_X1 U108 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U109 ( .A1(A[30]), .A2(n329), .B1(B[30]), .B2(n326), .ZN(n25) );
  AOI222_X1 U110 ( .A1(D[30]), .A2(n338), .B1(E[30]), .B2(n335), .C1(C[30]), 
        .C2(n332), .ZN(n26) );
  NAND2_X1 U111 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U112 ( .A1(A[31]), .A2(n330), .B1(B[31]), .B2(n327), .ZN(n23) );
  AOI222_X1 U113 ( .A1(D[31]), .A2(n339), .B1(E[31]), .B2(n336), .C1(C[31]), 
        .C2(n333), .ZN(n24) );
  INV_X1 U114 ( .A(Sel[1]), .ZN(n75) );
  NAND2_X1 U115 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U116 ( .A1(A[0]), .A2(n328), .B1(B[0]), .B2(n325), .ZN(n71) );
  AOI222_X1 U117 ( .A1(D[0]), .A2(n337), .B1(E[0]), .B2(n334), .C1(C[0]), .C2(
        n331), .ZN(n72) );
  NAND2_X1 U118 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U119 ( .A1(A[1]), .A2(n328), .B1(B[1]), .B2(n325), .ZN(n49) );
  AOI222_X1 U120 ( .A1(D[1]), .A2(n337), .B1(E[1]), .B2(n334), .C1(C[1]), .C2(
        n331), .ZN(n50) );
endmodule


module mux_N32_0 ( A, B, C, D, E, Sel, O );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] Sel;
  output [31:0] O;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286;

  OAI33_X1 U105 ( .A1(n73), .A2(n75), .A3(n76), .B1(Sel[0]), .B2(Sel[2]), .B3(
        Sel[1]), .ZN(n9) );
  BUF_X1 U1 ( .A(n10), .Z(n272) );
  BUF_X1 U2 ( .A(n10), .Z(n273) );
  BUF_X1 U3 ( .A(n10), .Z(n274) );
  BUF_X1 U4 ( .A(n6), .Z(n284) );
  BUF_X1 U5 ( .A(n6), .Z(n285) );
  BUF_X1 U6 ( .A(n9), .Z(n275) );
  BUF_X1 U7 ( .A(n9), .Z(n276) );
  BUF_X1 U8 ( .A(n7), .Z(n281) );
  BUF_X1 U9 ( .A(n7), .Z(n282) );
  BUF_X1 U10 ( .A(n9), .Z(n277) );
  BUF_X1 U11 ( .A(n8), .Z(n278) );
  BUF_X1 U12 ( .A(n8), .Z(n279) );
  BUF_X1 U13 ( .A(n7), .Z(n283) );
  BUF_X1 U14 ( .A(n8), .Z(n280) );
  BUF_X1 U15 ( .A(n6), .Z(n286) );
  AND2_X1 U16 ( .A1(n74), .A2(n73), .ZN(n10) );
  NOR3_X1 U17 ( .A1(Sel[0]), .A2(Sel[1]), .A3(n73), .ZN(n8) );
  NOR3_X1 U18 ( .A1(n75), .A2(Sel[2]), .A3(n76), .ZN(n6) );
  XNOR2_X1 U19 ( .A(n76), .B(Sel[1]), .ZN(n74) );
  NAND2_X1 U20 ( .A1(n61), .A2(n62), .ZN(O[14]) );
  AOI22_X1 U21 ( .A1(A[14]), .A2(n275), .B1(B[14]), .B2(n272), .ZN(n61) );
  AOI222_X1 U22 ( .A1(D[14]), .A2(n284), .B1(C[14]), .B2(n281), .C1(E[14]), 
        .C2(n278), .ZN(n62) );
  NAND2_X1 U23 ( .A1(n49), .A2(n50), .ZN(O[1]) );
  AOI22_X1 U24 ( .A1(A[1]), .A2(n275), .B1(B[1]), .B2(n272), .ZN(n49) );
  AOI222_X1 U25 ( .A1(D[1]), .A2(n284), .B1(C[1]), .B2(n281), .C1(E[1]), .C2(
        n278), .ZN(n50) );
  NAND2_X1 U26 ( .A1(n69), .A2(n70), .ZN(O[10]) );
  AOI22_X1 U27 ( .A1(A[10]), .A2(n275), .B1(B[10]), .B2(n272), .ZN(n69) );
  AOI222_X1 U28 ( .A1(D[10]), .A2(n284), .B1(C[10]), .B2(n281), .C1(E[10]), 
        .C2(n278), .ZN(n70) );
  NAND2_X1 U29 ( .A1(n19), .A2(n20), .ZN(O[4]) );
  AOI22_X1 U30 ( .A1(A[4]), .A2(n277), .B1(B[4]), .B2(n274), .ZN(n19) );
  AOI222_X1 U31 ( .A1(D[4]), .A2(n286), .B1(C[4]), .B2(n283), .C1(E[4]), .C2(
        n280), .ZN(n20) );
  NAND2_X1 U32 ( .A1(n71), .A2(n72), .ZN(O[0]) );
  AOI22_X1 U33 ( .A1(A[0]), .A2(n275), .B1(B[0]), .B2(n272), .ZN(n71) );
  AOI222_X1 U34 ( .A1(D[0]), .A2(n284), .B1(C[0]), .B2(n281), .C1(E[0]), .C2(
        n278), .ZN(n72) );
  NAND2_X1 U35 ( .A1(n11), .A2(n12), .ZN(O[8]) );
  AOI22_X1 U36 ( .A1(A[8]), .A2(n277), .B1(B[8]), .B2(n274), .ZN(n11) );
  AOI222_X1 U37 ( .A1(D[8]), .A2(n286), .B1(C[8]), .B2(n283), .C1(E[8]), .C2(
        n280), .ZN(n12) );
  NAND2_X1 U38 ( .A1(n27), .A2(n28), .ZN(O[2]) );
  AOI22_X1 U39 ( .A1(A[2]), .A2(n276), .B1(B[2]), .B2(n273), .ZN(n27) );
  AOI222_X1 U40 ( .A1(D[2]), .A2(n285), .B1(C[2]), .B2(n282), .C1(E[2]), .C2(
        n279), .ZN(n28) );
  INV_X1 U41 ( .A(Sel[2]), .ZN(n73) );
  NAND2_X1 U42 ( .A1(n63), .A2(n64), .ZN(O[13]) );
  AOI22_X1 U43 ( .A1(A[13]), .A2(n275), .B1(B[13]), .B2(n272), .ZN(n63) );
  AOI222_X1 U44 ( .A1(D[13]), .A2(n284), .B1(C[13]), .B2(n281), .C1(E[13]), 
        .C2(n278), .ZN(n64) );
  NAND2_X1 U45 ( .A1(n4), .A2(n5), .ZN(O[9]) );
  AOI22_X1 U46 ( .A1(A[9]), .A2(n277), .B1(B[9]), .B2(n274), .ZN(n4) );
  AOI222_X1 U47 ( .A1(D[9]), .A2(n286), .B1(C[9]), .B2(n283), .C1(E[9]), .C2(
        n280), .ZN(n5) );
  AND2_X1 U48 ( .A1(Sel[2]), .A2(n74), .ZN(n7) );
  NAND2_X1 U49 ( .A1(n21), .A2(n22), .ZN(O[3]) );
  AOI22_X1 U50 ( .A1(A[3]), .A2(n277), .B1(B[3]), .B2(n274), .ZN(n21) );
  AOI222_X1 U51 ( .A1(D[3]), .A2(n286), .B1(C[3]), .B2(n283), .C1(E[3]), .C2(
        n280), .ZN(n22) );
  NAND2_X1 U52 ( .A1(n13), .A2(n14), .ZN(O[7]) );
  AOI22_X1 U53 ( .A1(A[7]), .A2(n277), .B1(B[7]), .B2(n274), .ZN(n13) );
  AOI222_X1 U54 ( .A1(D[7]), .A2(n286), .B1(C[7]), .B2(n283), .C1(E[7]), .C2(
        n280), .ZN(n14) );
  NAND2_X1 U55 ( .A1(n59), .A2(n60), .ZN(O[15]) );
  AOI22_X1 U56 ( .A1(A[15]), .A2(n275), .B1(B[15]), .B2(n272), .ZN(n59) );
  AOI222_X1 U57 ( .A1(D[15]), .A2(n284), .B1(C[15]), .B2(n281), .C1(E[15]), 
        .C2(n278), .ZN(n60) );
  NAND2_X1 U58 ( .A1(n67), .A2(n68), .ZN(O[11]) );
  AOI22_X1 U59 ( .A1(A[11]), .A2(n275), .B1(B[11]), .B2(n272), .ZN(n67) );
  AOI222_X1 U60 ( .A1(D[11]), .A2(n284), .B1(C[11]), .B2(n281), .C1(E[11]), 
        .C2(n278), .ZN(n68) );
  NAND2_X1 U61 ( .A1(n65), .A2(n66), .ZN(O[12]) );
  AOI22_X1 U62 ( .A1(A[12]), .A2(n275), .B1(B[12]), .B2(n272), .ZN(n65) );
  AOI222_X1 U63 ( .A1(D[12]), .A2(n284), .B1(C[12]), .B2(n281), .C1(E[12]), 
        .C2(n278), .ZN(n66) );
  NAND2_X1 U64 ( .A1(n15), .A2(n16), .ZN(O[6]) );
  AOI22_X1 U65 ( .A1(A[6]), .A2(n277), .B1(B[6]), .B2(n274), .ZN(n15) );
  AOI222_X1 U66 ( .A1(D[6]), .A2(n286), .B1(C[6]), .B2(n283), .C1(E[6]), .C2(
        n280), .ZN(n16) );
  NAND2_X1 U67 ( .A1(n39), .A2(n40), .ZN(O[24]) );
  AOI22_X1 U68 ( .A1(A[24]), .A2(n276), .B1(B[24]), .B2(n273), .ZN(n39) );
  AOI222_X1 U69 ( .A1(D[24]), .A2(n285), .B1(C[24]), .B2(n282), .C1(E[24]), 
        .C2(n279), .ZN(n40) );
  NAND2_X1 U70 ( .A1(n47), .A2(n48), .ZN(O[20]) );
  AOI22_X1 U71 ( .A1(A[20]), .A2(n276), .B1(B[20]), .B2(n273), .ZN(n47) );
  AOI222_X1 U72 ( .A1(D[20]), .A2(n285), .B1(C[20]), .B2(n282), .C1(E[20]), 
        .C2(n279), .ZN(n48) );
  NAND2_X1 U73 ( .A1(n37), .A2(n38), .ZN(O[25]) );
  AOI22_X1 U74 ( .A1(A[25]), .A2(n276), .B1(B[25]), .B2(n273), .ZN(n37) );
  AOI222_X1 U75 ( .A1(D[25]), .A2(n285), .B1(C[25]), .B2(n282), .C1(E[25]), 
        .C2(n279), .ZN(n38) );
  NAND2_X1 U76 ( .A1(n45), .A2(n46), .ZN(O[21]) );
  AOI22_X1 U77 ( .A1(A[21]), .A2(n276), .B1(B[21]), .B2(n273), .ZN(n45) );
  AOI222_X1 U78 ( .A1(D[21]), .A2(n285), .B1(C[21]), .B2(n282), .C1(E[21]), 
        .C2(n279), .ZN(n46) );
  NAND2_X1 U79 ( .A1(n55), .A2(n56), .ZN(O[17]) );
  AOI22_X1 U80 ( .A1(A[17]), .A2(n275), .B1(B[17]), .B2(n272), .ZN(n55) );
  AOI222_X1 U81 ( .A1(D[17]), .A2(n284), .B1(C[17]), .B2(n281), .C1(E[17]), 
        .C2(n278), .ZN(n56) );
  NAND2_X1 U82 ( .A1(n35), .A2(n36), .ZN(O[26]) );
  AOI22_X1 U83 ( .A1(A[26]), .A2(n276), .B1(B[26]), .B2(n273), .ZN(n35) );
  AOI222_X1 U84 ( .A1(D[26]), .A2(n285), .B1(C[26]), .B2(n282), .C1(E[26]), 
        .C2(n279), .ZN(n36) );
  NAND2_X1 U85 ( .A1(n43), .A2(n44), .ZN(O[22]) );
  AOI22_X1 U86 ( .A1(A[22]), .A2(n276), .B1(B[22]), .B2(n273), .ZN(n43) );
  AOI222_X1 U87 ( .A1(D[22]), .A2(n285), .B1(C[22]), .B2(n282), .C1(E[22]), 
        .C2(n279), .ZN(n44) );
  NAND2_X1 U88 ( .A1(n53), .A2(n54), .ZN(O[18]) );
  AOI22_X1 U89 ( .A1(A[18]), .A2(n275), .B1(B[18]), .B2(n272), .ZN(n53) );
  AOI222_X1 U90 ( .A1(D[18]), .A2(n284), .B1(C[18]), .B2(n281), .C1(E[18]), 
        .C2(n278), .ZN(n54) );
  NAND2_X1 U91 ( .A1(n33), .A2(n34), .ZN(O[27]) );
  AOI22_X1 U92 ( .A1(A[27]), .A2(n276), .B1(B[27]), .B2(n273), .ZN(n33) );
  AOI222_X1 U93 ( .A1(D[27]), .A2(n285), .B1(C[27]), .B2(n282), .C1(E[27]), 
        .C2(n279), .ZN(n34) );
  NAND2_X1 U94 ( .A1(n41), .A2(n42), .ZN(O[23]) );
  AOI22_X1 U95 ( .A1(A[23]), .A2(n276), .B1(B[23]), .B2(n273), .ZN(n41) );
  AOI222_X1 U96 ( .A1(D[23]), .A2(n285), .B1(C[23]), .B2(n282), .C1(E[23]), 
        .C2(n279), .ZN(n42) );
  NAND2_X1 U97 ( .A1(n51), .A2(n52), .ZN(O[19]) );
  AOI22_X1 U98 ( .A1(A[19]), .A2(n275), .B1(B[19]), .B2(n272), .ZN(n51) );
  AOI222_X1 U99 ( .A1(D[19]), .A2(n284), .B1(C[19]), .B2(n281), .C1(E[19]), 
        .C2(n278), .ZN(n52) );
  NAND2_X1 U100 ( .A1(n31), .A2(n32), .ZN(O[28]) );
  AOI22_X1 U101 ( .A1(A[28]), .A2(n276), .B1(B[28]), .B2(n273), .ZN(n31) );
  AOI222_X1 U102 ( .A1(D[28]), .A2(n285), .B1(C[28]), .B2(n282), .C1(E[28]), 
        .C2(n279), .ZN(n32) );
  NAND2_X1 U103 ( .A1(n29), .A2(n30), .ZN(O[29]) );
  AOI22_X1 U104 ( .A1(A[29]), .A2(n276), .B1(B[29]), .B2(n273), .ZN(n29) );
  AOI222_X1 U106 ( .A1(D[29]), .A2(n285), .B1(C[29]), .B2(n282), .C1(E[29]), 
        .C2(n279), .ZN(n30) );
  NAND2_X1 U107 ( .A1(n25), .A2(n26), .ZN(O[30]) );
  AOI22_X1 U108 ( .A1(A[30]), .A2(n276), .B1(B[30]), .B2(n273), .ZN(n25) );
  AOI222_X1 U109 ( .A1(D[30]), .A2(n285), .B1(C[30]), .B2(n282), .C1(E[30]), 
        .C2(n279), .ZN(n26) );
  NAND2_X1 U110 ( .A1(n23), .A2(n24), .ZN(O[31]) );
  AOI22_X1 U111 ( .A1(A[31]), .A2(n277), .B1(B[31]), .B2(n274), .ZN(n23) );
  AOI222_X1 U112 ( .A1(D[31]), .A2(n286), .B1(C[31]), .B2(n283), .C1(E[31]), 
        .C2(n280), .ZN(n24) );
  NAND2_X1 U113 ( .A1(n57), .A2(n58), .ZN(O[16]) );
  AOI22_X1 U114 ( .A1(A[16]), .A2(n275), .B1(B[16]), .B2(n272), .ZN(n57) );
  AOI222_X1 U115 ( .A1(D[16]), .A2(n284), .B1(C[16]), .B2(n281), .C1(E[16]), 
        .C2(n278), .ZN(n58) );
  NAND2_X1 U116 ( .A1(n17), .A2(n18), .ZN(O[5]) );
  AOI22_X1 U117 ( .A1(A[5]), .A2(n277), .B1(B[5]), .B2(n274), .ZN(n17) );
  AOI222_X1 U118 ( .A1(D[5]), .A2(n286), .B1(C[5]), .B2(n283), .C1(E[5]), .C2(
        n280), .ZN(n18) );
  INV_X1 U119 ( .A(Sel[1]), .ZN(n75) );
  INV_X1 U120 ( .A(Sel[0]), .ZN(n76) );
endmodule


module shift_mul_N16_S14 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[14] , \A[13] , \A[11] , \A[9] , \A[7] , \A[5] , \A[4] , \A[3] ,
         \A[2] , \A[1] , \E[31] , \E[30] , \E[29] , \E[28] , \E[27] , \E[26] ,
         \E[25] , \E[24] , \E[23] , \E[22] , \E[21] , \E[20] , \E[19] ,
         \E[18] , \E[17] , \E[16] , \A[0] , \A[15] , n9, n10, n12, n13, n14,
         n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n62, n63, \D[21] ,
         n65, \D[23] , n67, \D[25] , n69, \D[27] , n71, n72;
  assign B[13] = 1'b0;
  assign B[12] = 1'b0;
  assign B[11] = 1'b0;
  assign B[10] = 1'b0;
  assign B[9] = 1'b0;
  assign B[8] = 1'b0;
  assign B[7] = 1'b0;
  assign B[6] = 1'b0;
  assign B[5] = 1'b0;
  assign B[4] = 1'b0;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[13] = 1'b0;
  assign C[12] = 1'b0;
  assign C[11] = 1'b0;
  assign C[10] = 1'b0;
  assign C[9] = 1'b0;
  assign C[8] = 1'b0;
  assign C[7] = 1'b0;
  assign C[6] = 1'b0;
  assign C[5] = 1'b0;
  assign C[4] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[14] = 1'b0;
  assign D[13] = 1'b0;
  assign D[12] = 1'b0;
  assign D[11] = 1'b0;
  assign D[10] = 1'b0;
  assign D[9] = 1'b0;
  assign D[8] = 1'b0;
  assign D[7] = 1'b0;
  assign D[6] = 1'b0;
  assign D[5] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[14] = 1'b0;
  assign E[13] = 1'b0;
  assign E[12] = 1'b0;
  assign E[11] = 1'b0;
  assign E[10] = 1'b0;
  assign E[9] = 1'b0;
  assign E[8] = 1'b0;
  assign E[7] = 1'b0;
  assign E[6] = 1'b0;
  assign E[5] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[28] = \A[14] ;
  assign D[29] = \A[14] ;
  assign \A[14]  = A[14];
  assign B[27] = \A[13] ;
  assign D[28] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[25] = \A[11] ;
  assign D[26] = \A[11] ;
  assign \A[11]  = A[11];
  assign B[23] = \A[9] ;
  assign D[24] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[21] = \A[7] ;
  assign D[22] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[19] = \A[5] ;
  assign D[20] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[18] = \A[4] ;
  assign D[19] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[17] = \A[3] ;
  assign D[18] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[16] = \A[2] ;
  assign D[17] = \A[2] ;
  assign \A[2]  = A[2];
  assign B[15] = \A[1] ;
  assign D[16] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[31] = \E[31] ;
  assign C[30] = \E[31] ;
  assign E[31] = \E[31] ;
  assign C[29] = \E[30] ;
  assign E[30] = \E[30] ;
  assign C[28] = \E[29] ;
  assign E[29] = \E[29] ;
  assign C[27] = \E[28] ;
  assign E[28] = \E[28] ;
  assign C[26] = \E[27] ;
  assign E[27] = \E[27] ;
  assign C[25] = \E[26] ;
  assign E[26] = \E[26] ;
  assign C[24] = \E[25] ;
  assign E[25] = \E[25] ;
  assign C[23] = \E[24] ;
  assign E[24] = \E[24] ;
  assign C[22] = \E[23] ;
  assign E[23] = \E[23] ;
  assign C[21] = \E[22] ;
  assign E[22] = \E[22] ;
  assign C[20] = \E[21] ;
  assign E[21] = \E[21] ;
  assign C[19] = \E[20] ;
  assign E[20] = \E[20] ;
  assign C[18] = \E[19] ;
  assign E[19] = \E[19] ;
  assign C[17] = \E[18] ;
  assign E[18] = \E[18] ;
  assign C[16] = \E[17] ;
  assign E[17] = \E[17] ;
  assign C[15] = \E[16] ;
  assign E[16] = \E[16] ;
  assign B[14] = \A[0] ;
  assign C[14] = \A[0] ;
  assign D[15] = \A[0] ;
  assign E[15] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[31] = \A[15] ;
  assign B[30] = \A[15] ;
  assign B[29] = \A[15] ;
  assign D[31] = \A[15] ;
  assign D[30] = \A[15] ;
  assign \A[15]  = A[15];
  assign B[20] = \D[21] ;
  assign D[21] = \D[21] ;
  assign B[22] = \D[23] ;
  assign D[23] = \D[23] ;
  assign B[24] = \D[25] ;
  assign D[25] = \D[25] ;
  assign B[26] = \D[27] ;
  assign D[27] = \D[27] ;

  XOR2_X1 U27 ( .A(n12), .B(\A[13] ), .Z(\E[28] ) );
  XOR2_X1 U28 ( .A(n14), .B(n71), .Z(\E[27] ) );
  XOR2_X1 U29 ( .A(n16), .B(\A[11] ), .Z(\E[26] ) );
  XOR2_X1 U30 ( .A(n17), .B(n69), .Z(\E[25] ) );
  XOR2_X1 U31 ( .A(n19), .B(\A[9] ), .Z(\E[24] ) );
  XOR2_X1 U32 ( .A(n20), .B(n67), .Z(\E[23] ) );
  XOR2_X1 U33 ( .A(n22), .B(\A[7] ), .Z(\E[22] ) );
  XOR2_X1 U34 ( .A(n23), .B(n65), .Z(\E[21] ) );
  XOR2_X1 U35 ( .A(n25), .B(\A[5] ), .Z(\E[20] ) );
  XOR2_X1 U36 ( .A(n26), .B(n63), .Z(\E[19] ) );
  XOR2_X1 U37 ( .A(n28), .B(\A[3] ), .Z(\E[18] ) );
  XOR2_X1 U38 ( .A(n29), .B(n62), .Z(\E[17] ) );
  XOR2_X1 U39 ( .A(\A[1] ), .B(\A[0] ), .Z(\E[16] ) );
  INV_X1 U2 ( .A(n9), .ZN(\E[31] ) );
  OAI21_X1 U3 ( .B1(n10), .B2(n72), .A(n9), .ZN(\E[30] ) );
  NAND2_X1 U4 ( .A1(n14), .A2(n71), .ZN(n12) );
  NAND2_X1 U5 ( .A1(n17), .A2(n69), .ZN(n16) );
  NAND2_X1 U6 ( .A1(n72), .A2(n10), .ZN(n9) );
  NAND2_X1 U7 ( .A1(n26), .A2(n63), .ZN(n25) );
  NAND2_X1 U8 ( .A1(n20), .A2(n67), .ZN(n19) );
  NAND2_X1 U9 ( .A1(n23), .A2(n65), .ZN(n22) );
  NOR2_X1 U10 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n29) );
  XNOR2_X1 U11 ( .A(\A[14] ), .B(n13), .ZN(\E[29] ) );
  NOR2_X1 U12 ( .A1(\A[13] ), .A2(n12), .ZN(n13) );
  NOR2_X1 U13 ( .A1(n19), .A2(\A[9] ), .ZN(n17) );
  NOR2_X1 U14 ( .A1(n28), .A2(\A[3] ), .ZN(n26) );
  NOR2_X1 U15 ( .A1(n22), .A2(\A[7] ), .ZN(n20) );
  NOR2_X1 U16 ( .A1(n25), .A2(\A[5] ), .ZN(n23) );
  NOR2_X1 U17 ( .A1(n16), .A2(\A[11] ), .ZN(n14) );
  INV_X1 U18 ( .A(A[8]), .ZN(n67) );
  INV_X1 U19 ( .A(A[12]), .ZN(n71) );
  INV_X1 U20 ( .A(A[10]), .ZN(n69) );
  INV_X1 U21 ( .A(A[6]), .ZN(n65) );
  INV_X1 U22 ( .A(\A[4] ), .ZN(n63) );
  INV_X1 U23 ( .A(\A[15] ), .ZN(n72) );
  OR3_X1 U24 ( .A1(\A[13] ), .A2(\A[14] ), .A3(n12), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n29), .A2(n62), .ZN(n28) );
  INV_X1 U26 ( .A(\A[2] ), .ZN(n62) );
  INV_X1 U40 ( .A(n65), .ZN(\D[21] ) );
  INV_X1 U41 ( .A(n67), .ZN(\D[23] ) );
  INV_X1 U42 ( .A(n69), .ZN(\D[25] ) );
  INV_X1 U43 ( .A(n71), .ZN(\D[27] ) );
endmodule


module shift_mul_N16_S12 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[14] , \A[13] , \A[11] , \A[10] , \A[9] , \A[7] , \A[6] , \A[5] ,
         \A[4] , \A[3] , \A[1] , \E[28] , \E[27] , \E[26] , \E[25] , \E[24] ,
         \E[23] , \E[22] , \E[21] , \E[20] , \E[19] , \E[18] , \E[17] ,
         \E[16] , \E[15] , \E[14] , \A[0] , \E[29] , \A[2] , n9, n10, n11, n13,
         n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n66, n67, n68,
         \D[21] , n70, n71, \D[25] , n73, n74, \D[28] ;
  assign B[11] = 1'b0;
  assign B[10] = 1'b0;
  assign B[9] = 1'b0;
  assign B[8] = 1'b0;
  assign B[7] = 1'b0;
  assign B[6] = 1'b0;
  assign B[5] = 1'b0;
  assign B[4] = 1'b0;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[11] = 1'b0;
  assign C[10] = 1'b0;
  assign C[9] = 1'b0;
  assign C[8] = 1'b0;
  assign C[7] = 1'b0;
  assign C[6] = 1'b0;
  assign C[5] = 1'b0;
  assign C[4] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[12] = 1'b0;
  assign D[11] = 1'b0;
  assign D[10] = 1'b0;
  assign D[9] = 1'b0;
  assign D[8] = 1'b0;
  assign D[7] = 1'b0;
  assign D[6] = 1'b0;
  assign D[5] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[12] = 1'b0;
  assign E[11] = 1'b0;
  assign E[10] = 1'b0;
  assign E[9] = 1'b0;
  assign E[8] = 1'b0;
  assign E[7] = 1'b0;
  assign E[6] = 1'b0;
  assign E[5] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[26] = \A[14] ;
  assign D[27] = \A[14] ;
  assign \A[14]  = A[14];
  assign B[25] = \A[13] ;
  assign D[26] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[23] = \A[11] ;
  assign D[24] = \A[11] ;
  assign \A[11]  = A[11];
  assign B[22] = \A[10] ;
  assign D[23] = \A[10] ;
  assign \A[10]  = A[10];
  assign B[21] = \A[9] ;
  assign D[22] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[19] = \A[7] ;
  assign D[20] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[18] = \A[6] ;
  assign D[19] = \A[6] ;
  assign \A[6]  = A[6];
  assign B[17] = \A[5] ;
  assign D[18] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[16] = \A[4] ;
  assign D[17] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[15] = \A[3] ;
  assign D[16] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[13] = \A[1] ;
  assign D[14] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[27] = \E[28] ;
  assign E[28] = \E[28] ;
  assign C[26] = \E[27] ;
  assign E[27] = \E[27] ;
  assign C[25] = \E[26] ;
  assign E[26] = \E[26] ;
  assign C[24] = \E[25] ;
  assign E[25] = \E[25] ;
  assign C[23] = \E[24] ;
  assign E[24] = \E[24] ;
  assign C[22] = \E[23] ;
  assign E[23] = \E[23] ;
  assign C[21] = \E[22] ;
  assign E[22] = \E[22] ;
  assign C[20] = \E[21] ;
  assign E[21] = \E[21] ;
  assign C[19] = \E[20] ;
  assign E[20] = \E[20] ;
  assign C[18] = \E[19] ;
  assign E[19] = \E[19] ;
  assign C[17] = \E[18] ;
  assign E[18] = \E[18] ;
  assign C[16] = \E[17] ;
  assign E[17] = \E[17] ;
  assign C[15] = \E[16] ;
  assign E[16] = \E[16] ;
  assign C[14] = \E[15] ;
  assign E[15] = \E[15] ;
  assign C[13] = \E[14] ;
  assign E[14] = \E[14] ;
  assign B[12] = \A[0] ;
  assign C[12] = \A[0] ;
  assign D[13] = \A[0] ;
  assign E[13] = \A[0] ;
  assign \A[0]  = A[0];
  assign C[31] = \E[29] ;
  assign C[30] = \E[29] ;
  assign C[29] = \E[29] ;
  assign C[28] = \E[29] ;
  assign E[31] = \E[29] ;
  assign E[30] = \E[29] ;
  assign E[29] = \E[29] ;
  assign B[14] = \A[2] ;
  assign D[15] = \A[2] ;
  assign \A[2]  = A[2];
  assign B[20] = \D[21] ;
  assign D[21] = \D[21] ;
  assign B[24] = \D[25] ;
  assign D[25] = \D[25] ;
  assign B[27] = \D[28] ;
  assign B[31] = \D[28] ;
  assign B[28] = \D[28] ;
  assign B[30] = \D[28] ;
  assign B[29] = \D[28] ;
  assign D[31] = \D[28] ;
  assign D[29] = \D[28] ;
  assign D[30] = \D[28] ;
  assign D[28] = \D[28] ;

  NAND3_X1 U25 ( .A1(n11), .A2(n74), .A3(\D[28] ), .ZN(n10) );
  XOR2_X1 U26 ( .A(n11), .B(n74), .Z(\E[27] ) );
  XOR2_X1 U27 ( .A(n13), .B(\A[13] ), .Z(\E[26] ) );
  XOR2_X1 U28 ( .A(n14), .B(n73), .Z(\E[25] ) );
  XOR2_X1 U29 ( .A(n16), .B(\A[11] ), .Z(\E[24] ) );
  XOR2_X1 U30 ( .A(n17), .B(n71), .Z(\E[23] ) );
  XOR2_X1 U31 ( .A(n19), .B(\A[9] ), .Z(\E[22] ) );
  XOR2_X1 U32 ( .A(n20), .B(n70), .Z(\E[21] ) );
  XOR2_X1 U33 ( .A(n22), .B(\A[7] ), .Z(\E[20] ) );
  XOR2_X1 U34 ( .A(n23), .B(n68), .Z(\E[19] ) );
  XOR2_X1 U35 ( .A(n25), .B(\A[5] ), .Z(\E[18] ) );
  XOR2_X1 U36 ( .A(n26), .B(n67), .Z(\E[17] ) );
  XOR2_X1 U37 ( .A(n28), .B(\A[3] ), .Z(\E[16] ) );
  XOR2_X1 U38 ( .A(n29), .B(n66), .Z(\E[15] ) );
  XOR2_X1 U39 ( .A(\A[1] ), .B(\A[0] ), .Z(\E[14] ) );
  AOI21_X1 U2 ( .B1(n74), .B2(n11), .A(\D[28] ), .ZN(\E[29] ) );
  NAND2_X1 U3 ( .A1(n9), .A2(n10), .ZN(\E[28] ) );
  INV_X1 U4 ( .A(\E[29] ), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n17), .A2(n71), .ZN(n16) );
  NAND2_X1 U6 ( .A1(n26), .A2(n67), .ZN(n25) );
  NAND2_X1 U7 ( .A1(n20), .A2(n70), .ZN(n19) );
  NAND2_X1 U8 ( .A1(n23), .A2(n68), .ZN(n22) );
  NAND2_X1 U9 ( .A1(n14), .A2(n73), .ZN(n13) );
  NOR2_X1 U10 ( .A1(n13), .A2(\A[13] ), .ZN(n11) );
  NOR2_X1 U11 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n29) );
  NOR2_X1 U12 ( .A1(n19), .A2(\A[9] ), .ZN(n17) );
  BUF_X1 U13 ( .A(A[15]), .Z(\D[28] ) );
  NOR2_X1 U14 ( .A1(n28), .A2(\A[3] ), .ZN(n26) );
  NOR2_X1 U15 ( .A1(n22), .A2(\A[7] ), .ZN(n20) );
  NOR2_X1 U16 ( .A1(n25), .A2(\A[5] ), .ZN(n23) );
  NOR2_X1 U17 ( .A1(n16), .A2(\A[11] ), .ZN(n14) );
  INV_X1 U18 ( .A(A[8]), .ZN(n70) );
  INV_X1 U19 ( .A(A[12]), .ZN(n73) );
  INV_X1 U20 ( .A(\A[10] ), .ZN(n71) );
  INV_X1 U21 ( .A(\A[6] ), .ZN(n68) );
  INV_X1 U22 ( .A(\A[4] ), .ZN(n67) );
  NAND2_X1 U23 ( .A1(n29), .A2(n66), .ZN(n28) );
  INV_X1 U24 ( .A(\A[2] ), .ZN(n66) );
  INV_X1 U40 ( .A(n70), .ZN(\D[21] ) );
  INV_X1 U41 ( .A(n73), .ZN(\D[25] ) );
  INV_X1 U42 ( .A(\A[14] ), .ZN(n74) );
endmodule


module shift_mul_N16_S10 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[8] , \A[7] , \A[5] ,
         \A[4] , \A[3] , \A[1] , \E[25] , \E[24] , \E[23] , \E[22] , \E[21] ,
         \E[20] , \E[19] , \E[18] , \E[17] , \E[16] , \E[15] , \E[14] ,
         \E[13] , \E[12] , \A[9] , \A[6] , \A[0] , \A[2] , \E[26] , \E[27] ,
         n9, n10, n12, n13, n14, n16, n17, n19, n20, n22, n23, n25, n26, n28,
         n29, n81, n82, n83, n84, n85, n86, \D[26] , n88;
  assign B[9] = 1'b0;
  assign B[8] = 1'b0;
  assign B[7] = 1'b0;
  assign B[6] = 1'b0;
  assign B[5] = 1'b0;
  assign B[4] = 1'b0;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[9] = 1'b0;
  assign C[8] = 1'b0;
  assign C[7] = 1'b0;
  assign C[6] = 1'b0;
  assign C[5] = 1'b0;
  assign C[4] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[10] = 1'b0;
  assign D[9] = 1'b0;
  assign D[8] = 1'b0;
  assign D[7] = 1'b0;
  assign D[6] = 1'b0;
  assign D[5] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[10] = 1'b0;
  assign E[9] = 1'b0;
  assign E[8] = 1'b0;
  assign E[7] = 1'b0;
  assign E[6] = 1'b0;
  assign E[5] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[24] = \A[14] ;
  assign D[25] = \A[14] ;
  assign \A[14]  = A[14];
  assign B[23] = \A[13] ;
  assign D[24] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[22] = \A[12] ;
  assign D[23] = \A[12] ;
  assign \A[12]  = A[12];
  assign B[21] = \A[11] ;
  assign D[22] = \A[11] ;
  assign \A[11]  = A[11];
  assign B[20] = \A[10] ;
  assign D[21] = \A[10] ;
  assign \A[10]  = A[10];
  assign B[18] = \A[8] ;
  assign D[19] = \A[8] ;
  assign \A[8]  = A[8];
  assign B[17] = \A[7] ;
  assign D[18] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[15] = \A[5] ;
  assign D[16] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[14] = \A[4] ;
  assign D[15] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[13] = \A[3] ;
  assign D[14] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[11] = \A[1] ;
  assign D[12] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[24] = \E[25] ;
  assign E[25] = \E[25] ;
  assign C[23] = \E[24] ;
  assign E[24] = \E[24] ;
  assign C[22] = \E[23] ;
  assign E[23] = \E[23] ;
  assign C[21] = \E[22] ;
  assign E[22] = \E[22] ;
  assign C[20] = \E[21] ;
  assign E[21] = \E[21] ;
  assign C[19] = \E[20] ;
  assign E[20] = \E[20] ;
  assign C[18] = \E[19] ;
  assign E[19] = \E[19] ;
  assign C[17] = \E[18] ;
  assign E[18] = \E[18] ;
  assign C[16] = \E[17] ;
  assign E[17] = \E[17] ;
  assign C[15] = \E[16] ;
  assign E[16] = \E[16] ;
  assign C[14] = \E[15] ;
  assign E[15] = \E[15] ;
  assign C[13] = \E[14] ;
  assign E[14] = \E[14] ;
  assign C[12] = \E[13] ;
  assign E[13] = \E[13] ;
  assign C[11] = \E[12] ;
  assign E[12] = \E[12] ;
  assign B[19] = \A[9] ;
  assign D[20] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[16] = \A[6] ;
  assign D[17] = \A[6] ;
  assign \A[6]  = A[6];
  assign B[10] = \A[0] ;
  assign C[10] = \A[0] ;
  assign D[11] = \A[0] ;
  assign E[11] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[12] = \A[2] ;
  assign D[13] = \A[2] ;
  assign \A[2]  = A[2];
  assign C[25] = \E[26] ;
  assign E[26] = \E[26] ;
  assign C[31] = \E[27] ;
  assign C[30] = \E[27] ;
  assign C[29] = \E[27] ;
  assign C[28] = \E[27] ;
  assign C[27] = \E[27] ;
  assign C[26] = \E[27] ;
  assign E[31] = \E[27] ;
  assign E[30] = \E[27] ;
  assign E[29] = \E[27] ;
  assign E[28] = \E[27] ;
  assign E[27] = \E[27] ;
  assign B[31] = \D[26] ;
  assign B[30] = \D[26] ;
  assign B[29] = \D[26] ;
  assign B[28] = \D[26] ;
  assign B[27] = \D[26] ;
  assign B[26] = \D[26] ;
  assign B[25] = \D[26] ;
  assign D[31] = \D[26] ;
  assign D[30] = \D[26] ;
  assign D[29] = \D[26] ;
  assign D[28] = \D[26] ;
  assign D[27] = \D[26] ;
  assign D[26] = \D[26] ;

  XOR2_X1 U27 ( .A(n12), .B(\A[13] ), .Z(\E[24] ) );
  XOR2_X1 U28 ( .A(n14), .B(n86), .Z(\E[23] ) );
  XOR2_X1 U29 ( .A(n16), .B(\A[11] ), .Z(\E[22] ) );
  XOR2_X1 U30 ( .A(n17), .B(n85), .Z(\E[21] ) );
  XOR2_X1 U31 ( .A(n19), .B(\A[9] ), .Z(\E[20] ) );
  XOR2_X1 U32 ( .A(n20), .B(n84), .Z(\E[19] ) );
  XOR2_X1 U33 ( .A(n22), .B(\A[7] ), .Z(\E[18] ) );
  XOR2_X1 U34 ( .A(n23), .B(n83), .Z(\E[17] ) );
  XOR2_X1 U35 ( .A(n25), .B(\A[5] ), .Z(\E[16] ) );
  XOR2_X1 U36 ( .A(n26), .B(n82), .Z(\E[15] ) );
  XOR2_X1 U37 ( .A(n28), .B(\A[3] ), .Z(\E[14] ) );
  XOR2_X1 U38 ( .A(n29), .B(n81), .Z(\E[13] ) );
  XOR2_X1 U39 ( .A(\A[1] ), .B(\A[0] ), .Z(\E[12] ) );
  INV_X1 U2 ( .A(n9), .ZN(\E[27] ) );
  INV_X1 U3 ( .A(n88), .ZN(\D[26] ) );
  OAI21_X1 U4 ( .B1(n10), .B2(n88), .A(n9), .ZN(\E[26] ) );
  NAND2_X1 U5 ( .A1(n14), .A2(n86), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n17), .A2(n85), .ZN(n16) );
  NAND2_X1 U7 ( .A1(n88), .A2(n10), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n26), .A2(n82), .ZN(n25) );
  NAND2_X1 U9 ( .A1(n20), .A2(n84), .ZN(n19) );
  NAND2_X1 U10 ( .A1(n23), .A2(n83), .ZN(n22) );
  NOR2_X1 U11 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n29) );
  XNOR2_X1 U12 ( .A(\A[14] ), .B(n13), .ZN(\E[25] ) );
  NOR2_X1 U13 ( .A1(\A[13] ), .A2(n12), .ZN(n13) );
  NOR2_X1 U14 ( .A1(n19), .A2(\A[9] ), .ZN(n17) );
  NOR2_X1 U15 ( .A1(n28), .A2(\A[3] ), .ZN(n26) );
  NOR2_X1 U16 ( .A1(n22), .A2(\A[7] ), .ZN(n20) );
  NOR2_X1 U17 ( .A1(n25), .A2(\A[5] ), .ZN(n23) );
  NOR2_X1 U18 ( .A1(n16), .A2(\A[11] ), .ZN(n14) );
  INV_X1 U19 ( .A(\A[8] ), .ZN(n84) );
  INV_X1 U20 ( .A(\A[12] ), .ZN(n86) );
  INV_X1 U21 ( .A(\A[10] ), .ZN(n85) );
  INV_X1 U22 ( .A(\A[6] ), .ZN(n83) );
  INV_X1 U23 ( .A(\A[4] ), .ZN(n82) );
  INV_X1 U24 ( .A(A[15]), .ZN(n88) );
  OR3_X1 U25 ( .A1(\A[13] ), .A2(\A[14] ), .A3(n12), .ZN(n10) );
  NAND2_X1 U26 ( .A1(n29), .A2(n81), .ZN(n28) );
  INV_X1 U40 ( .A(\A[2] ), .ZN(n81) );
endmodule


module shift_mul_N16_S8 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[13] , \A[12] , \A[8] , \A[7] , \A[5] , \A[3] , \A[1] , \E[25] ,
         \A[9] , \A[10] , \A[0] , \E[24] , n7, n8, n9, n11, n13, n15, n17, n18,
         n19, n21, n22, n24, n25, n95, n96, \D[11] , n98, \D[13] , n100,
         \D[15] , n102, \D[20] , n104, \D[23] , n106, \D[24] , \B[27] ;
  assign B[7] = 1'b0;
  assign B[6] = 1'b0;
  assign B[5] = 1'b0;
  assign B[4] = 1'b0;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[7] = 1'b0;
  assign C[6] = 1'b0;
  assign C[5] = 1'b0;
  assign C[4] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[8] = 1'b0;
  assign D[7] = 1'b0;
  assign D[6] = 1'b0;
  assign D[5] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[8] = 1'b0;
  assign E[7] = 1'b0;
  assign E[6] = 1'b0;
  assign E[5] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[21] = \A[13] ;
  assign D[22] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[20] = \A[12] ;
  assign D[21] = \A[12] ;
  assign \A[12]  = A[12];
  assign B[16] = \A[8] ;
  assign D[17] = \A[8] ;
  assign \A[8]  = A[8];
  assign B[15] = \A[7] ;
  assign D[16] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[13] = \A[5] ;
  assign D[14] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[11] = \A[3] ;
  assign D[12] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[9] = \A[1] ;
  assign D[10] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[22] = E[23];
  assign C[21] = E[22];
  assign C[20] = E[21];
  assign C[19] = E[20];
  assign C[18] = E[19];
  assign C[17] = E[18];
  assign C[16] = E[17];
  assign C[15] = E[16];
  assign C[14] = E[15];
  assign C[13] = E[14];
  assign C[12] = E[13];
  assign C[11] = E[12];
  assign C[10] = E[11];
  assign C[9] = E[10];
  assign C[31] = \E[25] ;
  assign C[30] = \E[25] ;
  assign C[29] = \E[25] ;
  assign C[28] = \E[25] ;
  assign C[27] = \E[25] ;
  assign C[26] = \E[25] ;
  assign C[25] = \E[25] ;
  assign C[24] = \E[25] ;
  assign E[31] = \E[25] ;
  assign E[30] = \E[25] ;
  assign E[29] = \E[25] ;
  assign E[28] = \E[25] ;
  assign E[27] = \E[25] ;
  assign E[26] = \E[25] ;
  assign E[25] = \E[25] ;
  assign B[17] = \A[9] ;
  assign D[18] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[18] = \A[10] ;
  assign D[19] = \A[10] ;
  assign \A[10]  = A[10];
  assign B[8] = \A[0] ;
  assign C[8] = \A[0] ;
  assign D[9] = \A[0] ;
  assign E[9] = \A[0] ;
  assign \A[0]  = A[0];
  assign C[23] = \E[24] ;
  assign E[24] = \E[24] ;
  assign B[10] = \D[11] ;
  assign D[11] = \D[11] ;
  assign B[12] = \D[13] ;
  assign D[13] = \D[13] ;
  assign B[14] = \D[15] ;
  assign D[15] = \D[15] ;
  assign B[19] = \D[20] ;
  assign D[20] = \D[20] ;
  assign B[22] = \D[23] ;
  assign D[23] = \D[23] ;
  assign B[26] = \D[24] ;
  assign B[25] = \D[24] ;
  assign B[24] = \D[24] ;
  assign B[23] = \D[24] ;
  assign D[31] = \D[24] ;
  assign D[30] = \D[24] ;
  assign D[29] = \D[24] ;
  assign D[28] = \D[24] ;
  assign D[27] = \D[24] ;
  assign D[26] = \D[24] ;
  assign D[25] = \D[24] ;
  assign D[24] = \D[24] ;
  assign B[31] = \B[27] ;
  assign B[30] = \B[27] ;
  assign B[29] = \B[27] ;
  assign B[28] = \B[27] ;
  assign B[27] = \B[27] ;

  NAND3_X1 U29 ( .A1(n9), .A2(n106), .A3(\B[27] ), .ZN(n8) );
  XOR2_X1 U31 ( .A(n11), .B(\A[12] ), .Z(E[21]) );
  XOR2_X1 U33 ( .A(n15), .B(\A[9] ), .Z(E[18]) );
  XOR2_X1 U34 ( .A(n17), .B(\A[7] ), .Z(E[16]) );
  XOR2_X1 U35 ( .A(n21), .B(\A[5] ), .Z(E[14]) );
  XOR2_X1 U36 ( .A(n24), .B(\A[3] ), .Z(E[12]) );
  XOR2_X1 U37 ( .A(\A[1] ), .B(\A[0] ), .Z(E[10]) );
  AOI21_X2 U2 ( .B1(n106), .B2(n9), .A(\B[27] ), .ZN(\E[25] ) );
  XNOR2_X1 U3 ( .A(n9), .B(\D[23] ), .ZN(E[23]) );
  XNOR2_X1 U4 ( .A(n13), .B(\D[20] ), .ZN(E[20]) );
  XNOR2_X1 U5 ( .A(n22), .B(\D[13] ), .ZN(E[13]) );
  XNOR2_X1 U6 ( .A(n25), .B(\D[11] ), .ZN(E[11]) );
  XNOR2_X1 U7 ( .A(n19), .B(\D[15] ), .ZN(E[15]) );
  NAND2_X1 U8 ( .A1(n13), .A2(n104), .ZN(n11) );
  NAND2_X1 U9 ( .A1(n19), .A2(n102), .ZN(n17) );
  NAND2_X1 U10 ( .A1(n7), .A2(n8), .ZN(\E[24] ) );
  INV_X1 U11 ( .A(\E[25] ), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n22), .A2(n100), .ZN(n21) );
  NOR3_X1 U13 ( .A1(\A[12] ), .A2(\A[13] ), .A3(n11), .ZN(n9) );
  XNOR2_X1 U14 ( .A(n95), .B(\A[13] ), .ZN(E[22]) );
  NOR2_X1 U15 ( .A1(n11), .A2(\A[12] ), .ZN(n95) );
  NOR3_X1 U16 ( .A1(\A[10] ), .A2(\A[9] ), .A3(n15), .ZN(n13) );
  XNOR2_X1 U17 ( .A(n96), .B(\A[10] ), .ZN(E[19]) );
  NOR2_X1 U18 ( .A1(n15), .A2(\A[9] ), .ZN(n96) );
  NOR2_X1 U19 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n25) );
  BUF_X1 U20 ( .A(A[15]), .Z(\D[24] ) );
  XNOR2_X1 U21 ( .A(\A[8] ), .B(n18), .ZN(E[17]) );
  NOR2_X1 U22 ( .A1(\A[7] ), .A2(n17), .ZN(n18) );
  NOR2_X1 U23 ( .A1(n24), .A2(\A[3] ), .ZN(n22) );
  NOR2_X1 U24 ( .A1(n21), .A2(\A[5] ), .ZN(n19) );
  BUF_X1 U25 ( .A(A[15]), .Z(\B[27] ) );
  NAND2_X1 U26 ( .A1(n25), .A2(n98), .ZN(n24) );
  OR3_X1 U27 ( .A1(\A[7] ), .A2(\A[8] ), .A3(n17), .ZN(n15) );
  INV_X1 U28 ( .A(n98), .ZN(\D[11] ) );
  INV_X1 U30 ( .A(A[2]), .ZN(n98) );
  INV_X1 U32 ( .A(n100), .ZN(\D[13] ) );
  INV_X1 U38 ( .A(A[4]), .ZN(n100) );
  INV_X1 U39 ( .A(n102), .ZN(\D[15] ) );
  INV_X1 U40 ( .A(A[6]), .ZN(n102) );
  INV_X1 U41 ( .A(n104), .ZN(\D[20] ) );
  INV_X1 U42 ( .A(A[11]), .ZN(n104) );
  INV_X1 U43 ( .A(n106), .ZN(\D[23] ) );
  INV_X1 U44 ( .A(A[14]), .ZN(n106) );
endmodule


module shift_mul_N16_S6 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[14] , \A[13] , \A[12] , \A[10] , \A[9] , \A[7] , \A[6] , \A[5] ,
         \A[4] , \A[3] , \A[2] , \A[1] , \E[21] , \E[20] , \E[19] , \E[18] ,
         \E[17] , \E[16] , \E[15] , \E[14] , \E[13] , \E[12] , \E[11] ,
         \E[10] , \E[9] , \E[8] , \A[0] , \E[23]_snps_wire , \A[8] , \E[22] ,
         n4, n6, n7, n9, n10, n11, n13, n15, n16, n17, n19, n20, n87, n88, n89,
         n90, \E[26] , \E[30] , \C[31] , \C[30] , \C[24] , \C[28] , \C[22] ,
         \C[26] , \E[27] , \D[18] , n101, n102, \D[22] , \B[23] ;
  assign B[5] = 1'b0;
  assign B[4] = 1'b0;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[5] = 1'b0;
  assign C[4] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[6] = 1'b0;
  assign D[5] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[6] = 1'b0;
  assign E[5] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[20] = \A[14] ;
  assign D[21] = \A[14] ;
  assign \A[14]  = A[14];
  assign B[19] = \A[13] ;
  assign D[20] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[18] = \A[12] ;
  assign D[19] = \A[12] ;
  assign \A[12]  = A[12];
  assign B[16] = \A[10] ;
  assign D[17] = \A[10] ;
  assign \A[10]  = A[10];
  assign B[15] = \A[9] ;
  assign D[16] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[13] = \A[7] ;
  assign D[14] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[12] = \A[6] ;
  assign D[13] = \A[6] ;
  assign \A[6]  = A[6];
  assign B[11] = \A[5] ;
  assign D[12] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[10] = \A[4] ;
  assign D[11] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[9] = \A[3] ;
  assign D[10] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[8] = \A[2] ;
  assign D[9] = \A[2] ;
  assign \A[2]  = A[2];
  assign B[7] = \A[1] ;
  assign D[8] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[20] = \E[21] ;
  assign E[21] = \E[21] ;
  assign C[19] = \E[20] ;
  assign E[20] = \E[20] ;
  assign C[18] = \E[19] ;
  assign E[19] = \E[19] ;
  assign C[17] = \E[18] ;
  assign E[18] = \E[18] ;
  assign C[16] = \E[17] ;
  assign E[17] = \E[17] ;
  assign C[15] = \E[16] ;
  assign E[16] = \E[16] ;
  assign C[14] = \E[15] ;
  assign E[15] = \E[15] ;
  assign C[13] = \E[14] ;
  assign E[14] = \E[14] ;
  assign C[12] = \E[13] ;
  assign E[13] = \E[13] ;
  assign C[11] = \E[12] ;
  assign E[12] = \E[12] ;
  assign C[10] = \E[11] ;
  assign E[11] = \E[11] ;
  assign C[9] = \E[10] ;
  assign E[10] = \E[10] ;
  assign C[8] = \E[9] ;
  assign E[9] = \E[9] ;
  assign C[7] = \E[8] ;
  assign E[8] = \E[8] ;
  assign B[6] = \A[0] ;
  assign C[6] = \A[0] ;
  assign D[7] = \A[0] ;
  assign E[7] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[14] = \A[8] ;
  assign D[15] = \A[8] ;
  assign \A[8]  = A[8];
  assign C[21] = \E[22] ;
  assign E[22] = \E[22] ;
  assign C[25] = \E[26] ;
  assign E[29] = \E[26] ;
  assign E[26] = \E[26] ;
  assign E[25] = \E[30] ;
  assign E[30] = \E[30] ;
  assign E[24] = \C[31] ;
  assign C[31] = \C[31] ;
  assign E[23] = \C[30] ;
  assign C[30] = \C[30] ;
  assign C[29] = \C[24] ;
  assign C[24] = \C[24] ;
  assign C[23] = \C[28] ;
  assign C[28] = \C[28] ;
  assign C[27] = \C[22] ;
  assign C[22] = \C[22] ;
  assign E[31] = \C[26] ;
  assign C[26] = \C[26] ;
  assign E[28] = \E[27] ;
  assign E[27] = \E[27] ;
  assign B[17] = \D[18] ;
  assign D[18] = \D[18] ;
  assign B[22] = \D[22] ;
  assign B[21] = \D[22] ;
  assign D[31] = \D[22] ;
  assign D[30] = \D[22] ;
  assign D[29] = \D[22] ;
  assign D[28] = \D[22] ;
  assign D[27] = \D[22] ;
  assign D[26] = \D[22] ;
  assign D[25] = \D[22] ;
  assign D[24] = \D[22] ;
  assign D[23] = \D[22] ;
  assign D[22] = \D[22] ;
  assign B[31] = \B[23] ;
  assign B[30] = \B[23] ;
  assign B[29] = \B[23] ;
  assign B[28] = \B[23] ;
  assign B[27] = \B[23] ;
  assign B[26] = \B[23] ;
  assign B[25] = \B[23] ;
  assign B[24] = \B[23] ;
  assign B[23] = \B[23] ;

  XOR2_X1 U24 ( .A(n4), .B(\A[2] ), .Z(\E[9] ) );
  XOR2_X1 U25 ( .A(\A[1] ), .B(\A[0] ), .Z(\E[8] ) );
  NAND3_X1 U26 ( .A1(n7), .A2(n102), .A3(\B[23] ), .ZN(n6) );
  XOR2_X1 U27 ( .A(n9), .B(\A[13] ), .Z(\E[20] ) );
  XOR2_X1 U28 ( .A(n10), .B(\A[12] ), .Z(\E[19] ) );
  XOR2_X1 U30 ( .A(n13), .B(\A[9] ), .Z(\E[16] ) );
  XOR2_X1 U31 ( .A(n15), .B(\A[7] ), .Z(\E[14] ) );
  XOR2_X1 U33 ( .A(n17), .B(\A[5] ), .Z(\E[12] ) );
  XOR2_X1 U34 ( .A(n19), .B(\A[3] ), .Z(\E[10] ) );
  AOI21_X1 U2 ( .B1(n102), .B2(n7), .A(\B[23] ), .ZN(\E[23]_snps_wire ) );
  XNOR2_X1 U3 ( .A(n7), .B(\A[14] ), .ZN(\E[21] ) );
  XNOR2_X1 U4 ( .A(n11), .B(\D[18] ), .ZN(\E[18] ) );
  NAND2_X1 U5 ( .A1(n11), .A2(n101), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n90), .A2(n6), .ZN(\E[22] ) );
  NOR3_X1 U7 ( .A1(\A[10] ), .A2(\A[9] ), .A3(n13), .ZN(n11) );
  XNOR2_X1 U8 ( .A(n87), .B(\A[10] ), .ZN(\E[17] ) );
  NOR2_X1 U9 ( .A1(n13), .A2(\A[9] ), .ZN(n87) );
  XNOR2_X1 U10 ( .A(n88), .B(\A[6] ), .ZN(\E[13] ) );
  NOR2_X1 U11 ( .A1(n17), .A2(\A[5] ), .ZN(n88) );
  NOR2_X1 U12 ( .A1(n9), .A2(\A[13] ), .ZN(n7) );
  BUF_X1 U13 ( .A(A[15]), .Z(\D[22] ) );
  XNOR2_X1 U14 ( .A(\A[8] ), .B(n16), .ZN(\E[15] ) );
  NOR2_X1 U15 ( .A1(\A[7] ), .A2(n15), .ZN(n16) );
  BUF_X1 U16 ( .A(A[15]), .Z(\B[23] ) );
  XNOR2_X1 U17 ( .A(\A[4] ), .B(n20), .ZN(\E[11] ) );
  NOR2_X1 U18 ( .A1(\A[3] ), .A2(n19), .ZN(n20) );
  OR3_X1 U19 ( .A1(\A[3] ), .A2(\A[4] ), .A3(n19), .ZN(n17) );
  OR3_X1 U20 ( .A1(\A[5] ), .A2(\A[6] ), .A3(n17), .ZN(n15) );
  OR3_X1 U21 ( .A1(\A[7] ), .A2(\A[8] ), .A3(n15), .ZN(n13) );
  OR2_X1 U22 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n4) );
  OR2_X1 U23 ( .A1(n10), .A2(\A[12] ), .ZN(n9) );
  OR2_X1 U29 ( .A1(n4), .A2(\A[2] ), .ZN(n19) );
  INV_X1 U32 ( .A(\E[23]_snps_wire ), .ZN(n89) );
  INV_X1 U35 ( .A(\E[23]_snps_wire ), .ZN(n90) );
  INV_X1 U36 ( .A(n89), .ZN(\E[26] ) );
  INV_X1 U37 ( .A(n89), .ZN(\E[30] ) );
  INV_X1 U38 ( .A(n89), .ZN(\C[31] ) );
  INV_X1 U39 ( .A(n89), .ZN(\C[30] ) );
  INV_X1 U40 ( .A(n90), .ZN(\C[24] ) );
  INV_X1 U41 ( .A(n90), .ZN(\C[28] ) );
  INV_X1 U42 ( .A(n90), .ZN(\C[22] ) );
  INV_X1 U43 ( .A(n90), .ZN(\C[26] ) );
  INV_X1 U44 ( .A(n89), .ZN(\E[27] ) );
  INV_X1 U45 ( .A(n101), .ZN(\D[18] ) );
  INV_X1 U46 ( .A(A[11]), .ZN(n101) );
  INV_X1 U47 ( .A(\A[14] ), .ZN(n102) );
endmodule


module shift_mul_N16_S4 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[13] , \A[12] , \A[10] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] ,
         \A[3] , \A[2] , \A[1] , \E[20] , \E[19] , \E[18] , \E[17] , \E[16] ,
         \E[15] , \E[14] , \E[13] , \E[12] , \E[11] , \E[10] , \E[9] , \E[8] ,
         \E[7] , \E[6] , \A[0] , \A[11] , \A[9] , \E[23] , \E[21] , n6, n7, n8,
         n10, n12, n13, n14, n15, n16, n19, n21, n22, n24, n25, n105, n106,
         n107, n108, n109, \D[19] , n111, \D[20] , \B[19] , n114;
  assign B[3] = 1'b0;
  assign B[2] = 1'b0;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[3] = 1'b0;
  assign C[2] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[4] = 1'b0;
  assign D[3] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[4] = 1'b0;
  assign E[3] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[17] = \A[13] ;
  assign D[18] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[16] = \A[12] ;
  assign D[17] = \A[12] ;
  assign \A[12]  = A[12];
  assign B[14] = \A[10] ;
  assign D[15] = \A[10] ;
  assign \A[10]  = A[10];
  assign B[12] = \A[8] ;
  assign D[13] = \A[8] ;
  assign \A[8]  = A[8];
  assign B[11] = \A[7] ;
  assign D[12] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[10] = \A[6] ;
  assign D[11] = \A[6] ;
  assign \A[6]  = A[6];
  assign B[9] = \A[5] ;
  assign D[10] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[8] = \A[4] ;
  assign D[9] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[7] = \A[3] ;
  assign D[8] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[6] = \A[2] ;
  assign D[7] = \A[2] ;
  assign \A[2]  = A[2];
  assign B[5] = \A[1] ;
  assign D[6] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[19] = \E[20] ;
  assign E[20] = \E[20] ;
  assign C[18] = \E[19] ;
  assign E[19] = \E[19] ;
  assign C[17] = \E[18] ;
  assign E[18] = \E[18] ;
  assign C[16] = \E[17] ;
  assign E[17] = \E[17] ;
  assign C[15] = \E[16] ;
  assign E[16] = \E[16] ;
  assign C[14] = \E[15] ;
  assign E[15] = \E[15] ;
  assign C[13] = \E[14] ;
  assign E[14] = \E[14] ;
  assign C[12] = \E[13] ;
  assign E[13] = \E[13] ;
  assign C[11] = \E[12] ;
  assign E[12] = \E[12] ;
  assign C[10] = \E[11] ;
  assign E[11] = \E[11] ;
  assign C[9] = \E[10] ;
  assign E[10] = \E[10] ;
  assign C[8] = \E[9] ;
  assign E[9] = \E[9] ;
  assign C[7] = \E[8] ;
  assign E[8] = \E[8] ;
  assign C[6] = \E[7] ;
  assign E[7] = \E[7] ;
  assign C[5] = \E[6] ;
  assign E[6] = \E[6] ;
  assign B[4] = \A[0] ;
  assign C[4] = \A[0] ;
  assign D[5] = \A[0] ;
  assign E[5] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[15] = \A[11] ;
  assign D[16] = \A[11] ;
  assign \A[11]  = A[11];
  assign B[13] = \A[9] ;
  assign D[14] = \A[9] ;
  assign \A[9]  = A[9];
  assign C[27] = \E[23] ;
  assign C[26] = \E[23] ;
  assign C[23] = \E[23] ;
  assign C[22] = \E[23] ;
  assign C[21] = \E[23] ;
  assign C[20] = \E[23] ;
  assign E[31] = \E[23] ;
  assign E[30] = \E[23] ;
  assign E[29] = \E[23] ;
  assign E[27] = \E[23] ;
  assign E[26] = \E[23] ;
  assign E[25] = \E[23] ;
  assign E[24] = \E[23] ;
  assign E[23] = \E[23] ;
  assign C[31] = \E[21] ;
  assign C[30] = \E[21] ;
  assign C[29] = \E[21] ;
  assign C[28] = \E[21] ;
  assign C[25] = \E[21] ;
  assign C[24] = \E[21] ;
  assign E[28] = \E[21] ;
  assign E[22] = \E[21] ;
  assign E[21] = \E[21] ;
  assign B[18] = \D[19] ;
  assign D[19] = \D[19] ;
  assign D[31] = \D[20] ;
  assign D[30] = \D[20] ;
  assign D[29] = \D[20] ;
  assign D[28] = \D[20] ;
  assign D[27] = \D[20] ;
  assign D[26] = \D[20] ;
  assign D[25] = \D[20] ;
  assign D[24] = \D[20] ;
  assign D[23] = \D[20] ;
  assign D[22] = \D[20] ;
  assign D[21] = \D[20] ;
  assign D[20] = \D[20] ;
  assign B[30] = \B[19] ;
  assign B[29] = \B[19] ;
  assign B[28] = \B[19] ;
  assign B[27] = \B[19] ;
  assign B[31] = \B[19] ;
  assign B[25] = \B[19] ;
  assign B[24] = \B[19] ;
  assign B[23] = \B[19] ;
  assign B[22] = \B[19] ;
  assign B[21] = \B[19] ;
  assign B[20] = \B[19] ;
  assign B[26] = \B[19] ;
  assign B[19] = \B[19] ;

  XOR2_X1 U26 ( .A(n6), .B(\A[4] ), .Z(\E[9] ) );
  XOR2_X1 U27 ( .A(n7), .B(\A[3] ), .Z(\E[8] ) );
  XOR2_X1 U28 ( .A(n8), .B(n107), .Z(\E[7] ) );
  XOR2_X1 U29 ( .A(\A[1] ), .B(\A[0] ), .Z(\E[6] ) );
  NAND3_X1 U30 ( .A1(n14), .A2(n15), .A3(n114), .ZN(n13) );
  XOR2_X1 U32 ( .A(\A[12] ), .B(n16), .Z(\E[17] ) );
  XOR2_X1 U33 ( .A(n15), .B(n109), .Z(\E[16] ) );
  XOR2_X1 U35 ( .A(n19), .B(\A[9] ), .Z(\E[14] ) );
  XOR2_X1 U36 ( .A(n21), .B(\A[8] ), .Z(\E[13] ) );
  XOR2_X1 U37 ( .A(n22), .B(n108), .Z(\E[12] ) );
  XOR2_X1 U38 ( .A(n24), .B(\A[5] ), .Z(\E[10] ) );
  AOI21_X1 U2 ( .B1(n15), .B2(n14), .A(n114), .ZN(\E[21] ) );
  AOI21_X2 U3 ( .B1(n10), .B2(n111), .A(n114), .ZN(\E[23] ) );
  XNOR2_X1 U4 ( .A(n10), .B(\D[19] ), .ZN(\E[19] ) );
  NAND2_X1 U5 ( .A1(n15), .A2(n109), .ZN(n16) );
  NAND2_X1 U6 ( .A1(n22), .A2(n108), .ZN(n21) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(\E[20] ) );
  INV_X1 U8 ( .A(\E[21] ), .ZN(n12) );
  NOR3_X1 U9 ( .A1(\A[10] ), .A2(\A[9] ), .A3(n19), .ZN(n15) );
  NOR3_X1 U10 ( .A1(\A[12] ), .A2(\A[13] ), .A3(n16), .ZN(n10) );
  NOR4_X1 U11 ( .A1(\A[11] ), .A2(\A[12] ), .A3(\A[13] ), .A4(\D[19] ), .ZN(
        n14) );
  XNOR2_X1 U12 ( .A(n105), .B(\A[13] ), .ZN(\E[18] ) );
  NOR2_X1 U13 ( .A1(n16), .A2(\A[12] ), .ZN(n105) );
  XNOR2_X1 U14 ( .A(n106), .B(\A[10] ), .ZN(\E[15] ) );
  NOR2_X1 U15 ( .A1(n19), .A2(\A[9] ), .ZN(n106) );
  NOR3_X1 U16 ( .A1(\A[5] ), .A2(\A[6] ), .A3(n24), .ZN(n22) );
  BUF_X1 U17 ( .A(A[15]), .Z(\B[19] ) );
  BUF_X1 U18 ( .A(A[15]), .Z(\D[20] ) );
  NOR2_X1 U19 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n8) );
  XNOR2_X1 U20 ( .A(\A[6] ), .B(n25), .ZN(\E[11] ) );
  NOR2_X1 U21 ( .A1(\A[5] ), .A2(n24), .ZN(n25) );
  INV_X1 U22 ( .A(\A[7] ), .ZN(n108) );
  INV_X1 U23 ( .A(\A[11] ), .ZN(n109) );
  OR2_X1 U24 ( .A1(n6), .A2(\A[4] ), .ZN(n24) );
  OR2_X1 U25 ( .A1(n21), .A2(\A[8] ), .ZN(n19) );
  BUF_X1 U31 ( .A(A[15]), .Z(n114) );
  NAND2_X1 U34 ( .A1(n8), .A2(n107), .ZN(n7) );
  OR2_X1 U39 ( .A1(n7), .A2(\A[3] ), .ZN(n6) );
  INV_X1 U40 ( .A(\A[2] ), .ZN(n107) );
  INV_X1 U41 ( .A(n111), .ZN(\D[19] ) );
  INV_X1 U42 ( .A(A[14]), .ZN(n111) );
endmodule


module shift_mul_N16_S2 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   \A[14] , \A[13] , \A[11] , \A[9] , \A[8] , \A[7] , \A[4] , \A[3] ,
         \A[1] , \C[22] , \A[2] , \A[0] , \A[5] , \A[6] , n7, n8, n9, n11, n12,
         n15, n16, n17, n18, n19, n20, n21, n23, n24, n26, n27, n28, \E[23] ,
         n118, n119, n120, \D[13] , n122, \D[15] , n124, \D[18] , \D[30] ,
         \B[29] ;
  assign B[1] = 1'b0;
  assign B[0] = 1'b0;
  assign C[1] = 1'b0;
  assign C[0] = 1'b0;
  assign D[2] = 1'b0;
  assign D[1] = 1'b0;
  assign D[0] = 1'b0;
  assign E[2] = 1'b0;
  assign E[1] = 1'b0;
  assign E[0] = 1'b0;
  assign B[16] = \A[14] ;
  assign D[17] = \A[14] ;
  assign \A[14]  = A[14];
  assign B[15] = \A[13] ;
  assign D[16] = \A[13] ;
  assign \A[13]  = A[13];
  assign B[13] = \A[11] ;
  assign D[14] = \A[11] ;
  assign \A[11]  = A[11];
  assign B[11] = \A[9] ;
  assign D[12] = \A[9] ;
  assign \A[9]  = A[9];
  assign B[10] = \A[8] ;
  assign D[11] = \A[8] ;
  assign \A[8]  = A[8];
  assign B[9] = \A[7] ;
  assign D[10] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[6] = \A[4] ;
  assign D[7] = \A[4] ;
  assign \A[4]  = A[4];
  assign B[5] = \A[3] ;
  assign D[6] = \A[3] ;
  assign \A[3]  = A[3];
  assign B[3] = \A[1] ;
  assign D[4] = \A[1] ;
  assign \A[1]  = A[1];
  assign C[17] = E[18];
  assign C[16] = E[17];
  assign C[15] = E[16];
  assign C[14] = E[15];
  assign C[13] = E[14];
  assign C[12] = E[13];
  assign C[11] = E[12];
  assign C[10] = E[11];
  assign C[9] = E[10];
  assign C[8] = E[9];
  assign C[7] = E[8];
  assign C[6] = E[7];
  assign C[5] = E[6];
  assign C[4] = E[5];
  assign C[3] = E[4];
  assign C[31] = \C[22] ;
  assign E[30] = \C[22] ;
  assign E[31] = \C[22] ;
  assign E[28] = \C[22] ;
  assign C[19] = \C[22] ;
  assign C[28] = \C[22] ;
  assign C[27] = \C[22] ;
  assign C[26] = \C[22] ;
  assign C[25] = \C[22] ;
  assign C[29] = \C[22] ;
  assign C[23] = \C[22] ;
  assign C[22] = \C[22] ;
  assign B[4] = \A[2] ;
  assign D[5] = \A[2] ;
  assign \A[2]  = A[2];
  assign B[2] = \A[0] ;
  assign C[2] = \A[0] ;
  assign D[3] = \A[0] ;
  assign E[3] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[7] = \A[5] ;
  assign D[8] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[8] = \A[6] ;
  assign D[9] = \A[6] ;
  assign \A[6]  = A[6];
  assign C[21] = \E[23] ;
  assign C[20] = \E[23] ;
  assign C[24] = \E[23] ;
  assign C[18] = \E[23] ;
  assign C[30] = \E[23] ;
  assign E[29] = \E[23] ;
  assign E[26] = \E[23] ;
  assign E[27] = \E[23] ;
  assign E[24] = \E[23] ;
  assign E[25] = \E[23] ;
  assign E[22] = \E[23] ;
  assign E[21] = \E[23] ;
  assign E[20] = \E[23] ;
  assign E[19] = \E[23] ;
  assign E[23] = \E[23] ;
  assign B[12] = \D[13] ;
  assign D[13] = \D[13] ;
  assign B[14] = \D[15] ;
  assign D[15] = \D[15] ;
  assign D[29] = \D[18] ;
  assign D[28] = \D[18] ;
  assign D[27] = \D[18] ;
  assign D[26] = \D[18] ;
  assign D[25] = \D[18] ;
  assign D[24] = \D[18] ;
  assign D[23] = \D[18] ;
  assign D[22] = \D[18] ;
  assign D[21] = \D[18] ;
  assign D[20] = \D[18] ;
  assign D[19] = \D[18] ;
  assign D[18] = \D[18] ;
  assign B[25] = \D[30] ;
  assign B[24] = \D[30] ;
  assign B[26] = \D[30] ;
  assign B[22] = \D[30] ;
  assign B[21] = \D[30] ;
  assign B[23] = \D[30] ;
  assign B[19] = \D[30] ;
  assign B[18] = \D[30] ;
  assign B[20] = \D[30] ;
  assign B[17] = \D[30] ;
  assign D[31] = \D[30] ;
  assign D[30] = \D[30] ;
  assign B[30] = \B[29] ;
  assign B[31] = \B[29] ;
  assign B[28] = \B[29] ;
  assign B[27] = \B[29] ;
  assign B[29] = \B[29] ;

  XOR2_X1 U27 ( .A(n7), .B(\A[6] ), .Z(E[9]) );
  XOR2_X1 U28 ( .A(n8), .B(\A[5] ), .Z(E[8]) );
  XOR2_X1 U29 ( .A(n9), .B(n120), .Z(E[7]) );
  XOR2_X1 U30 ( .A(n11), .B(\A[3] ), .Z(E[6]) );
  XOR2_X1 U31 ( .A(n12), .B(n119), .Z(E[5]) );
  XOR2_X1 U32 ( .A(\A[1] ), .B(\A[0] ), .Z(E[4]) );
  NAND3_X1 U33 ( .A1(n16), .A2(n17), .A3(\B[29] ), .ZN(n15) );
  XOR2_X1 U34 ( .A(n20), .B(\A[13] ), .Z(E[16]) );
  XOR2_X1 U35 ( .A(n124), .B(n21), .Z(E[15]) );
  XOR2_X1 U36 ( .A(n23), .B(\A[11] ), .Z(E[14]) );
  XOR2_X1 U37 ( .A(n122), .B(n24), .Z(E[13]) );
  XOR2_X1 U38 ( .A(n26), .B(\A[9] ), .Z(E[12]) );
  XOR2_X1 U39 ( .A(n27), .B(\A[7] ), .Z(E[10]) );
  INV_X1 U2 ( .A(n118), .ZN(\E[23] ) );
  INV_X1 U3 ( .A(\C[22] ), .ZN(n118) );
  AOI21_X1 U4 ( .B1(n17), .B2(n16), .A(\B[29] ), .ZN(\C[22] ) );
  NAND2_X1 U5 ( .A1(n118), .A2(n15), .ZN(E[18]) );
  INV_X1 U6 ( .A(n16), .ZN(n26) );
  NAND2_X1 U7 ( .A1(n24), .A2(n122), .ZN(n23) );
  NAND2_X1 U8 ( .A1(n21), .A2(n124), .ZN(n20) );
  NAND2_X1 U9 ( .A1(n9), .A2(n120), .ZN(n8) );
  NOR3_X1 U10 ( .A1(\A[7] ), .A2(\A[8] ), .A3(n27), .ZN(n16) );
  NOR4_X1 U11 ( .A1(\A[11] ), .A2(\D[15] ), .A3(\D[13] ), .A4(n18), .ZN(n17)
         );
  OR3_X1 U12 ( .A1(\A[13] ), .A2(\A[9] ), .A3(\A[14] ), .ZN(n18) );
  BUF_X1 U13 ( .A(A[15]), .Z(\D[18] ) );
  BUF_X1 U14 ( .A(A[15]), .Z(\D[30] ) );
  XNOR2_X1 U15 ( .A(\A[8] ), .B(n28), .ZN(E[11]) );
  NOR2_X1 U16 ( .A1(\A[7] ), .A2(n27), .ZN(n28) );
  NOR2_X1 U17 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n12) );
  XNOR2_X1 U18 ( .A(\A[14] ), .B(n19), .ZN(E[17]) );
  NOR2_X1 U19 ( .A1(\A[13] ), .A2(n20), .ZN(n19) );
  NOR2_X1 U20 ( .A1(n26), .A2(\A[9] ), .ZN(n24) );
  NOR2_X1 U21 ( .A1(n11), .A2(\A[3] ), .ZN(n9) );
  NOR2_X1 U22 ( .A1(n23), .A2(\A[11] ), .ZN(n21) );
  INV_X1 U23 ( .A(A[12]), .ZN(n124) );
  INV_X1 U24 ( .A(A[10]), .ZN(n122) );
  BUF_X1 U25 ( .A(A[15]), .Z(\B[29] ) );
  INV_X1 U26 ( .A(\A[4] ), .ZN(n120) );
  OR2_X1 U40 ( .A1(n7), .A2(\A[6] ), .ZN(n27) );
  NAND2_X1 U41 ( .A1(n12), .A2(n119), .ZN(n11) );
  OR2_X1 U42 ( .A1(n8), .A2(\A[5] ), .ZN(n7) );
  INV_X1 U43 ( .A(\A[2] ), .ZN(n119) );
  INV_X1 U44 ( .A(n122), .ZN(\D[13] ) );
  INV_X1 U45 ( .A(n124), .ZN(\D[15] ) );
endmodule


module shift_mul_N16_S0 ( A, B, C, D, E );
  input [15:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [31:0] E;
  wire   net25272, \A[1] , \A[12] , \E[4] , \A[7] , \A[6] , \A[5] , \A[0] ,
         \A[15] , n6, n8, n9, n10, n11, n12, n13, n14, n16, n18, n19, n21, n22,
         n99, n100, \C[20] , \D[3] , n103, n104, \D[12] , n106, \D[28] , n108;
  assign D[0] = 1'b0;
  assign E[0] = 1'b0;
  assign B[14] = A[14];
  assign D[15] = A[14];
  assign B[13] = A[13];
  assign D[14] = A[13];
  assign B[10] = A[10];
  assign D[11] = A[10];
  assign B[9] = A[9];
  assign D[10] = A[9];
  assign B[8] = A[8];
  assign D[9] = A[8];
  assign B[4] = A[4];
  assign D[5] = A[4];
  assign B[3] = A[3];
  assign D[4] = A[3];
  assign C[15] = E[16];
  assign C[14] = E[15];
  assign C[13] = E[14];
  assign C[12] = E[13];
  assign C[11] = E[12];
  assign C[10] = E[11];
  assign C[9] = E[10];
  assign C[8] = E[9];
  assign C[7] = E[8];
  assign C[6] = E[7];
  assign C[5] = E[6];
  assign C[4] = E[5];
  assign C[2] = E[3];
  assign C[1] = E[2];
  assign B[1] = \A[1] ;
  assign D[2] = \A[1] ;
  assign \A[1]  = A[1];
  assign B[12] = \A[12] ;
  assign D[13] = \A[12] ;
  assign \A[12]  = A[12];
  assign C[3] = \E[4] ;
  assign E[4] = \E[4] ;
  assign B[7] = \A[7] ;
  assign D[8] = \A[7] ;
  assign \A[7]  = A[7];
  assign B[6] = \A[6] ;
  assign D[7] = \A[6] ;
  assign \A[6]  = A[6];
  assign B[5] = \A[5] ;
  assign D[6] = \A[5] ;
  assign \A[5]  = A[5];
  assign B[0] = \A[0] ;
  assign C[0] = \A[0] ;
  assign D[1] = \A[0] ;
  assign E[1] = \A[0] ;
  assign \A[0]  = A[0];
  assign B[31] = \A[15] ;
  assign B[27] = \A[15] ;
  assign D[27] = \A[15] ;
  assign D[25] = \A[15] ;
  assign D[23] = \A[15] ;
  assign D[21] = \A[15] ;
  assign D[19] = \A[15] ;
  assign D[17] = \A[15] ;
  assign \A[15]  = A[15];
  assign E[17] = \C[20] ;
  assign E[22] = \C[20] ;
  assign E[25] = \C[20] ;
  assign E[18] = \C[20] ;
  assign E[19] = \C[20] ;
  assign C[27] = \C[20] ;
  assign E[21] = \C[20] ;
  assign E[23] = \C[20] ;
  assign E[24] = \C[20] ;
  assign E[20] = \C[20] ;
  assign E[26] = \C[20] ;
  assign E[27] = \C[20] ;
  assign E[28] = \C[20] ;
  assign E[29] = \C[20] ;
  assign E[30] = \C[20] ;
  assign E[31] = \C[20] ;
  assign C[16] = \C[20] ;
  assign C[31] = \C[20] ;
  assign C[17] = \C[20] ;
  assign C[18] = \C[20] ;
  assign C[19] = \C[20] ;
  assign C[22] = \C[20] ;
  assign C[21] = \C[20] ;
  assign C[24] = \C[20] ;
  assign C[23] = \C[20] ;
  assign C[26] = \C[20] ;
  assign C[25] = \C[20] ;
  assign C[28] = \C[20] ;
  assign C[30] = \C[20] ;
  assign C[29] = \C[20] ;
  assign C[20] = \C[20] ;
  assign B[2] = \D[3] ;
  assign D[3] = \D[3] ;
  assign B[11] = \D[12] ;
  assign D[12] = \D[12] ;
  assign B[29] = \D[28] ;
  assign B[25] = \D[28] ;
  assign D[26] = \D[28] ;
  assign D[24] = \D[28] ;
  assign D[22] = \D[28] ;
  assign D[20] = \D[28] ;
  assign D[18] = \D[28] ;
  assign D[16] = \D[28] ;
  assign B[30] = \D[28] ;
  assign B[28] = \D[28] ;
  assign B[26] = \D[28] ;
  assign B[24] = \D[28] ;
  assign B[23] = \D[28] ;
  assign B[22] = \D[28] ;
  assign B[21] = \D[28] ;
  assign B[20] = \D[28] ;
  assign B[19] = \D[28] ;
  assign B[18] = \D[28] ;
  assign B[17] = \D[28] ;
  assign B[16] = \D[28] ;
  assign B[15] = \D[28] ;
  assign D[31] = \D[28] ;
  assign D[30] = \D[28] ;
  assign D[29] = \D[28] ;
  assign D[28] = \D[28] ;

  XOR2_X1 U29 ( .A(n8), .B(\A[7] ), .Z(E[8]) );
  XOR2_X1 U30 ( .A(n9), .B(\A[6] ), .Z(E[7]) );
  XOR2_X1 U31 ( .A(n12), .B(A[3]), .Z(\E[4] ) );
  XOR2_X1 U32 ( .A(\A[1] ), .B(\A[0] ), .Z(E[2]) );
  XOR2_X1 U34 ( .A(n16), .B(A[13]), .Z(E[14]) );
  XOR2_X1 U35 ( .A(n18), .B(\A[12] ), .Z(E[13]) );
  XOR2_X1 U36 ( .A(n21), .B(A[9]), .Z(E[10]) );
  BUF_X2 U2 ( .A(net25272), .Z(\C[20] ) );
  INV_X1 U3 ( .A(n6), .ZN(net25272) );
  INV_X1 U4 ( .A(n108), .ZN(\D[28] ) );
  XNOR2_X1 U5 ( .A(n19), .B(\D[12] ), .ZN(E[12]) );
  XNOR2_X1 U6 ( .A(n10), .B(\A[5] ), .ZN(E[6]) );
  XNOR2_X1 U7 ( .A(n13), .B(\D[3] ), .ZN(E[3]) );
  OAI21_X1 U8 ( .B1(n14), .B2(n108), .A(n6), .ZN(E[16]) );
  NAND2_X1 U9 ( .A1(n10), .A2(n104), .ZN(n9) );
  NAND2_X1 U10 ( .A1(n19), .A2(n106), .ZN(n18) );
  NAND2_X1 U11 ( .A1(n108), .A2(n14), .ZN(n6) );
  NOR3_X1 U12 ( .A1(A[3]), .A2(A[4]), .A3(n12), .ZN(n10) );
  NOR3_X1 U13 ( .A1(A[10]), .A2(A[9]), .A3(n21), .ZN(n19) );
  XNOR2_X1 U14 ( .A(n99), .B(A[8]), .ZN(E[9]) );
  NOR2_X1 U15 ( .A1(n8), .A2(\A[7] ), .ZN(n99) );
  XNOR2_X1 U16 ( .A(n100), .B(A[14]), .ZN(E[15]) );
  NOR2_X1 U17 ( .A1(n16), .A2(A[13]), .ZN(n100) );
  NOR2_X1 U18 ( .A1(\A[1] ), .A2(\A[0] ), .ZN(n13) );
  XNOR2_X1 U19 ( .A(A[10]), .B(n22), .ZN(E[11]) );
  NOR2_X1 U20 ( .A1(A[9]), .A2(n21), .ZN(n22) );
  XNOR2_X1 U21 ( .A(A[4]), .B(n11), .ZN(E[5]) );
  NOR2_X1 U22 ( .A1(A[3]), .A2(n12), .ZN(n11) );
  NAND2_X1 U23 ( .A1(n13), .A2(n103), .ZN(n12) );
  OR3_X1 U24 ( .A1(\A[7] ), .A2(A[8]), .A3(n8), .ZN(n21) );
  OR3_X1 U25 ( .A1(A[13]), .A2(A[14]), .A3(n16), .ZN(n14) );
  OR2_X1 U26 ( .A1(n18), .A2(\A[12] ), .ZN(n16) );
  OR2_X1 U27 ( .A1(n9), .A2(\A[6] ), .ZN(n8) );
  INV_X1 U28 ( .A(n103), .ZN(\D[3] ) );
  INV_X1 U33 ( .A(A[2]), .ZN(n103) );
  INV_X1 U37 ( .A(\A[5] ), .ZN(n104) );
  INV_X1 U38 ( .A(n106), .ZN(\D[12] ) );
  INV_X1 U39 ( .A(A[11]), .ZN(n106) );
  INV_X1 U40 ( .A(\A[15] ), .ZN(n108) );
endmodule


module cla_adder_N32_0 ( A, B, Ci, Cout, Sum );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Ci;
  output Cout;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50;
  wire   [8:0] Carry;
  assign n3 = A[5];
  assign n4 = B[6];
  assign n5 = A[2];
  assign n6 = A[12];
  assign n7 = A[0];
  assign n8 = B[10];
  assign n9 = B[26];
  assign n10 = B[5];
  assign n11 = B[22];
  assign n12 = B[3];
  assign n13 = A[1];
  assign n14 = A[6];
  assign n15 = A[18];
  assign n16 = A[7];
  assign n17 = B[7];
  assign n18 = B[11];
  assign n19 = A[19];
  assign n20 = A[3];
  assign n21 = B[9];
  assign n22 = A[29];
  assign n23 = B[12];
  assign n24 = A[10];
  assign n25 = B[18];
  assign n26 = B[14];
  assign n27 = A[11];
  assign n28 = A[22];
  assign n29 = B[19];
  assign n30 = A[17];
  assign n31 = B[15];
  assign n32 = A[9];
  assign n33 = B[17];
  assign n34 = A[25];
  assign n35 = A[26];
  assign n36 = B[29];
  assign n37 = A[21];
  assign n38 = B[13];
  assign n39 = A[13];
  assign n40 = A[14];
  assign n41 = A[15];
  assign n42 = B[24];
  assign n43 = B[27];
  assign n44 = B[28];
  assign n45 = A[27];
  assign n46 = B[21];
  assign n47 = A[28];
  assign n48 = A[24];
  assign n49 = B[23];
  assign n50 = A[23];

  carry_generator_N32_Nblocks8_0 CG ( .A({A[31:30], n22, n47, n45, n35, n34, 
        n48, n50, n28, n37, A[20], n19, n15, n30, A[16], n41, n40, n39, n6, 
        n27, n24, n32, A[8], n16, n14, n3, A[4], n20, n5, n13, n7}), .B({
        B[31:30], n36, n44, n43, n9, B[25], n42, n49, n11, n46, B[20], n29, 
        n25, n33, B[16], n31, n26, n38, n23, n18, n8, n21, B[8], n17, n4, n10, 
        B[4], n12, B[2:0]}), .Ci(Ci), .Cout(Carry) );
  sum_generator_Nbits32_Nblocks8_0 SG ( .A({A[31:30], n22, n47, n45, n35, n34, 
        n48, n50, n28, n37, A[20], n19, n15, n30, A[16], n41, n40, n39, n6, 
        n27, n24, n32, A[8], n16, n14, n3, A[4], n20, n5, n13, n7}), .B({
        B[31:30], n36, n44, n43, n9, B[25], n42, n49, n11, n46, B[20], n29, 
        n25, n33, B[16], n31, n26, n38, n23, n18, n8, n21, B[8], n17, n4, n10, 
        B[4], n12, B[2:0]}), .Carry(Carry), .S(Sum), .Cout(Cout) );
endmodule


module generic_xor_N32 ( A, B, Y );
  input [31:0] A;
  output [31:0] Y;
  input B;
  wire   n1, n2, n3;

  xor_gate_0 X_gate_0 ( .A(A[0]), .B(n3), .Y(Y[0]) );
  xor_gate_31 X_gate_1 ( .A(A[1]), .B(n1), .Y(Y[1]) );
  xor_gate_30 X_gate_2 ( .A(A[2]), .B(n1), .Y(Y[2]) );
  xor_gate_29 X_gate_3 ( .A(A[3]), .B(n1), .Y(Y[3]) );
  xor_gate_28 X_gate_4 ( .A(A[4]), .B(n1), .Y(Y[4]) );
  xor_gate_27 X_gate_5 ( .A(A[5]), .B(n1), .Y(Y[5]) );
  xor_gate_26 X_gate_6 ( .A(A[6]), .B(n1), .Y(Y[6]) );
  xor_gate_25 X_gate_7 ( .A(A[7]), .B(n1), .Y(Y[7]) );
  xor_gate_24 X_gate_8 ( .A(A[8]), .B(n1), .Y(Y[8]) );
  xor_gate_23 X_gate_9 ( .A(A[9]), .B(n1), .Y(Y[9]) );
  xor_gate_22 X_gate_10 ( .A(A[10]), .B(n1), .Y(Y[10]) );
  xor_gate_21 X_gate_11 ( .A(A[11]), .B(n1), .Y(Y[11]) );
  xor_gate_20 X_gate_12 ( .A(A[12]), .B(n1), .Y(Y[12]) );
  xor_gate_19 X_gate_13 ( .A(A[13]), .B(n2), .Y(Y[13]) );
  xor_gate_18 X_gate_14 ( .A(A[14]), .B(n2), .Y(Y[14]) );
  xor_gate_17 X_gate_15 ( .A(A[15]), .B(n2), .Y(Y[15]) );
  xor_gate_16 X_gate_16 ( .A(A[16]), .B(n2), .Y(Y[16]) );
  xor_gate_15 X_gate_17 ( .A(A[17]), .B(n2), .Y(Y[17]) );
  xor_gate_14 X_gate_18 ( .A(A[18]), .B(n2), .Y(Y[18]) );
  xor_gate_13 X_gate_19 ( .A(A[19]), .B(n2), .Y(Y[19]) );
  xor_gate_12 X_gate_20 ( .A(A[20]), .B(n2), .Y(Y[20]) );
  xor_gate_11 X_gate_21 ( .A(A[21]), .B(n2), .Y(Y[21]) );
  xor_gate_10 X_gate_22 ( .A(A[22]), .B(n2), .Y(Y[22]) );
  xor_gate_9 X_gate_23 ( .A(A[23]), .B(n2), .Y(Y[23]) );
  xor_gate_8 X_gate_24 ( .A(A[24]), .B(n2), .Y(Y[24]) );
  xor_gate_7 X_gate_25 ( .A(A[25]), .B(n3), .Y(Y[25]) );
  xor_gate_6 X_gate_26 ( .A(A[26]), .B(n3), .Y(Y[26]) );
  xor_gate_5 X_gate_27 ( .A(A[27]), .B(n3), .Y(Y[27]) );
  xor_gate_4 X_gate_28 ( .A(A[28]), .B(n3), .Y(Y[28]) );
  xor_gate_3 X_gate_29 ( .A(A[29]), .B(n3), .Y(Y[29]) );
  xor_gate_2 X_gate_30 ( .A(A[30]), .B(n3), .Y(Y[30]) );
  xor_gate_1 X_gate_31 ( .A(A[31]), .B(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(B), .Z(n1) );
  BUF_X1 U2 ( .A(B), .Z(n2) );
  BUF_X1 U3 ( .A(B), .Z(n3) );
endmodule


module counter_DW01_dec_0 ( A, SUM );
  input [30:0] A;
  output [30:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n60, n61, n62,
         n63, n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;

  XOR2_X1 U48 ( .A(A[30]), .B(n34), .Z(SUM[30]) );
  OR2_X2 U3 ( .A1(n29), .A2(A[6]), .ZN(n1) );
  OR2_X1 U1 ( .A1(n6), .A2(A[4]), .ZN(n7) );
  OR2_X1 U2 ( .A1(n38), .A2(A[3]), .ZN(n6) );
  AND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(n69) );
  INV_X1 U5 ( .A(n12), .ZN(n57) );
  INV_X1 U6 ( .A(n50), .ZN(n51) );
  NAND2_X1 U7 ( .A1(n57), .A2(n15), .ZN(n14) );
  OR2_X1 U8 ( .A1(n77), .A2(n5), .ZN(n73) );
  AND2_X1 U9 ( .A1(n52), .A2(n53), .ZN(n50) );
  OAI21_X1 U10 ( .B1(n57), .B2(n15), .A(n14), .ZN(SUM[20]) );
  INV_X1 U11 ( .A(A[6]), .ZN(n26) );
  OAI21_X1 U12 ( .B1(n55), .B2(n56), .A(n54), .ZN(SUM[21]) );
  INV_X1 U13 ( .A(A[21]), .ZN(n56) );
  INV_X1 U14 ( .A(n14), .ZN(n55) );
  OAI21_X1 U15 ( .B1(n74), .B2(n75), .A(n73), .ZN(SUM[12]) );
  INV_X1 U16 ( .A(A[12]), .ZN(n75) );
  NOR2_X1 U17 ( .A1(n77), .A2(A[11]), .ZN(n74) );
  NOR2_X1 U18 ( .A1(n73), .A2(A[13]), .ZN(n71) );
  NOR2_X1 U19 ( .A1(n14), .A2(A[21]), .ZN(n52) );
  INV_X1 U20 ( .A(n76), .ZN(SUM[11]) );
  AOI21_X1 U21 ( .B1(n77), .B2(A[11]), .A(n74), .ZN(n76) );
  AND2_X1 U22 ( .A1(n79), .A2(n80), .ZN(n60) );
  NOR2_X1 U23 ( .A1(n10), .A2(A[16]), .ZN(n79) );
  NOR2_X1 U24 ( .A1(A[18]), .A2(A[17]), .ZN(n80) );
  NOR2_X1 U25 ( .A1(n42), .A2(A[27]), .ZN(n39) );
  NOR2_X1 U26 ( .A1(n1), .A2(A[7]), .ZN(n22) );
  NOR2_X1 U27 ( .A1(n87), .A2(A[17]), .ZN(n62) );
  OR2_X1 U28 ( .A1(n16), .A2(A[24]), .ZN(n81) );
  NOR2_X1 U29 ( .A1(A[29]), .A2(n35), .ZN(n34) );
  NOR2_X1 U30 ( .A1(A[14]), .A2(A[13]), .ZN(n3) );
  NOR2_X1 U31 ( .A1(n4), .A2(n5), .ZN(n2) );
  OR2_X1 U32 ( .A1(A[1]), .A2(A[0]), .ZN(n88) );
  INV_X1 U33 ( .A(n45), .ZN(SUM[25]) );
  INV_X1 U34 ( .A(n41), .ZN(SUM[27]) );
  INV_X1 U35 ( .A(A[20]), .ZN(n15) );
  NOR2_X1 U36 ( .A1(n82), .A2(n83), .ZN(n43) );
  NAND2_X1 U37 ( .A1(n50), .A2(n17), .ZN(n82) );
  OR2_X1 U38 ( .A1(A[25]), .A2(A[24]), .ZN(n83) );
  OAI21_X1 U39 ( .B1(n47), .B2(n48), .A(n81), .ZN(SUM[24]) );
  INV_X1 U40 ( .A(A[24]), .ZN(n48) );
  INV_X1 U41 ( .A(A[10]), .ZN(n78) );
  INV_X1 U42 ( .A(A[16]), .ZN(n68) );
  OR2_X1 U43 ( .A1(A[12]), .A2(A[11]), .ZN(n5) );
  INV_X1 U44 ( .A(A[17]), .ZN(n65) );
  OAI21_X1 U45 ( .B1(n71), .B2(n9), .A(n70), .ZN(SUM[14]) );
  INV_X1 U46 ( .A(A[14]), .ZN(n9) );
  INV_X1 U47 ( .A(n69), .ZN(n70) );
  INV_X1 U49 ( .A(A[8]), .ZN(n23) );
  INV_X1 U50 ( .A(n24), .ZN(SUM[7]) );
  INV_X1 U51 ( .A(n19), .ZN(SUM[9]) );
  INV_X1 U52 ( .A(n72), .ZN(SUM[13]) );
  AOI21_X1 U53 ( .B1(n73), .B2(A[13]), .A(n71), .ZN(n72) );
  INV_X1 U54 ( .A(A[18]), .ZN(n8) );
  INV_X1 U55 ( .A(A[22]), .ZN(n53) );
  INV_X1 U56 ( .A(A[19]), .ZN(n13) );
  INV_X1 U57 ( .A(A[15]), .ZN(n11) );
  INV_X1 U58 ( .A(A[1]), .ZN(n58) );
  INV_X1 U59 ( .A(A[3]), .ZN(n33) );
  INV_X1 U60 ( .A(A[5]), .ZN(n28) );
  INV_X1 U61 ( .A(n7), .ZN(n27) );
  INV_X1 U62 ( .A(A[2]), .ZN(n37) );
  INV_X1 U63 ( .A(n88), .ZN(n36) );
  OAI21_X1 U64 ( .B1(n30), .B2(n31), .A(n7), .ZN(SUM[4]) );
  INV_X1 U65 ( .A(A[4]), .ZN(n31) );
  INV_X1 U66 ( .A(n6), .ZN(n30) );
  INV_X1 U67 ( .A(A[23]), .ZN(n17) );
  INV_X1 U68 ( .A(A[28]), .ZN(n40) );
  INV_X1 U69 ( .A(A[26]), .ZN(n44) );
  OAI21_X1 U70 ( .B1(n39), .B2(n40), .A(n35), .ZN(SUM[28]) );
  OAI21_X1 U71 ( .B1(n60), .B2(n13), .A(n12), .ZN(SUM[19]) );
  INV_X1 U72 ( .A(n60), .ZN(n61) );
  AOI21_X1 U73 ( .B1(n42), .B2(A[27]), .A(n39), .ZN(n41) );
  NAND2_X1 U74 ( .A1(n39), .A2(n40), .ZN(n35) );
  OAI21_X1 U75 ( .B1(SUM[0]), .B2(n58), .A(n88), .ZN(SUM[1]) );
  OR2_X1 U76 ( .A1(n10), .A2(A[16]), .ZN(n87) );
  NOR2_X1 U77 ( .A1(n88), .A2(A[2]), .ZN(n32) );
  NOR2_X1 U78 ( .A1(n7), .A2(A[5]), .ZN(n25) );
  NAND2_X1 U79 ( .A1(n60), .A2(n13), .ZN(n12) );
  NOR2_X1 U80 ( .A1(n1), .A2(A[7]), .ZN(n84) );
  AND2_X2 U81 ( .A1(n84), .A2(n85), .ZN(n21) );
  AND2_X1 U82 ( .A1(n86), .A2(n23), .ZN(n85) );
  INV_X1 U83 ( .A(A[9]), .ZN(n86) );
  XNOR2_X1 U84 ( .A(A[29]), .B(n35), .ZN(SUM[29]) );
  NAND2_X1 U85 ( .A1(n69), .A2(n11), .ZN(n10) );
  OAI21_X1 U86 ( .B1(n69), .B2(n11), .A(n10), .ZN(SUM[15]) );
  OAI21_X1 U87 ( .B1(n43), .B2(n44), .A(n42), .ZN(SUM[26]) );
  OAI21_X1 U88 ( .B1(n32), .B2(n33), .A(n6), .ZN(SUM[3]) );
  INV_X1 U89 ( .A(n10), .ZN(n67) );
  AOI21_X1 U90 ( .B1(n81), .B2(A[25]), .A(n43), .ZN(n45) );
  NAND2_X1 U91 ( .A1(n43), .A2(n44), .ZN(n42) );
  INV_X1 U92 ( .A(n32), .ZN(n38) );
  NAND2_X1 U93 ( .A1(n50), .A2(n17), .ZN(n16) );
  OAI21_X1 U94 ( .B1(n25), .B2(n26), .A(n1), .ZN(SUM[6]) );
  OAI21_X1 U95 ( .B1(n67), .B2(n68), .A(n87), .ZN(SUM[16]) );
  OAI21_X1 U96 ( .B1(n50), .B2(n17), .A(n16), .ZN(SUM[23]) );
  OAI21_X1 U97 ( .B1(n27), .B2(n28), .A(n29), .ZN(SUM[5]) );
  INV_X1 U98 ( .A(n16), .ZN(n47) );
  INV_X1 U99 ( .A(n25), .ZN(n29) );
  OAI21_X1 U100 ( .B1(n36), .B2(n37), .A(n38), .ZN(SUM[2]) );
  OAI21_X1 U101 ( .B1(n79), .B2(n65), .A(n63), .ZN(SUM[17]) );
  INV_X1 U102 ( .A(A[0]), .ZN(SUM[0]) );
  OAI21_X1 U103 ( .B1(n22), .B2(n23), .A(n20), .ZN(SUM[8]) );
  OAI21_X1 U104 ( .B1(n62), .B2(n8), .A(n61), .ZN(SUM[18]) );
  INV_X1 U105 ( .A(n62), .ZN(n63) );
  OAI21_X1 U106 ( .B1(n52), .B2(n53), .A(n51), .ZN(SUM[22]) );
  AOI21_X1 U107 ( .B1(n20), .B2(A[9]), .A(n21), .ZN(n19) );
  AOI21_X1 U108 ( .B1(n1), .B2(A[7]), .A(n22), .ZN(n24) );
  OAI21_X1 U109 ( .B1(n21), .B2(n78), .A(n77), .ZN(SUM[10]) );
  INV_X1 U110 ( .A(n52), .ZN(n54) );
  NAND2_X1 U111 ( .A1(n21), .A2(n78), .ZN(n77) );
  NAND2_X1 U112 ( .A1(n21), .A2(n78), .ZN(n4) );
  NAND2_X1 U113 ( .A1(n22), .A2(n23), .ZN(n20) );
endmodule


module PC_incr_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U5 ( .A(A[28]), .B(n13), .Z(SUM[28]) );
  XOR2_X1 U6 ( .A(A[27]), .B(n14), .Z(SUM[27]) );
  XOR2_X1 U7 ( .A(A[26]), .B(n15), .Z(SUM[26]) );
  XOR2_X1 U8 ( .A(A[25]), .B(n16), .Z(SUM[25]) );
  XOR2_X1 U9 ( .A(A[24]), .B(n17), .Z(SUM[24]) );
  XOR2_X1 U10 ( .A(A[23]), .B(n18), .Z(SUM[23]) );
  XOR2_X1 U11 ( .A(A[21]), .B(n19), .Z(SUM[21]) );
  XOR2_X1 U12 ( .A(A[20]), .B(n21), .Z(SUM[20]) );
  XOR2_X1 U13 ( .A(A[19]), .B(n22), .Z(SUM[19]) );
  XOR2_X1 U14 ( .A(A[18]), .B(n23), .Z(SUM[18]) );
  XOR2_X1 U15 ( .A(A[29]), .B(n11), .Z(SUM[29]) );
  XOR2_X1 U16 ( .A(n10), .B(A[30]), .Z(SUM[30]) );
  XOR2_X1 U34 ( .A(A[7]), .B(n6), .Z(SUM[7]) );
  XOR2_X1 U35 ( .A(A[17]), .B(n24), .Z(SUM[17]) );
  XOR2_X1 U36 ( .A(A[13]), .B(n40), .Z(SUM[13]) );
  XOR2_X1 U37 ( .A(A[12]), .B(n43), .Z(SUM[12]) );
  XOR2_X1 U38 ( .A(n2), .B(A[16]), .Z(SUM[16]) );
  XOR2_X1 U39 ( .A(A[10]), .B(n46), .Z(SUM[10]) );
  XOR2_X1 U40 ( .A(A[9]), .B(n4), .Z(SUM[9]) );
  XOR2_X1 U41 ( .A(A[8]), .B(n5), .Z(SUM[8]) );
  XOR2_X1 U42 ( .A(A[5]), .B(n7), .Z(SUM[5]) );
  XOR2_X1 U43 ( .A(A[4]), .B(n33), .Z(SUM[4]) );
  INV_X1 U2 ( .A(n33), .ZN(n8) );
  INV_X1 U3 ( .A(n5), .ZN(n44) );
  XNOR2_X1 U4 ( .A(n41), .B(n38), .ZN(SUM[14]) );
  NOR2_X1 U17 ( .A1(n50), .A2(SUM[2]), .ZN(n33) );
  NOR2_X1 U18 ( .A1(n35), .A2(n39), .ZN(n38) );
  INV_X1 U19 ( .A(n40), .ZN(n39) );
  NOR2_X1 U20 ( .A1(n8), .A2(n34), .ZN(n5) );
  NOR2_X1 U21 ( .A1(n44), .A2(n31), .ZN(n43) );
  NOR2_X1 U22 ( .A1(n29), .A2(n42), .ZN(n40) );
  INV_X1 U23 ( .A(n43), .ZN(n42) );
  NOR2_X1 U24 ( .A1(n30), .A2(n31), .ZN(n27) );
  NAND2_X1 U25 ( .A1(n32), .A2(n33), .ZN(n30) );
  INV_X1 U26 ( .A(n34), .ZN(n32) );
  XOR2_X1 U27 ( .A(n51), .B(A[15]), .Z(SUM[15]) );
  AND2_X1 U28 ( .A1(n38), .A2(A[14]), .ZN(n51) );
  XNOR2_X1 U29 ( .A(n1), .B(A[6]), .ZN(SUM[6]) );
  XNOR2_X1 U30 ( .A(n45), .B(A[11]), .ZN(SUM[11]) );
  NAND2_X1 U31 ( .A1(n46), .A2(A[10]), .ZN(n45) );
  XNOR2_X1 U32 ( .A(n9), .B(A[31]), .ZN(SUM[31]) );
  NAND2_X1 U33 ( .A1(n10), .A2(A[30]), .ZN(n9) );
  XNOR2_X1 U44 ( .A(A[22]), .B(n3), .ZN(SUM[22]) );
  NAND4_X1 U45 ( .A1(A[7]), .A2(A[6]), .A3(A[5]), .A4(A[4]), .ZN(n34) );
  NAND4_X1 U46 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n31) );
  NOR2_X1 U47 ( .A1(n8), .A2(n48), .ZN(n7) );
  INV_X1 U48 ( .A(A[4]), .ZN(n48) );
  NOR2_X1 U49 ( .A1(n20), .A2(n3), .ZN(n18) );
  INV_X1 U50 ( .A(A[22]), .ZN(n20) );
  NOR2_X1 U51 ( .A1(n44), .A2(n47), .ZN(n4) );
  INV_X1 U52 ( .A(A[8]), .ZN(n47) );
  INV_X1 U53 ( .A(A[2]), .ZN(SUM[2]) );
  NAND2_X1 U54 ( .A1(A[21]), .A2(n19), .ZN(n3) );
  NAND2_X1 U55 ( .A1(A[5]), .A2(n7), .ZN(n1) );
  NOR2_X1 U56 ( .A1(n49), .A2(n1), .ZN(n6) );
  INV_X1 U57 ( .A(A[6]), .ZN(n49) );
  INV_X1 U58 ( .A(A[3]), .ZN(n50) );
  INV_X1 U59 ( .A(A[14]), .ZN(n41) );
  AND2_X1 U60 ( .A1(A[20]), .A2(n21), .ZN(n19) );
  AND2_X1 U61 ( .A1(n4), .A2(A[9]), .ZN(n46) );
  INV_X1 U62 ( .A(A[13]), .ZN(n35) );
  INV_X1 U63 ( .A(A[12]), .ZN(n29) );
  AND2_X1 U64 ( .A1(A[29]), .A2(n11), .ZN(n10) );
  AND2_X1 U65 ( .A1(A[23]), .A2(n18), .ZN(n17) );
  AND2_X1 U66 ( .A1(A[16]), .A2(n2), .ZN(n24) );
  AND2_X1 U67 ( .A1(A[17]), .A2(n24), .ZN(n23) );
  AND2_X1 U68 ( .A1(A[18]), .A2(n23), .ZN(n22) );
  AND2_X1 U69 ( .A1(A[19]), .A2(n22), .ZN(n21) );
  AND2_X1 U70 ( .A1(A[24]), .A2(n17), .ZN(n16) );
  AND2_X1 U71 ( .A1(A[25]), .A2(n16), .ZN(n15) );
  AND2_X1 U72 ( .A1(A[26]), .A2(n15), .ZN(n14) );
  AND2_X1 U73 ( .A1(A[27]), .A2(n14), .ZN(n13) );
  AND2_X1 U74 ( .A1(A[28]), .A2(n13), .ZN(n11) );
  AND2_X1 U75 ( .A1(n25), .A2(A[15]), .ZN(n2) );
  NOR2_X1 U76 ( .A1(n26), .A2(n41), .ZN(n25) );
  NAND2_X1 U77 ( .A1(n27), .A2(n28), .ZN(n26) );
  NOR2_X1 U78 ( .A1(n29), .A2(n35), .ZN(n28) );
  XNOR2_X1 U79 ( .A(A[2]), .B(n50), .ZN(SUM[3]) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_665 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_664 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA_X1 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(\carry[5] ), .B(A[5]), .Z(SUM[5]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module w_reg_file_M8_N8_F4_Nbit32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI;
  output CO;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U3 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule


module w_reg_file_M8_N8_F4_Nbit32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI;
  output CO;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U3 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule


module sum_generator_Nbits32_Nblocks8 ( A, B, Carry, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Carry;
  output [31:0] S;
  output Cout;

  assign Cout = Carry[8];

  carry_select_N4 CS_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Carry[0]), .S(S[3:0]) );
  carry_select_N4 CS_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Carry[1]), .S(S[7:4]) );
  carry_select_N4 CS_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Carry[2]), .S(S[11:8])
         );
  carry_select_N4 CS_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Carry[3]), .S(
        S[15:12]) );
  carry_select_N4 CS_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Carry[4]), .S(
        S[19:16]) );
  carry_select_N4 CS_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Carry[5]), .S(
        S[23:20]) );
  carry_select_N4 CS_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Carry[6]), .S(
        S[27:24]) );
  carry_select_N4 CS_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Carry[7]), .S(
        S[31:28]) );
endmodule


module carry_generator_N32_Nblocks8 ( A, B, Ci, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Ci;
  wire   g_cin, p_cin, \Gsignal[1][31] , \Gsignal[1][30] , \Gsignal[1][29] ,
         \Gsignal[1][28] , \Gsignal[1][27] , \Gsignal[1][26] ,
         \Gsignal[1][25] , \Gsignal[1][24] , \Gsignal[1][23] ,
         \Gsignal[1][22] , \Gsignal[1][21] , \Gsignal[1][20] ,
         \Gsignal[1][19] , \Gsignal[1][18] , \Gsignal[1][17] ,
         \Gsignal[1][16] , \Gsignal[1][15] , \Gsignal[1][14] ,
         \Gsignal[1][13] , \Gsignal[1][12] , \Gsignal[1][11] ,
         \Gsignal[1][10] , \Gsignal[1][9] , \Gsignal[1][8] , \Gsignal[1][7] ,
         \Gsignal[1][6] , \Gsignal[1][5] , \Gsignal[1][4] , \Gsignal[1][3] ,
         \Gsignal[1][2] , \Gsignal[1][1] , \Gsignal[1][0] , \Gsignal[2][31] ,
         \Gsignal[2][29] , \Gsignal[2][27] , \Gsignal[2][25] ,
         \Gsignal[2][23] , \Gsignal[2][21] , \Gsignal[2][19] ,
         \Gsignal[2][17] , \Gsignal[2][15] , \Gsignal[2][13] ,
         \Gsignal[2][11] , \Gsignal[2][9] , \Gsignal[2][7] , \Gsignal[2][5] ,
         \Gsignal[2][3] , \Gsignal[2][1] , \Gsignal[3][31] , \Gsignal[3][27] ,
         \Gsignal[3][23] , \Gsignal[3][19] , \Gsignal[3][15] ,
         \Gsignal[3][11] , \Gsignal[3][7] , \Gsignal[4][31] , \Gsignal[4][23] ,
         \Gsignal[4][15] , \Gsignal[5][31] , \Gsignal[5][27] ,
         \Psignal[1][31] , \Psignal[1][30] , \Psignal[1][29] ,
         \Psignal[1][28] , \Psignal[1][27] , \Psignal[1][26] ,
         \Psignal[1][25] , \Psignal[1][24] , \Psignal[1][23] ,
         \Psignal[1][22] , \Psignal[1][21] , \Psignal[1][20] ,
         \Psignal[1][19] , \Psignal[1][18] , \Psignal[1][17] ,
         \Psignal[1][16] , \Psignal[1][15] , \Psignal[1][14] ,
         \Psignal[1][13] , \Psignal[1][12] , \Psignal[1][11] ,
         \Psignal[1][10] , \Psignal[1][9] , \Psignal[1][8] , \Psignal[1][7] ,
         \Psignal[1][6] , \Psignal[1][5] , \Psignal[1][4] , \Psignal[1][3] ,
         \Psignal[1][2] , \Psignal[1][1] , \Psignal[2][31] , \Psignal[2][29] ,
         \Psignal[2][27] , \Psignal[2][25] , \Psignal[2][23] ,
         \Psignal[2][21] , \Psignal[2][19] , \Psignal[2][17] ,
         \Psignal[2][15] , \Psignal[2][13] , \Psignal[2][11] , \Psignal[2][9] ,
         \Psignal[2][7] , \Psignal[2][5] , \Psignal[2][3] , \Psignal[3][31] ,
         \Psignal[3][27] , \Psignal[3][23] , \Psignal[3][19] ,
         \Psignal[3][15] , \Psignal[3][11] , \Psignal[3][7] , \Psignal[4][31] ,
         \Psignal[4][23] , \Psignal[4][15] , \Psignal[5][31] ,
         \Psignal[5][27] ;
  assign Cout[0] = Ci;

  PGnet_block PGnet_Cin_0 ( .A(A[0]), .B(B[0]), .pout(p_cin), .gout(g_cin) );
  G GCin_0 ( .gleft(g_cin), .gright(Cout[0]), .pleft(p_cin), .gout(
        \Gsignal[1][0] ) );
  PGnet_block PGnet_1 ( .A(A[1]), .B(B[1]), .pout(\Psignal[1][1] ), .gout(
        \Gsignal[1][1] ) );
  PGnet_block PGnet_2 ( .A(A[2]), .B(B[2]), .pout(\Psignal[1][2] ), .gout(
        \Gsignal[1][2] ) );
  PGnet_block PGnet_3 ( .A(A[3]), .B(B[3]), .pout(\Psignal[1][3] ), .gout(
        \Gsignal[1][3] ) );
  PGnet_block PGnet_4 ( .A(A[4]), .B(B[4]), .pout(\Psignal[1][4] ), .gout(
        \Gsignal[1][4] ) );
  PGnet_block PGnet_5 ( .A(A[5]), .B(B[5]), .pout(\Psignal[1][5] ), .gout(
        \Gsignal[1][5] ) );
  PGnet_block PGnet_6 ( .A(A[6]), .B(B[6]), .pout(\Psignal[1][6] ), .gout(
        \Gsignal[1][6] ) );
  PGnet_block PGnet_7 ( .A(A[7]), .B(B[7]), .pout(\Psignal[1][7] ), .gout(
        \Gsignal[1][7] ) );
  PGnet_block PGnet_8 ( .A(A[8]), .B(B[8]), .pout(\Psignal[1][8] ), .gout(
        \Gsignal[1][8] ) );
  PGnet_block PGnet_9 ( .A(A[9]), .B(B[9]), .pout(\Psignal[1][9] ), .gout(
        \Gsignal[1][9] ) );
  PGnet_block PGnet_10 ( .A(A[10]), .B(B[10]), .pout(\Psignal[1][10] ), .gout(
        \Gsignal[1][10] ) );
  PGnet_block PGnet_11 ( .A(A[11]), .B(B[11]), .pout(\Psignal[1][11] ), .gout(
        \Gsignal[1][11] ) );
  PGnet_block PGnet_12 ( .A(A[12]), .B(B[12]), .pout(\Psignal[1][12] ), .gout(
        \Gsignal[1][12] ) );
  PGnet_block PGnet_13 ( .A(A[13]), .B(B[13]), .pout(\Psignal[1][13] ), .gout(
        \Gsignal[1][13] ) );
  PGnet_block PGnet_14 ( .A(A[14]), .B(B[14]), .pout(\Psignal[1][14] ), .gout(
        \Gsignal[1][14] ) );
  PGnet_block PGnet_15 ( .A(A[15]), .B(B[15]), .pout(\Psignal[1][15] ), .gout(
        \Gsignal[1][15] ) );
  PGnet_block PGnet_16 ( .A(A[16]), .B(B[16]), .pout(\Psignal[1][16] ), .gout(
        \Gsignal[1][16] ) );
  PGnet_block PGnet_17 ( .A(A[17]), .B(B[17]), .pout(\Psignal[1][17] ), .gout(
        \Gsignal[1][17] ) );
  PGnet_block PGnet_18 ( .A(A[18]), .B(B[18]), .pout(\Psignal[1][18] ), .gout(
        \Gsignal[1][18] ) );
  PGnet_block PGnet_19 ( .A(A[19]), .B(B[19]), .pout(\Psignal[1][19] ), .gout(
        \Gsignal[1][19] ) );
  PGnet_block PGnet_20 ( .A(A[20]), .B(B[20]), .pout(\Psignal[1][20] ), .gout(
        \Gsignal[1][20] ) );
  PGnet_block PGnet_21 ( .A(A[21]), .B(B[21]), .pout(\Psignal[1][21] ), .gout(
        \Gsignal[1][21] ) );
  PGnet_block PGnet_22 ( .A(A[22]), .B(B[22]), .pout(\Psignal[1][22] ), .gout(
        \Gsignal[1][22] ) );
  PGnet_block PGnet_23 ( .A(A[23]), .B(B[23]), .pout(\Psignal[1][23] ), .gout(
        \Gsignal[1][23] ) );
  PGnet_block PGnet_24 ( .A(A[24]), .B(B[24]), .pout(\Psignal[1][24] ), .gout(
        \Gsignal[1][24] ) );
  PGnet_block PGnet_25 ( .A(A[25]), .B(B[25]), .pout(\Psignal[1][25] ), .gout(
        \Gsignal[1][25] ) );
  PGnet_block PGnet_26 ( .A(A[26]), .B(B[26]), .pout(\Psignal[1][26] ), .gout(
        \Gsignal[1][26] ) );
  PGnet_block PGnet_27 ( .A(A[27]), .B(B[27]), .pout(\Psignal[1][27] ), .gout(
        \Gsignal[1][27] ) );
  PGnet_block PGnet_28 ( .A(A[28]), .B(B[28]), .pout(\Psignal[1][28] ), .gout(
        \Gsignal[1][28] ) );
  PGnet_block PGnet_29 ( .A(A[29]), .B(B[29]), .pout(\Psignal[1][29] ), .gout(
        \Gsignal[1][29] ) );
  PGnet_block PGnet_30 ( .A(A[30]), .B(B[30]), .pout(\Psignal[1][30] ), .gout(
        \Gsignal[1][30] ) );
  PGnet_block PGnet_31 ( .A(A[31]), .B(B[31]), .pout(\Psignal[1][31] ), .gout(
        \Gsignal[1][31] ) );
  G Gblock_1_1 ( .gleft(\Gsignal[1][1] ), .gright(\Gsignal[1][0] ), .pleft(
        \Psignal[1][1] ), .gout(\Gsignal[2][1] ) );
  PG PGblock_1_3 ( .gleft(\Gsignal[1][3] ), .gright(\Gsignal[1][2] ), .pleft(
        \Psignal[1][3] ), .pright(\Psignal[1][2] ), .pout(\Psignal[2][3] ), 
        .gout(\Gsignal[2][3] ) );
  PG PGblock_1_5 ( .gleft(\Gsignal[1][5] ), .gright(\Gsignal[1][4] ), .pleft(
        \Psignal[1][5] ), .pright(\Psignal[1][4] ), .pout(\Psignal[2][5] ), 
        .gout(\Gsignal[2][5] ) );
  PG PGblock_1_7 ( .gleft(\Gsignal[1][7] ), .gright(\Gsignal[1][6] ), .pleft(
        \Psignal[1][7] ), .pright(\Psignal[1][6] ), .pout(\Psignal[2][7] ), 
        .gout(\Gsignal[2][7] ) );
  PG PGblock_1_9 ( .gleft(\Gsignal[1][9] ), .gright(\Gsignal[1][8] ), .pleft(
        \Psignal[1][9] ), .pright(\Psignal[1][8] ), .pout(\Psignal[2][9] ), 
        .gout(\Gsignal[2][9] ) );
  PG PGblock_1_11 ( .gleft(\Gsignal[1][11] ), .gright(\Gsignal[1][10] ), 
        .pleft(\Psignal[1][11] ), .pright(\Psignal[1][10] ), .pout(
        \Psignal[2][11] ), .gout(\Gsignal[2][11] ) );
  PG PGblock_1_13 ( .gleft(\Gsignal[1][13] ), .gright(\Gsignal[1][12] ), 
        .pleft(\Psignal[1][13] ), .pright(\Psignal[1][12] ), .pout(
        \Psignal[2][13] ), .gout(\Gsignal[2][13] ) );
  PG PGblock_1_15 ( .gleft(\Gsignal[1][15] ), .gright(\Gsignal[1][14] ), 
        .pleft(\Psignal[1][15] ), .pright(\Psignal[1][14] ), .pout(
        \Psignal[2][15] ), .gout(\Gsignal[2][15] ) );
  PG PGblock_1_17 ( .gleft(\Gsignal[1][17] ), .gright(\Gsignal[1][16] ), 
        .pleft(\Psignal[1][17] ), .pright(\Psignal[1][16] ), .pout(
        \Psignal[2][17] ), .gout(\Gsignal[2][17] ) );
  PG PGblock_1_19 ( .gleft(\Gsignal[1][19] ), .gright(\Gsignal[1][18] ), 
        .pleft(\Psignal[1][19] ), .pright(\Psignal[1][18] ), .pout(
        \Psignal[2][19] ), .gout(\Gsignal[2][19] ) );
  PG PGblock_1_21 ( .gleft(\Gsignal[1][21] ), .gright(\Gsignal[1][20] ), 
        .pleft(\Psignal[1][21] ), .pright(\Psignal[1][20] ), .pout(
        \Psignal[2][21] ), .gout(\Gsignal[2][21] ) );
  PG PGblock_1_23 ( .gleft(\Gsignal[1][23] ), .gright(\Gsignal[1][22] ), 
        .pleft(\Psignal[1][23] ), .pright(\Psignal[1][22] ), .pout(
        \Psignal[2][23] ), .gout(\Gsignal[2][23] ) );
  PG PGblock_1_25 ( .gleft(\Gsignal[1][25] ), .gright(\Gsignal[1][24] ), 
        .pleft(\Psignal[1][25] ), .pright(\Psignal[1][24] ), .pout(
        \Psignal[2][25] ), .gout(\Gsignal[2][25] ) );
  PG PGblock_1_27 ( .gleft(\Gsignal[1][27] ), .gright(\Gsignal[1][26] ), 
        .pleft(\Psignal[1][27] ), .pright(\Psignal[1][26] ), .pout(
        \Psignal[2][27] ), .gout(\Gsignal[2][27] ) );
  PG PGblock_1_29 ( .gleft(\Gsignal[1][29] ), .gright(\Gsignal[1][28] ), 
        .pleft(\Psignal[1][29] ), .pright(\Psignal[1][28] ), .pout(
        \Psignal[2][29] ), .gout(\Gsignal[2][29] ) );
  PG PGblock_1_31 ( .gleft(\Gsignal[1][31] ), .gright(\Gsignal[1][30] ), 
        .pleft(\Psignal[1][31] ), .pright(\Psignal[1][30] ), .pout(
        \Psignal[2][31] ), .gout(\Gsignal[2][31] ) );
  G Gblock_2_3 ( .gleft(\Gsignal[2][3] ), .gright(\Gsignal[2][1] ), .pleft(
        \Psignal[2][3] ), .gout(Cout[1]) );
  PG PGblock_2_7 ( .gleft(\Gsignal[2][7] ), .gright(\Gsignal[2][5] ), .pleft(
        \Psignal[2][7] ), .pright(\Psignal[2][5] ), .pout(\Psignal[3][7] ), 
        .gout(\Gsignal[3][7] ) );
  PG PGblock_2_11 ( .gleft(\Gsignal[2][11] ), .gright(\Gsignal[2][9] ), 
        .pleft(\Psignal[2][11] ), .pright(\Psignal[2][9] ), .pout(
        \Psignal[3][11] ), .gout(\Gsignal[3][11] ) );
  PG PGblock_2_15 ( .gleft(\Gsignal[2][15] ), .gright(\Gsignal[2][13] ), 
        .pleft(\Psignal[2][15] ), .pright(\Psignal[2][13] ), .pout(
        \Psignal[3][15] ), .gout(\Gsignal[3][15] ) );
  PG PGblock_2_19 ( .gleft(\Gsignal[2][19] ), .gright(\Gsignal[2][17] ), 
        .pleft(\Psignal[2][19] ), .pright(\Psignal[2][17] ), .pout(
        \Psignal[3][19] ), .gout(\Gsignal[3][19] ) );
  PG PGblock_2_23 ( .gleft(\Gsignal[2][23] ), .gright(\Gsignal[2][21] ), 
        .pleft(\Psignal[2][23] ), .pright(\Psignal[2][21] ), .pout(
        \Psignal[3][23] ), .gout(\Gsignal[3][23] ) );
  PG PGblock_2_27 ( .gleft(\Gsignal[2][27] ), .gright(\Gsignal[2][25] ), 
        .pleft(\Psignal[2][27] ), .pright(\Psignal[2][25] ), .pout(
        \Psignal[3][27] ), .gout(\Gsignal[3][27] ) );
  PG PGblock_2_31 ( .gleft(\Gsignal[2][31] ), .gright(\Gsignal[2][29] ), 
        .pleft(\Psignal[2][31] ), .pright(\Psignal[2][29] ), .pout(
        \Psignal[3][31] ), .gout(\Gsignal[3][31] ) );
  G Gblock_3_7 ( .gleft(\Gsignal[3][7] ), .gright(Cout[1]), .pleft(
        \Psignal[3][7] ), .gout(Cout[2]) );
  PG PGblock_3_15 ( .gleft(\Gsignal[3][15] ), .gright(\Gsignal[3][11] ), 
        .pleft(\Psignal[3][15] ), .pright(\Psignal[3][11] ), .pout(
        \Psignal[4][15] ), .gout(\Gsignal[4][15] ) );
  PG PGblock_3_23 ( .gleft(\Gsignal[3][23] ), .gright(\Gsignal[3][19] ), 
        .pleft(\Psignal[3][23] ), .pright(\Psignal[3][19] ), .pout(
        \Psignal[4][23] ), .gout(\Gsignal[4][23] ) );
  PG PGblock_3_31 ( .gleft(\Gsignal[3][31] ), .gright(\Gsignal[3][27] ), 
        .pleft(\Psignal[3][31] ), .pright(\Psignal[3][27] ), .pout(
        \Psignal[4][31] ), .gout(\Gsignal[4][31] ) );
  G Gblock_4_11 ( .gleft(\Gsignal[3][11] ), .gright(Cout[2]), .pleft(
        \Psignal[3][11] ), .gout(Cout[3]) );
  G Gblock_4_15 ( .gleft(\Gsignal[4][15] ), .gright(Cout[2]), .pleft(
        \Psignal[4][15] ), .gout(Cout[4]) );
  PG PGblock_4_27 ( .gleft(\Gsignal[3][27] ), .gright(\Gsignal[4][23] ), 
        .pleft(\Psignal[3][27] ), .pright(\Psignal[4][23] ), .pout(
        \Psignal[5][27] ), .gout(\Gsignal[5][27] ) );
  PG PGblock_4_31 ( .gleft(\Gsignal[4][31] ), .gright(\Gsignal[4][23] ), 
        .pleft(\Psignal[4][31] ), .pright(\Psignal[4][23] ), .pout(
        \Psignal[5][31] ), .gout(\Gsignal[5][31] ) );
  G Gblock_5_19 ( .gleft(\Gsignal[3][19] ), .gright(Cout[4]), .pleft(
        \Psignal[3][19] ), .gout(Cout[5]) );
  G Gblock_5_23 ( .gleft(\Gsignal[4][23] ), .gright(Cout[4]), .pleft(
        \Psignal[4][23] ), .gout(Cout[6]) );
  G Gblock_5_27 ( .gleft(\Gsignal[5][27] ), .gright(Cout[4]), .pleft(
        \Psignal[5][27] ), .gout(Cout[7]) );
  G Gblock_5_31 ( .gleft(\Gsignal[5][31] ), .gright(Cout[4]), .pleft(
        \Psignal[5][31] ), .gout(Cout[8]) );
endmodule


module mux_alu ( addsub, mul, log, shift, lhi, gt, get, lt, let, eq, neq, 
    .sel({\sel[4] , \sel[3] , \sel[2] , \sel[1] , \sel[0] }), out_mux );
  input [31:0] addsub;
  input [31:0] mul;
  input [31:0] log;
  input [31:0] shift;
  input [31:0] lhi;
  output [31:0] out_mux;
  input gt, get, lt, let, eq, neq, \sel[4] , \sel[3] , \sel[2] , \sel[1] ,
         \sel[0] ;
  wire   n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n145, n146, n147, n148, n149, n150, n151, n152, n153, n2, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n144;
  tri   [31:0] out_mux;

  OAI33_X1 U128 ( .A1(n101), .A2(n30), .A3(n102), .B1(n103), .B2(sel[4]), .B3(
        sel[2]), .ZN(n16) );
  TBUF_X1 \out_mux_tri[0]  ( .A(n153), .EN(n119), .Z(out_mux[0]) );
  TBUF_X1 \out_mux_tri[1]  ( .A(n152), .EN(n119), .Z(out_mux[1]) );
  TBUF_X1 \out_mux_tri[2]  ( .A(n151), .EN(n119), .Z(out_mux[2]) );
  TBUF_X1 \out_mux_tri[3]  ( .A(n150), .EN(n119), .Z(out_mux[3]) );
  TBUF_X1 \out_mux_tri[4]  ( .A(n149), .EN(n119), .Z(out_mux[4]) );
  TBUF_X1 \out_mux_tri[5]  ( .A(n148), .EN(n119), .Z(out_mux[5]) );
  TBUF_X1 \out_mux_tri[6]  ( .A(n147), .EN(n119), .Z(out_mux[6]) );
  TBUF_X1 \out_mux_tri[7]  ( .A(n146), .EN(n119), .Z(out_mux[7]) );
  TBUF_X1 \out_mux_tri[8]  ( .A(n145), .EN(n119), .Z(out_mux[8]) );
  TBUF_X1 \out_mux_tri[9]  ( .A(n143), .EN(n119), .Z(out_mux[9]) );
  TBUF_X1 \out_mux_tri[10]  ( .A(n142), .EN(n119), .Z(out_mux[10]) );
  TBUF_X1 \out_mux_tri[11]  ( .A(n141), .EN(n119), .Z(out_mux[11]) );
  TBUF_X1 \out_mux_tri[12]  ( .A(n140), .EN(n120), .Z(out_mux[12]) );
  TBUF_X1 \out_mux_tri[13]  ( .A(n139), .EN(n120), .Z(out_mux[13]) );
  TBUF_X1 \out_mux_tri[14]  ( .A(n138), .EN(n120), .Z(out_mux[14]) );
  TBUF_X1 \out_mux_tri[15]  ( .A(n137), .EN(n120), .Z(out_mux[15]) );
  TBUF_X1 \out_mux_tri[16]  ( .A(n136), .EN(n120), .Z(out_mux[16]) );
  TBUF_X1 \out_mux_tri[17]  ( .A(n135), .EN(n120), .Z(out_mux[17]) );
  TBUF_X1 \out_mux_tri[18]  ( .A(n134), .EN(n120), .Z(out_mux[18]) );
  TBUF_X1 \out_mux_tri[19]  ( .A(n133), .EN(n120), .Z(out_mux[19]) );
  TBUF_X1 \out_mux_tri[20]  ( .A(n132), .EN(n120), .Z(out_mux[20]) );
  TBUF_X1 \out_mux_tri[21]  ( .A(n131), .EN(n120), .Z(out_mux[21]) );
  TBUF_X1 \out_mux_tri[22]  ( .A(n130), .EN(n120), .Z(out_mux[22]) );
  TBUF_X1 \out_mux_tri[23]  ( .A(n129), .EN(n120), .Z(out_mux[23]) );
  TBUF_X1 \out_mux_tri[24]  ( .A(n128), .EN(n144), .Z(out_mux[24]) );
  TBUF_X1 \out_mux_tri[25]  ( .A(n127), .EN(n144), .Z(out_mux[25]) );
  TBUF_X1 \out_mux_tri[26]  ( .A(n126), .EN(n144), .Z(out_mux[26]) );
  TBUF_X1 \out_mux_tri[27]  ( .A(n125), .EN(n144), .Z(out_mux[27]) );
  TBUF_X1 \out_mux_tri[28]  ( .A(n124), .EN(n144), .Z(out_mux[28]) );
  TBUF_X1 \out_mux_tri[29]  ( .A(n123), .EN(n144), .Z(out_mux[29]) );
  TBUF_X1 \out_mux_tri[30]  ( .A(n122), .EN(n144), .Z(out_mux[30]) );
  TBUF_X1 \out_mux_tri[31]  ( .A(n121), .EN(n144), .Z(out_mux[31]) );
  BUF_X1 U2 ( .A(n38), .Z(n104) );
  BUF_X1 U3 ( .A(n38), .Z(n105) );
  BUF_X1 U4 ( .A(n38), .Z(n106) );
  NOR3_X1 U5 ( .A1(n30), .A2(n25), .A3(n101), .ZN(n38) );
  BUF_X1 U6 ( .A(n17), .Z(n113) );
  BUF_X1 U7 ( .A(n17), .Z(n114) );
  BUF_X1 U8 ( .A(n37), .Z(n107) );
  BUF_X1 U9 ( .A(n37), .Z(n108) );
  BUF_X1 U10 ( .A(n16), .Z(n116) );
  BUF_X1 U11 ( .A(n16), .Z(n117) );
  BUF_X1 U12 ( .A(n36), .Z(n110) );
  BUF_X1 U13 ( .A(n36), .Z(n111) );
  BUF_X1 U14 ( .A(n16), .Z(n118) );
  BUF_X1 U15 ( .A(n36), .Z(n112) );
  AOI22_X1 U16 ( .A1(n24), .A2(gt), .B1(n25), .B2(let), .ZN(n23) );
  BUF_X1 U17 ( .A(n2), .Z(n120) );
  BUF_X1 U18 ( .A(n2), .Z(n119) );
  INV_X1 U19 ( .A(n102), .ZN(n25) );
  BUF_X1 U20 ( .A(n2), .Z(n144) );
  BUF_X1 U21 ( .A(n17), .Z(n115) );
  NAND2_X1 U22 ( .A1(n10), .A2(n12), .ZN(n101) );
  BUF_X1 U23 ( .A(n37), .Z(n109) );
  INV_X1 U24 ( .A(n24), .ZN(n13) );
  INV_X1 U25 ( .A(n35), .ZN(n29) );
  AOI22_X1 U26 ( .A1(get), .A2(n25), .B1(n26), .B2(gt), .ZN(n35) );
  NAND2_X1 U27 ( .A1(sel[3]), .A2(n28), .ZN(n103) );
  NOR4_X1 U28 ( .A1(n13), .A2(n12), .A3(n30), .A4(sel[3]), .ZN(n17) );
  NOR4_X1 U29 ( .A1(n101), .A2(n25), .A3(n24), .A4(sel[2]), .ZN(n36) );
  NAND2_X1 U30 ( .A1(n87), .A2(n88), .ZN(n127) );
  AOI22_X1 U31 ( .A1(log[25]), .A2(n104), .B1(addsub[25]), .B2(n110), .ZN(n87)
         );
  AOI222_X1 U32 ( .A1(mul[25]), .A2(n108), .B1(shift[25]), .B2(n116), .C1(
        lhi[25]), .C2(n114), .ZN(n88) );
  NAND2_X1 U33 ( .A1(n85), .A2(n86), .ZN(n128) );
  AOI22_X1 U34 ( .A1(log[24]), .A2(n104), .B1(addsub[24]), .B2(n110), .ZN(n85)
         );
  AOI222_X1 U35 ( .A1(mul[24]), .A2(n108), .B1(shift[24]), .B2(n116), .C1(
        lhi[24]), .C2(n114), .ZN(n86) );
  NAND2_X1 U36 ( .A1(n83), .A2(n84), .ZN(n129) );
  AOI22_X1 U37 ( .A1(log[23]), .A2(n104), .B1(addsub[23]), .B2(n110), .ZN(n83)
         );
  AOI222_X1 U38 ( .A1(mul[23]), .A2(n108), .B1(shift[23]), .B2(n116), .C1(
        lhi[23]), .C2(n114), .ZN(n84) );
  NAND2_X1 U39 ( .A1(n81), .A2(n82), .ZN(n130) );
  AOI22_X1 U40 ( .A1(log[22]), .A2(n104), .B1(addsub[22]), .B2(n110), .ZN(n81)
         );
  AOI222_X1 U41 ( .A1(mul[22]), .A2(n108), .B1(shift[22]), .B2(n116), .C1(
        lhi[22]), .C2(n114), .ZN(n82) );
  NAND2_X1 U42 ( .A1(n79), .A2(n80), .ZN(n131) );
  AOI22_X1 U43 ( .A1(log[21]), .A2(n104), .B1(addsub[21]), .B2(n110), .ZN(n79)
         );
  AOI222_X1 U44 ( .A1(mul[21]), .A2(n108), .B1(shift[21]), .B2(n116), .C1(
        lhi[21]), .C2(n114), .ZN(n80) );
  NAND2_X1 U45 ( .A1(n77), .A2(n78), .ZN(n132) );
  AOI22_X1 U46 ( .A1(log[20]), .A2(n104), .B1(addsub[20]), .B2(n110), .ZN(n77)
         );
  AOI222_X1 U47 ( .A1(mul[20]), .A2(n108), .B1(shift[20]), .B2(n116), .C1(
        lhi[20]), .C2(n114), .ZN(n78) );
  NAND2_X1 U48 ( .A1(n75), .A2(n76), .ZN(n133) );
  AOI22_X1 U49 ( .A1(log[19]), .A2(n105), .B1(addsub[19]), .B2(n111), .ZN(n75)
         );
  AOI222_X1 U50 ( .A1(mul[19]), .A2(n108), .B1(shift[19]), .B2(n117), .C1(
        lhi[19]), .C2(n114), .ZN(n76) );
  NAND2_X1 U51 ( .A1(n73), .A2(n74), .ZN(n134) );
  AOI22_X1 U52 ( .A1(log[18]), .A2(n105), .B1(addsub[18]), .B2(n111), .ZN(n73)
         );
  AOI222_X1 U53 ( .A1(mul[18]), .A2(n108), .B1(shift[18]), .B2(n117), .C1(
        lhi[18]), .C2(n114), .ZN(n74) );
  NAND2_X1 U54 ( .A1(n71), .A2(n72), .ZN(n135) );
  AOI22_X1 U55 ( .A1(log[17]), .A2(n105), .B1(addsub[17]), .B2(n111), .ZN(n71)
         );
  AOI222_X1 U56 ( .A1(mul[17]), .A2(n108), .B1(shift[17]), .B2(n117), .C1(
        lhi[17]), .C2(n114), .ZN(n72) );
  NAND2_X1 U57 ( .A1(n69), .A2(n70), .ZN(n136) );
  AOI22_X1 U58 ( .A1(log[16]), .A2(n105), .B1(addsub[16]), .B2(n111), .ZN(n69)
         );
  AOI222_X1 U59 ( .A1(mul[16]), .A2(n108), .B1(shift[16]), .B2(n117), .C1(
        lhi[16]), .C2(n114), .ZN(n70) );
  NAND2_X1 U60 ( .A1(n67), .A2(n68), .ZN(n137) );
  AOI22_X1 U61 ( .A1(log[15]), .A2(n105), .B1(addsub[15]), .B2(n111), .ZN(n67)
         );
  AOI222_X1 U62 ( .A1(mul[15]), .A2(n108), .B1(shift[15]), .B2(n117), .C1(
        lhi[15]), .C2(n114), .ZN(n68) );
  NAND2_X1 U63 ( .A1(n65), .A2(n66), .ZN(n138) );
  AOI22_X1 U64 ( .A1(log[14]), .A2(n105), .B1(addsub[14]), .B2(n111), .ZN(n65)
         );
  AOI222_X1 U65 ( .A1(mul[14]), .A2(n108), .B1(shift[14]), .B2(n117), .C1(
        lhi[14]), .C2(n114), .ZN(n66) );
  NAND2_X1 U66 ( .A1(n63), .A2(n64), .ZN(n139) );
  AOI22_X1 U67 ( .A1(log[13]), .A2(n105), .B1(addsub[13]), .B2(n111), .ZN(n63)
         );
  AOI222_X1 U68 ( .A1(mul[13]), .A2(n108), .B1(shift[13]), .B2(n117), .C1(
        lhi[13]), .C2(n114), .ZN(n64) );
  NOR3_X1 U69 ( .A1(n102), .A2(sel[2]), .A3(n101), .ZN(n37) );
  NOR2_X1 U70 ( .A1(sel[1]), .A2(sel[0]), .ZN(n24) );
  AOI21_X1 U71 ( .B1(n10), .B2(n11), .A(n12), .ZN(n2) );
  NAND2_X1 U72 ( .A1(sel[2]), .A2(n13), .ZN(n11) );
  NOR2_X1 U73 ( .A1(n28), .A2(sel[0]), .ZN(n26) );
  INV_X1 U74 ( .A(sel[2]), .ZN(n30) );
  AOI21_X1 U75 ( .B1(n26), .B2(lt), .A(n27), .ZN(n22) );
  AND3_X1 U76 ( .A1(get), .A2(n28), .A3(sel[0]), .ZN(n27) );
  AOI21_X1 U77 ( .B1(n32), .B2(n33), .A(n30), .ZN(n31) );
  AOI21_X1 U78 ( .B1(eq), .B2(n26), .A(n34), .ZN(n33) );
  AOI22_X1 U79 ( .A1(neq), .A2(n25), .B1(n24), .B2(lt), .ZN(n32) );
  AND3_X1 U80 ( .A1(let), .A2(n28), .A3(sel[0]), .ZN(n34) );
  INV_X1 U81 ( .A(sel[4]), .ZN(n12) );
  OAI21_X1 U82 ( .B1(n19), .B2(n10), .A(n20), .ZN(n18) );
  INV_X1 U83 ( .A(n21), .ZN(n20) );
  AOI21_X1 U84 ( .B1(n29), .B2(n30), .A(n31), .ZN(n19) );
  AOI211_X1 U85 ( .C1(n22), .C2(n23), .A(sel[2]), .B(n12), .ZN(n21) );
  NAND2_X1 U86 ( .A1(sel[1]), .A2(sel[0]), .ZN(n102) );
  INV_X1 U87 ( .A(sel[1]), .ZN(n28) );
  NAND2_X1 U88 ( .A1(n14), .A2(n15), .ZN(n153) );
  AOI222_X1 U89 ( .A1(addsub[0]), .A2(n112), .B1(mul[0]), .B2(n107), .C1(
        log[0]), .C2(n106), .ZN(n14) );
  AOI221_X1 U90 ( .B1(shift[0]), .B2(n118), .C1(lhi[0]), .C2(n113), .A(n18), 
        .ZN(n15) );
  INV_X1 U91 ( .A(sel[3]), .ZN(n10) );
  NAND2_X1 U92 ( .A1(n51), .A2(n52), .ZN(n146) );
  AOI22_X1 U93 ( .A1(log[7]), .A2(n106), .B1(addsub[7]), .B2(n112), .ZN(n51)
         );
  AOI222_X1 U94 ( .A1(mul[7]), .A2(n107), .B1(shift[7]), .B2(n118), .C1(lhi[7]), .C2(n113), .ZN(n52) );
  NAND2_X1 U95 ( .A1(n49), .A2(n50), .ZN(n147) );
  AOI22_X1 U96 ( .A1(log[6]), .A2(n106), .B1(addsub[6]), .B2(n112), .ZN(n49)
         );
  AOI222_X1 U97 ( .A1(mul[6]), .A2(n107), .B1(shift[6]), .B2(n118), .C1(lhi[6]), .C2(n113), .ZN(n50) );
  NAND2_X1 U98 ( .A1(n47), .A2(n48), .ZN(n148) );
  AOI22_X1 U99 ( .A1(log[5]), .A2(n106), .B1(addsub[5]), .B2(n112), .ZN(n47)
         );
  AOI222_X1 U100 ( .A1(mul[5]), .A2(n107), .B1(shift[5]), .B2(n118), .C1(
        lhi[5]), .C2(n113), .ZN(n48) );
  NAND2_X1 U101 ( .A1(n45), .A2(n46), .ZN(n149) );
  AOI22_X1 U102 ( .A1(log[4]), .A2(n106), .B1(addsub[4]), .B2(n112), .ZN(n45)
         );
  AOI222_X1 U103 ( .A1(mul[4]), .A2(n107), .B1(shift[4]), .B2(n118), .C1(
        lhi[4]), .C2(n113), .ZN(n46) );
  NAND2_X1 U104 ( .A1(n43), .A2(n44), .ZN(n150) );
  AOI22_X1 U105 ( .A1(log[3]), .A2(n106), .B1(addsub[3]), .B2(n112), .ZN(n43)
         );
  AOI222_X1 U106 ( .A1(mul[3]), .A2(n107), .B1(shift[3]), .B2(n118), .C1(
        lhi[3]), .C2(n113), .ZN(n44) );
  NAND2_X1 U107 ( .A1(n41), .A2(n42), .ZN(n151) );
  AOI22_X1 U108 ( .A1(log[2]), .A2(n106), .B1(addsub[2]), .B2(n112), .ZN(n41)
         );
  AOI222_X1 U109 ( .A1(mul[2]), .A2(n107), .B1(shift[2]), .B2(n118), .C1(
        lhi[2]), .C2(n113), .ZN(n42) );
  NAND2_X1 U110 ( .A1(n39), .A2(n40), .ZN(n152) );
  AOI22_X1 U111 ( .A1(log[1]), .A2(n106), .B1(addsub[1]), .B2(n112), .ZN(n39)
         );
  AOI222_X1 U112 ( .A1(mul[1]), .A2(n107), .B1(shift[1]), .B2(n118), .C1(
        lhi[1]), .C2(n113), .ZN(n40) );
  NAND2_X1 U113 ( .A1(n99), .A2(n100), .ZN(n121) );
  AOI22_X1 U114 ( .A1(log[31]), .A2(n104), .B1(addsub[31]), .B2(n110), .ZN(n99) );
  AOI222_X1 U115 ( .A1(mul[31]), .A2(n109), .B1(shift[31]), .B2(n116), .C1(
        lhi[31]), .C2(n115), .ZN(n100) );
  NAND2_X1 U116 ( .A1(n97), .A2(n98), .ZN(n122) );
  AOI22_X1 U117 ( .A1(log[30]), .A2(n104), .B1(addsub[30]), .B2(n110), .ZN(n97) );
  AOI222_X1 U118 ( .A1(mul[30]), .A2(n109), .B1(shift[30]), .B2(n116), .C1(
        lhi[30]), .C2(n115), .ZN(n98) );
  NAND2_X1 U119 ( .A1(n95), .A2(n96), .ZN(n123) );
  AOI22_X1 U120 ( .A1(log[29]), .A2(n104), .B1(addsub[29]), .B2(n110), .ZN(n95) );
  AOI222_X1 U121 ( .A1(mul[29]), .A2(n109), .B1(shift[29]), .B2(n116), .C1(
        lhi[29]), .C2(n115), .ZN(n96) );
  NAND2_X1 U122 ( .A1(n93), .A2(n94), .ZN(n124) );
  AOI22_X1 U123 ( .A1(log[28]), .A2(n104), .B1(addsub[28]), .B2(n110), .ZN(n93) );
  AOI222_X1 U124 ( .A1(mul[28]), .A2(n109), .B1(shift[28]), .B2(n116), .C1(
        lhi[28]), .C2(n115), .ZN(n94) );
  NAND2_X1 U125 ( .A1(n91), .A2(n92), .ZN(n125) );
  AOI22_X1 U126 ( .A1(log[27]), .A2(n104), .B1(addsub[27]), .B2(n110), .ZN(n91) );
  AOI222_X1 U127 ( .A1(mul[27]), .A2(n109), .B1(shift[27]), .B2(n116), .C1(
        lhi[27]), .C2(n115), .ZN(n92) );
  NAND2_X1 U129 ( .A1(n89), .A2(n90), .ZN(n126) );
  AOI22_X1 U130 ( .A1(log[26]), .A2(n104), .B1(addsub[26]), .B2(n110), .ZN(n89) );
  AOI222_X1 U131 ( .A1(mul[26]), .A2(n109), .B1(shift[26]), .B2(n116), .C1(
        lhi[26]), .C2(n115), .ZN(n90) );
  NAND2_X1 U132 ( .A1(n61), .A2(n62), .ZN(n140) );
  AOI22_X1 U133 ( .A1(log[12]), .A2(n105), .B1(addsub[12]), .B2(n111), .ZN(n61) );
  AOI222_X1 U134 ( .A1(mul[12]), .A2(n107), .B1(shift[12]), .B2(n117), .C1(
        lhi[12]), .C2(n113), .ZN(n62) );
  NAND2_X1 U135 ( .A1(n59), .A2(n60), .ZN(n141) );
  AOI22_X1 U136 ( .A1(log[11]), .A2(n105), .B1(addsub[11]), .B2(n111), .ZN(n59) );
  AOI222_X1 U137 ( .A1(mul[11]), .A2(n107), .B1(shift[11]), .B2(n117), .C1(
        lhi[11]), .C2(n113), .ZN(n60) );
  NAND2_X1 U138 ( .A1(n57), .A2(n58), .ZN(n142) );
  AOI22_X1 U139 ( .A1(log[10]), .A2(n105), .B1(addsub[10]), .B2(n111), .ZN(n57) );
  AOI222_X1 U140 ( .A1(mul[10]), .A2(n107), .B1(shift[10]), .B2(n117), .C1(
        lhi[10]), .C2(n113), .ZN(n58) );
  NAND2_X1 U141 ( .A1(n55), .A2(n56), .ZN(n143) );
  AOI22_X1 U142 ( .A1(log[9]), .A2(n105), .B1(addsub[9]), .B2(n111), .ZN(n55)
         );
  AOI222_X1 U143 ( .A1(mul[9]), .A2(n107), .B1(shift[9]), .B2(n117), .C1(
        lhi[9]), .C2(n113), .ZN(n56) );
  NAND2_X1 U144 ( .A1(n53), .A2(n54), .ZN(n145) );
  AOI22_X1 U145 ( .A1(log[8]), .A2(n105), .B1(addsub[8]), .B2(n111), .ZN(n53)
         );
  AOI222_X1 U146 ( .A1(mul[8]), .A2(n107), .B1(shift[8]), .B2(n117), .C1(
        lhi[8]), .C2(n113), .ZN(n54) );
endmodule


module comparator ( C, Sum, sign, gt, get, lt, let, eq, neq );
  input [31:0] Sum;
  input C, sign;
  output gt, get, lt, let, eq, neq;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  XOR2_X1 U16 ( .A(sign), .B(C), .Z(get) );
  INV_X1 U1 ( .A(gt), .ZN(let) );
  INV_X1 U2 ( .A(eq), .ZN(neq) );
  NOR4_X1 U3 ( .A1(Sum[23]), .A2(Sum[22]), .A3(Sum[21]), .A4(Sum[20]), .ZN(n9)
         );
  NOR4_X1 U4 ( .A1(Sum[9]), .A2(Sum[8]), .A3(Sum[7]), .A4(Sum[6]), .ZN(n13) );
  NOR4_X1 U5 ( .A1(Sum[16]), .A2(Sum[15]), .A3(Sum[14]), .A4(Sum[13]), .ZN(n7)
         );
  NOR2_X1 U6 ( .A1(lt), .A2(eq), .ZN(gt) );
  NOR2_X1 U7 ( .A1(n4), .A2(n5), .ZN(eq) );
  NAND4_X1 U8 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n4) );
  NAND4_X1 U9 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  NOR4_X1 U10 ( .A1(Sum[27]), .A2(Sum[26]), .A3(Sum[25]), .A4(Sum[24]), .ZN(
        n10) );
  NOR4_X1 U11 ( .A1(Sum[1]), .A2(Sum[19]), .A3(Sum[18]), .A4(Sum[17]), .ZN(n8)
         );
  NOR4_X1 U12 ( .A1(Sum[5]), .A2(Sum[4]), .A3(Sum[3]), .A4(Sum[31]), .ZN(n12)
         );
  NOR4_X1 U13 ( .A1(Sum[30]), .A2(Sum[2]), .A3(Sum[29]), .A4(Sum[28]), .ZN(n11) );
  NOR4_X1 U14 ( .A1(Sum[12]), .A2(Sum[11]), .A3(Sum[10]), .A4(Sum[0]), .ZN(n6)
         );
  INV_X1 U15 ( .A(get), .ZN(lt) );
endmodule


module shifter ( A, B, sel, C );
  input [31:0] A;
  input [31:0] B;
  input [1:0] sel;
  output [31:0] C;
  wire   n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [2:0] s3;
  wire   [38:0] m0;
  wire   [38:0] m8;
  wire   [38:0] m16;
  wire   [38:0] y;

  shift_firstLevel IL ( .A(A), .sel(sel), .mask00(m0), .mask08(m8), .mask16(
        m16) );
  shift_secondLevel IIL ( .sel(B[4:3]), .mask00(m0), .mask08(m8), .mask16(m16), 
        .Y(y) );
  shift_thirdLevel IIIL ( .sel(s3), .A(y), .Y(C) );
  AOI221_X1 U1 ( .B1(n6), .B2(n7), .C1(sel[0]), .C2(B[2]), .A(n8), .ZN(s3[2])
         );
  INV_X1 U2 ( .A(n6), .ZN(n11) );
  INV_X1 U3 ( .A(B[2]), .ZN(n7) );
  INV_X1 U4 ( .A(n9), .ZN(n8) );
  OAI21_X1 U5 ( .B1(B[2]), .B2(sel[0]), .A(sel[1]), .ZN(n9) );
  OAI22_X1 U6 ( .A1(B[0]), .A2(n10), .B1(n11), .B2(n13), .ZN(s3[0]) );
  INV_X1 U7 ( .A(B[0]), .ZN(n13) );
  OAI22_X1 U8 ( .A1(B[1]), .A2(n10), .B1(n11), .B2(n12), .ZN(s3[1]) );
  INV_X1 U9 ( .A(B[1]), .ZN(n12) );
  XNOR2_X1 U10 ( .A(sel[1]), .B(sel[0]), .ZN(n10) );
  NOR2_X1 U11 ( .A1(sel[0]), .A2(sel[1]), .ZN(n6) );
endmodule


module logical ( A, B, sel, Y );
  input [31:0] A;
  input [31:0] B;
  input [3:0] sel;
  output [31:0] Y;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201;

  OAI22_X1 U1 ( .A1(n121), .A2(n122), .B1(B[25]), .B2(n123), .ZN(Y[25]) );
  OAI22_X1 U2 ( .A1(n125), .A2(n126), .B1(B[24]), .B2(n127), .ZN(Y[24]) );
  OAI22_X1 U3 ( .A1(n129), .A2(n130), .B1(B[23]), .B2(n131), .ZN(Y[23]) );
  OAI22_X1 U4 ( .A1(n133), .A2(n134), .B1(B[22]), .B2(n135), .ZN(Y[22]) );
  OAI22_X1 U5 ( .A1(n137), .A2(n138), .B1(B[21]), .B2(n139), .ZN(Y[21]) );
  OAI22_X1 U6 ( .A1(n141), .A2(n142), .B1(B[20]), .B2(n143), .ZN(Y[20]) );
  OAI22_X1 U7 ( .A1(n149), .A2(n150), .B1(B[19]), .B2(n151), .ZN(Y[19]) );
  OAI22_X1 U8 ( .A1(n153), .A2(n154), .B1(B[18]), .B2(n155), .ZN(Y[18]) );
  OAI22_X1 U9 ( .A1(n157), .A2(n158), .B1(B[17]), .B2(n159), .ZN(Y[17]) );
  OAI22_X1 U10 ( .A1(n161), .A2(n162), .B1(B[16]), .B2(n163), .ZN(Y[16]) );
  OAI22_X1 U11 ( .A1(n165), .A2(n166), .B1(B[15]), .B2(n167), .ZN(Y[15]) );
  OAI22_X1 U12 ( .A1(n169), .A2(n170), .B1(B[14]), .B2(n171), .ZN(Y[14]) );
  OAI22_X1 U13 ( .A1(n173), .A2(n174), .B1(B[13]), .B2(n175), .ZN(Y[13]) );
  OAI22_X1 U14 ( .A1(n73), .A2(n74), .B1(B[7]), .B2(n75), .ZN(Y[7]) );
  OAI22_X1 U15 ( .A1(n77), .A2(n78), .B1(B[6]), .B2(n79), .ZN(Y[6]) );
  OAI22_X1 U16 ( .A1(n81), .A2(n82), .B1(B[5]), .B2(n83), .ZN(Y[5]) );
  OAI22_X1 U17 ( .A1(n85), .A2(n86), .B1(B[4]), .B2(n87), .ZN(Y[4]) );
  OAI22_X1 U18 ( .A1(n89), .A2(n90), .B1(B[3]), .B2(n91), .ZN(Y[3]) );
  OAI22_X1 U19 ( .A1(n101), .A2(n102), .B1(B[2]), .B2(n103), .ZN(Y[2]) );
  OAI22_X1 U20 ( .A1(n145), .A2(n146), .B1(B[1]), .B2(n147), .ZN(Y[1]) );
  OAI22_X1 U21 ( .A1(n93), .A2(n94), .B1(B[31]), .B2(n95), .ZN(Y[31]) );
  OAI22_X1 U22 ( .A1(n97), .A2(n98), .B1(B[30]), .B2(n99), .ZN(Y[30]) );
  OAI22_X1 U23 ( .A1(n105), .A2(n106), .B1(B[29]), .B2(n107), .ZN(Y[29]) );
  OAI22_X1 U24 ( .A1(n109), .A2(n110), .B1(B[28]), .B2(n111), .ZN(Y[28]) );
  OAI22_X1 U25 ( .A1(n113), .A2(n114), .B1(B[27]), .B2(n115), .ZN(Y[27]) );
  OAI22_X1 U26 ( .A1(n117), .A2(n118), .B1(B[26]), .B2(n119), .ZN(Y[26]) );
  OAI22_X1 U27 ( .A1(n177), .A2(n178), .B1(B[12]), .B2(n179), .ZN(Y[12]) );
  OAI22_X1 U28 ( .A1(n181), .A2(n182), .B1(B[11]), .B2(n183), .ZN(Y[11]) );
  OAI22_X1 U29 ( .A1(n185), .A2(n186), .B1(B[10]), .B2(n187), .ZN(Y[10]) );
  OAI22_X1 U30 ( .A1(n65), .A2(n66), .B1(B[9]), .B2(n67), .ZN(Y[9]) );
  OAI22_X1 U31 ( .A1(n69), .A2(n70), .B1(B[8]), .B2(n71), .ZN(Y[8]) );
  BUF_X1 U32 ( .A(sel[1]), .Z(n197) );
  BUF_X1 U33 ( .A(sel[0]), .Z(n194) );
  BUF_X1 U34 ( .A(sel[1]), .Z(n196) );
  BUF_X1 U35 ( .A(sel[0]), .Z(n193) );
  OAI22_X1 U36 ( .A1(n189), .A2(n190), .B1(B[0]), .B2(n191), .ZN(Y[0]) );
  INV_X1 U37 ( .A(B[0]), .ZN(n190) );
  AOI22_X1 U38 ( .A1(n199), .A2(n192), .B1(A[0]), .B2(n193), .ZN(n189) );
  AOI22_X1 U39 ( .A1(sel[3]), .A2(n192), .B1(A[0]), .B2(n196), .ZN(n191) );
  BUF_X1 U40 ( .A(sel[2]), .Z(n200) );
  BUF_X1 U41 ( .A(sel[2]), .Z(n199) );
  BUF_X1 U42 ( .A(sel[1]), .Z(n198) );
  BUF_X1 U43 ( .A(sel[0]), .Z(n195) );
  BUF_X1 U44 ( .A(sel[2]), .Z(n201) );
  AOI22_X1 U45 ( .A1(sel[3]), .A2(n96), .B1(A[31]), .B2(n198), .ZN(n95) );
  AOI22_X1 U46 ( .A1(sel[3]), .A2(n72), .B1(A[8]), .B2(n198), .ZN(n71) );
  AOI22_X1 U47 ( .A1(sel[3]), .A2(n76), .B1(A[7]), .B2(n198), .ZN(n75) );
  AOI22_X1 U48 ( .A1(sel[3]), .A2(n80), .B1(A[6]), .B2(n198), .ZN(n79) );
  AOI22_X1 U49 ( .A1(sel[3]), .A2(n84), .B1(A[5]), .B2(n198), .ZN(n83) );
  AOI22_X1 U50 ( .A1(sel[3]), .A2(n88), .B1(A[4]), .B2(n198), .ZN(n87) );
  AOI22_X1 U51 ( .A1(sel[3]), .A2(n92), .B1(A[3]), .B2(n198), .ZN(n91) );
  AOI22_X1 U52 ( .A1(sel[3]), .A2(n68), .B1(n198), .B2(A[9]), .ZN(n67) );
  AOI22_X1 U53 ( .A1(sel[3]), .A2(n100), .B1(A[30]), .B2(n197), .ZN(n99) );
  AOI22_X1 U54 ( .A1(sel[3]), .A2(n108), .B1(A[29]), .B2(n197), .ZN(n107) );
  AOI22_X1 U55 ( .A1(sel[3]), .A2(n112), .B1(A[28]), .B2(n197), .ZN(n111) );
  AOI22_X1 U56 ( .A1(sel[3]), .A2(n116), .B1(A[27]), .B2(n197), .ZN(n115) );
  AOI22_X1 U57 ( .A1(sel[3]), .A2(n120), .B1(A[26]), .B2(n197), .ZN(n119) );
  AOI22_X1 U58 ( .A1(sel[3]), .A2(n124), .B1(A[25]), .B2(n197), .ZN(n123) );
  AOI22_X1 U59 ( .A1(sel[3]), .A2(n128), .B1(A[24]), .B2(n197), .ZN(n127) );
  AOI22_X1 U60 ( .A1(sel[3]), .A2(n132), .B1(A[23]), .B2(n197), .ZN(n131) );
  AOI22_X1 U61 ( .A1(sel[3]), .A2(n136), .B1(A[22]), .B2(n197), .ZN(n135) );
  AOI22_X1 U62 ( .A1(sel[3]), .A2(n140), .B1(A[21]), .B2(n197), .ZN(n139) );
  AOI22_X1 U63 ( .A1(sel[3]), .A2(n144), .B1(A[20]), .B2(n197), .ZN(n143) );
  AOI22_X1 U64 ( .A1(sel[3]), .A2(n152), .B1(A[19]), .B2(n196), .ZN(n151) );
  AOI22_X1 U65 ( .A1(sel[3]), .A2(n156), .B1(A[18]), .B2(n196), .ZN(n155) );
  AOI22_X1 U66 ( .A1(sel[3]), .A2(n160), .B1(A[17]), .B2(n196), .ZN(n159) );
  AOI22_X1 U67 ( .A1(sel[3]), .A2(n164), .B1(A[16]), .B2(n196), .ZN(n163) );
  AOI22_X1 U68 ( .A1(sel[3]), .A2(n168), .B1(A[15]), .B2(n196), .ZN(n167) );
  AOI22_X1 U69 ( .A1(sel[3]), .A2(n172), .B1(A[14]), .B2(n196), .ZN(n171) );
  AOI22_X1 U70 ( .A1(sel[3]), .A2(n176), .B1(A[13]), .B2(n196), .ZN(n175) );
  AOI22_X1 U71 ( .A1(sel[3]), .A2(n180), .B1(A[12]), .B2(n196), .ZN(n179) );
  AOI22_X1 U72 ( .A1(sel[3]), .A2(n184), .B1(A[11]), .B2(n196), .ZN(n183) );
  AOI22_X1 U73 ( .A1(sel[3]), .A2(n188), .B1(A[10]), .B2(n196), .ZN(n187) );
  AOI22_X1 U74 ( .A1(sel[3]), .A2(n104), .B1(A[2]), .B2(n197), .ZN(n103) );
  AOI22_X1 U75 ( .A1(sel[3]), .A2(n148), .B1(A[1]), .B2(n196), .ZN(n147) );
  AOI22_X1 U76 ( .A1(n201), .A2(n96), .B1(A[31]), .B2(n195), .ZN(n93) );
  AOI22_X1 U77 ( .A1(n201), .A2(n72), .B1(A[8]), .B2(n195), .ZN(n69) );
  AOI22_X1 U78 ( .A1(n201), .A2(n76), .B1(A[7]), .B2(n195), .ZN(n73) );
  AOI22_X1 U79 ( .A1(n201), .A2(n80), .B1(A[6]), .B2(n195), .ZN(n77) );
  AOI22_X1 U80 ( .A1(n201), .A2(n84), .B1(A[5]), .B2(n195), .ZN(n81) );
  AOI22_X1 U81 ( .A1(n201), .A2(n88), .B1(A[4]), .B2(n195), .ZN(n85) );
  AOI22_X1 U82 ( .A1(n201), .A2(n92), .B1(A[3]), .B2(n195), .ZN(n89) );
  AOI22_X1 U83 ( .A1(n201), .A2(n68), .B1(n195), .B2(A[9]), .ZN(n65) );
  AOI22_X1 U84 ( .A1(n200), .A2(n100), .B1(A[30]), .B2(n194), .ZN(n97) );
  AOI22_X1 U85 ( .A1(n200), .A2(n108), .B1(A[29]), .B2(n194), .ZN(n105) );
  AOI22_X1 U86 ( .A1(n200), .A2(n112), .B1(A[28]), .B2(n194), .ZN(n109) );
  AOI22_X1 U87 ( .A1(n200), .A2(n116), .B1(A[27]), .B2(n194), .ZN(n113) );
  AOI22_X1 U88 ( .A1(n200), .A2(n120), .B1(A[26]), .B2(n194), .ZN(n117) );
  AOI22_X1 U89 ( .A1(n200), .A2(n124), .B1(A[25]), .B2(n194), .ZN(n121) );
  AOI22_X1 U90 ( .A1(n200), .A2(n128), .B1(A[24]), .B2(n194), .ZN(n125) );
  AOI22_X1 U91 ( .A1(n200), .A2(n132), .B1(A[23]), .B2(n194), .ZN(n129) );
  AOI22_X1 U92 ( .A1(n200), .A2(n136), .B1(A[22]), .B2(n194), .ZN(n133) );
  AOI22_X1 U93 ( .A1(n200), .A2(n140), .B1(A[21]), .B2(n194), .ZN(n137) );
  AOI22_X1 U94 ( .A1(n200), .A2(n144), .B1(A[20]), .B2(n194), .ZN(n141) );
  AOI22_X1 U95 ( .A1(n199), .A2(n152), .B1(A[19]), .B2(n193), .ZN(n149) );
  AOI22_X1 U96 ( .A1(n199), .A2(n156), .B1(A[18]), .B2(n193), .ZN(n153) );
  AOI22_X1 U97 ( .A1(n199), .A2(n160), .B1(A[17]), .B2(n193), .ZN(n157) );
  AOI22_X1 U98 ( .A1(n199), .A2(n164), .B1(A[16]), .B2(n193), .ZN(n161) );
  AOI22_X1 U99 ( .A1(n199), .A2(n168), .B1(A[15]), .B2(n193), .ZN(n165) );
  AOI22_X1 U100 ( .A1(n199), .A2(n172), .B1(A[14]), .B2(n193), .ZN(n169) );
  AOI22_X1 U101 ( .A1(n199), .A2(n176), .B1(A[13]), .B2(n193), .ZN(n173) );
  AOI22_X1 U102 ( .A1(n199), .A2(n180), .B1(A[12]), .B2(n193), .ZN(n177) );
  AOI22_X1 U103 ( .A1(n199), .A2(n184), .B1(A[11]), .B2(n193), .ZN(n181) );
  AOI22_X1 U104 ( .A1(n199), .A2(n188), .B1(A[10]), .B2(n193), .ZN(n185) );
  AOI22_X1 U105 ( .A1(n200), .A2(n104), .B1(A[2]), .B2(n194), .ZN(n101) );
  AOI22_X1 U106 ( .A1(n199), .A2(n148), .B1(A[1]), .B2(n193), .ZN(n145) );
  INV_X1 U107 ( .A(A[9]), .ZN(n68) );
  INV_X1 U108 ( .A(A[31]), .ZN(n96) );
  INV_X1 U109 ( .A(A[30]), .ZN(n100) );
  INV_X1 U110 ( .A(A[29]), .ZN(n108) );
  INV_X1 U111 ( .A(A[28]), .ZN(n112) );
  INV_X1 U112 ( .A(A[27]), .ZN(n116) );
  INV_X1 U113 ( .A(A[26]), .ZN(n120) );
  INV_X1 U114 ( .A(A[25]), .ZN(n124) );
  INV_X1 U115 ( .A(A[24]), .ZN(n128) );
  INV_X1 U116 ( .A(A[23]), .ZN(n132) );
  INV_X1 U117 ( .A(A[22]), .ZN(n136) );
  INV_X1 U118 ( .A(A[21]), .ZN(n140) );
  INV_X1 U119 ( .A(A[20]), .ZN(n144) );
  INV_X1 U120 ( .A(A[19]), .ZN(n152) );
  INV_X1 U121 ( .A(A[18]), .ZN(n156) );
  INV_X1 U122 ( .A(A[17]), .ZN(n160) );
  INV_X1 U123 ( .A(A[16]), .ZN(n164) );
  INV_X1 U124 ( .A(A[15]), .ZN(n168) );
  INV_X1 U125 ( .A(A[14]), .ZN(n172) );
  INV_X1 U126 ( .A(A[13]), .ZN(n176) );
  INV_X1 U127 ( .A(A[12]), .ZN(n180) );
  INV_X1 U128 ( .A(A[11]), .ZN(n184) );
  INV_X1 U129 ( .A(A[10]), .ZN(n188) );
  INV_X1 U130 ( .A(A[8]), .ZN(n72) );
  INV_X1 U131 ( .A(A[7]), .ZN(n76) );
  INV_X1 U132 ( .A(A[6]), .ZN(n80) );
  INV_X1 U133 ( .A(A[5]), .ZN(n84) );
  INV_X1 U134 ( .A(A[4]), .ZN(n88) );
  INV_X1 U135 ( .A(A[3]), .ZN(n92) );
  INV_X1 U136 ( .A(A[2]), .ZN(n104) );
  INV_X1 U137 ( .A(A[1]), .ZN(n148) );
  INV_X1 U138 ( .A(A[0]), .ZN(n192) );
  INV_X1 U139 ( .A(B[31]), .ZN(n94) );
  INV_X1 U140 ( .A(B[30]), .ZN(n98) );
  INV_X1 U141 ( .A(B[29]), .ZN(n106) );
  INV_X1 U142 ( .A(B[28]), .ZN(n110) );
  INV_X1 U143 ( .A(B[27]), .ZN(n114) );
  INV_X1 U144 ( .A(B[26]), .ZN(n118) );
  INV_X1 U145 ( .A(B[25]), .ZN(n122) );
  INV_X1 U146 ( .A(B[24]), .ZN(n126) );
  INV_X1 U147 ( .A(B[23]), .ZN(n130) );
  INV_X1 U148 ( .A(B[22]), .ZN(n134) );
  INV_X1 U149 ( .A(B[21]), .ZN(n138) );
  INV_X1 U150 ( .A(B[20]), .ZN(n142) );
  INV_X1 U151 ( .A(B[19]), .ZN(n150) );
  INV_X1 U152 ( .A(B[18]), .ZN(n154) );
  INV_X1 U153 ( .A(B[17]), .ZN(n158) );
  INV_X1 U154 ( .A(B[16]), .ZN(n162) );
  INV_X1 U155 ( .A(B[15]), .ZN(n166) );
  INV_X1 U156 ( .A(B[14]), .ZN(n170) );
  INV_X1 U157 ( .A(B[13]), .ZN(n174) );
  INV_X1 U158 ( .A(B[12]), .ZN(n178) );
  INV_X1 U159 ( .A(B[11]), .ZN(n182) );
  INV_X1 U160 ( .A(B[10]), .ZN(n186) );
  INV_X1 U161 ( .A(B[9]), .ZN(n66) );
  INV_X1 U162 ( .A(B[8]), .ZN(n70) );
  INV_X1 U163 ( .A(B[7]), .ZN(n74) );
  INV_X1 U164 ( .A(B[6]), .ZN(n78) );
  INV_X1 U165 ( .A(B[5]), .ZN(n82) );
  INV_X1 U166 ( .A(B[4]), .ZN(n86) );
  INV_X1 U167 ( .A(B[3]), .ZN(n90) );
  INV_X1 U168 ( .A(B[2]), .ZN(n102) );
  INV_X1 U169 ( .A(B[1]), .ZN(n146) );
endmodule


module booth_mul_N16 ( A, B, Y );
  input [15:0] A;
  input [15:0] B;
  output [31:0] Y;
  wire   \muxInE[7][31] , \muxInE[7][30] , \muxInE[7][29] , \muxInE[7][28] ,
         \muxInE[7][27] , \muxInE[7][26] , \muxInE[7][25] , \muxInE[7][24] ,
         \muxInE[7][23] , \muxInE[7][22] , \muxInE[7][21] , \muxInE[7][20] ,
         \muxInE[7][19] , \muxInE[7][18] , \muxInE[7][17] , \muxInE[7][16] ,
         \muxInE[7][15] , \muxInE[6][31] , \muxInE[6][30] , \muxInE[6][29] ,
         \muxInE[6][28] , \muxInE[6][27] , \muxInE[6][26] , \muxInE[6][25] ,
         \muxInE[6][24] , \muxInE[6][23] , \muxInE[6][22] , \muxInE[6][21] ,
         \muxInE[6][20] , \muxInE[6][19] , \muxInE[6][18] , \muxInE[6][17] ,
         \muxInE[6][16] , \muxInE[6][15] , \muxInE[6][14] , \muxInE[6][13] ,
         \muxInE[5][31] , \muxInE[5][30] , \muxInE[5][29] , \muxInE[5][28] ,
         \muxInE[5][27] , \muxInE[5][26] , \muxInE[5][25] , \muxInE[5][24] ,
         \muxInE[5][23] , \muxInE[5][22] , \muxInE[5][21] , \muxInE[5][20] ,
         \muxInE[5][19] , \muxInE[5][18] , \muxInE[5][17] , \muxInE[5][16] ,
         \muxInE[5][15] , \muxInE[5][14] , \muxInE[5][13] , \muxInE[5][12] ,
         \muxInE[5][11] , \muxInE[4][31] , \muxInE[4][30] , \muxInE[4][29] ,
         \muxInE[4][28] , \muxInE[4][27] , \muxInE[4][26] , \muxInE[4][25] ,
         \muxInE[4][24] , \muxInE[4][23] , \muxInE[4][22] , \muxInE[4][21] ,
         \muxInE[4][20] , \muxInE[4][19] , \muxInE[4][18] , \muxInE[4][17] ,
         \muxInE[4][16] , \muxInE[4][15] , \muxInE[4][14] , \muxInE[4][13] ,
         \muxInE[4][12] , \muxInE[4][11] , \muxInE[4][10] , \muxInE[4][9] ,
         \muxInE[3][31] , \muxInE[3][30] , \muxInE[3][29] , \muxInE[3][28] ,
         \muxInE[3][27] , \muxInE[3][26] , \muxInE[3][25] , \muxInE[3][24] ,
         \muxInE[3][23] , \muxInE[3][22] , \muxInE[3][21] , \muxInE[3][20] ,
         \muxInE[3][19] , \muxInE[3][18] , \muxInE[3][17] , \muxInE[3][16] ,
         \muxInE[3][15] , \muxInE[3][14] , \muxInE[3][13] , \muxInE[3][12] ,
         \muxInE[3][11] , \muxInE[3][10] , \muxInE[3][9] , \muxInE[3][8] ,
         \muxInE[3][7] , \muxInE[2][31] , \muxInE[2][30] , \muxInE[2][29] ,
         \muxInE[2][28] , \muxInE[2][27] , \muxInE[2][26] , \muxInE[2][25] ,
         \muxInE[2][24] , \muxInE[2][23] , \muxInE[2][22] , \muxInE[2][21] ,
         \muxInE[2][19] , \muxInE[2][18] , \muxInE[2][17] , \muxInE[2][16] ,
         \muxInE[2][15] , \muxInE[2][14] , \muxInE[2][13] , \muxInE[2][12] ,
         \muxInE[2][11] , \muxInE[2][10] , \muxInE[2][9] , \muxInE[2][8] ,
         \muxInE[2][7] , \muxInE[2][6] , \muxInE[2][5] , \muxInE[1][31] ,
         \muxInE[1][30] , \muxInE[1][29] , \muxInE[1][28] , \muxInE[1][27] ,
         \muxInE[1][26] , \muxInE[1][25] , \muxInE[1][24] , \muxInE[1][23] ,
         \muxInE[1][22] , \muxInE[1][21] , \muxInE[1][20] , \muxInE[1][19] ,
         \muxInE[1][18] , \muxInE[1][17] , \muxInE[1][16] , \muxInE[1][15] ,
         \muxInE[1][14] , \muxInE[1][13] , \muxInE[1][12] , \muxInE[1][11] ,
         \muxInE[1][10] , \muxInE[1][9] , \muxInE[1][8] , \muxInE[1][7] ,
         \muxInE[1][6] , \muxInE[1][5] , \muxInE[1][4] , \muxInE[1][3] ,
         \muxInE[0][31] , \muxInE[0][30] , \muxInE[0][29] , \muxInE[0][28] ,
         \muxInE[0][27] , \muxInE[0][26] , \muxInE[0][24] , \muxInE[0][23] ,
         \muxInE[0][21] , \muxInE[0][20] , \muxInE[0][19] , \muxInE[0][18] ,
         \muxInE[0][16] , \muxInE[0][15] , \muxInE[0][14] , \muxInE[0][13] ,
         \muxInE[0][12] , \muxInE[0][11] , \muxInE[0][10] , \muxInE[0][9] ,
         \muxInE[0][8] , \muxInE[0][7] , \muxInE[0][6] , \muxInE[0][5] ,
         \muxInE[0][4] , \muxInE[0][3] , \muxInE[0][2] , \muxInE[0][1] ,
         \muxInD[7][31] , \muxInD[7][30] , \muxInD[7][29] , \muxInD[7][28] ,
         \muxInD[7][27] , \muxInD[7][26] , \muxInD[7][25] , \muxInD[7][24] ,
         \muxInD[7][23] , \muxInD[7][22] , \muxInD[7][21] , \muxInD[7][20] ,
         \muxInD[7][19] , \muxInD[7][18] , \muxInD[7][17] , \muxInD[7][16] ,
         \muxInD[7][15] , \muxInD[6][31] , \muxInD[6][30] , \muxInD[6][29] ,
         \muxInD[6][28] , \muxInD[6][27] , \muxInD[6][26] , \muxInD[6][25] ,
         \muxInD[6][24] , \muxInD[6][23] , \muxInD[6][22] , \muxInD[6][21] ,
         \muxInD[6][20] , \muxInD[6][19] , \muxInD[6][18] , \muxInD[6][17] ,
         \muxInD[6][16] , \muxInD[6][15] , \muxInD[6][14] , \muxInD[6][13] ,
         \muxInD[5][31] , \muxInD[5][30] , \muxInD[5][29] , \muxInD[5][28] ,
         \muxInD[5][27] , \muxInD[5][26] , \muxInD[5][25] , \muxInD[5][24] ,
         \muxInD[5][23] , \muxInD[5][22] , \muxInD[5][21] , \muxInD[5][20] ,
         \muxInD[5][19] , \muxInD[5][18] , \muxInD[5][17] , \muxInD[5][16] ,
         \muxInD[5][15] , \muxInD[5][14] , \muxInD[5][13] , \muxInD[5][12] ,
         \muxInD[5][11] , \muxInD[4][31] , \muxInD[4][30] , \muxInD[4][29] ,
         \muxInD[4][28] , \muxInD[4][27] , \muxInD[4][26] , \muxInD[4][25] ,
         \muxInD[4][24] , \muxInD[4][23] , \muxInD[4][22] , \muxInD[4][21] ,
         \muxInD[4][20] , \muxInD[4][19] , \muxInD[4][18] , \muxInD[4][17] ,
         \muxInD[4][16] , \muxInD[4][15] , \muxInD[4][14] , \muxInD[4][13] ,
         \muxInD[4][12] , \muxInD[4][11] , \muxInD[4][10] , \muxInD[4][9] ,
         \muxInD[3][31] , \muxInD[3][30] , \muxInD[3][29] , \muxInD[3][28] ,
         \muxInD[3][27] , \muxInD[3][26] , \muxInD[3][25] , \muxInD[3][24] ,
         \muxInD[3][23] , \muxInD[3][22] , \muxInD[3][21] , \muxInD[3][20] ,
         \muxInD[3][19] , \muxInD[3][18] , \muxInD[3][17] , \muxInD[3][16] ,
         \muxInD[3][15] , \muxInD[3][14] , \muxInD[3][13] , \muxInD[3][12] ,
         \muxInD[3][11] , \muxInD[3][10] , \muxInD[3][9] , \muxInD[3][8] ,
         \muxInD[3][7] , \muxInD[2][31] , \muxInD[2][30] , \muxInD[2][29] ,
         \muxInD[2][28] , \muxInD[2][27] , \muxInD[2][26] , \muxInD[2][25] ,
         \muxInD[2][24] , \muxInD[2][23] , \muxInD[2][22] , \muxInD[2][21] ,
         \muxInD[2][20] , \muxInD[2][19] , \muxInD[2][18] , \muxInD[2][17] ,
         \muxInD[2][16] , \muxInD[2][15] , \muxInD[2][14] , \muxInD[2][13] ,
         \muxInD[2][12] , \muxInD[2][11] , \muxInD[2][10] , \muxInD[2][9] ,
         \muxInD[2][8] , \muxInD[2][7] , \muxInD[2][6] , \muxInD[2][5] ,
         \muxInD[1][31] , \muxInD[1][30] , \muxInD[1][29] , \muxInD[1][28] ,
         \muxInD[1][27] , \muxInD[1][26] , \muxInD[1][25] , \muxInD[1][24] ,
         \muxInD[1][23] , \muxInD[1][22] , \muxInD[1][21] , \muxInD[1][20] ,
         \muxInD[1][19] , \muxInD[1][18] , \muxInD[1][17] , \muxInD[1][16] ,
         \muxInD[1][15] , \muxInD[1][14] , \muxInD[1][13] , \muxInD[1][12] ,
         \muxInD[1][11] , \muxInD[1][10] , \muxInD[1][9] , \muxInD[1][8] ,
         \muxInD[1][7] , \muxInD[1][6] , \muxInD[1][5] , \muxInD[1][4] ,
         \muxInD[1][3] , \muxInD[0][31] , \muxInD[0][30] , \muxInD[0][29] ,
         \muxInD[0][28] , \muxInD[0][27] , \muxInD[0][26] , \muxInD[0][25] ,
         \muxInD[0][24] , \muxInD[0][23] , \muxInD[0][22] , \muxInD[0][21] ,
         \muxInD[0][20] , \muxInD[0][19] , \muxInD[0][18] , \muxInD[0][17] ,
         \muxInD[0][16] , \muxInD[0][15] , \muxInD[0][14] , \muxInD[0][13] ,
         \muxInD[0][12] , \muxInD[0][11] , \muxInD[0][10] , \muxInD[0][9] ,
         \muxInD[0][8] , \muxInD[0][7] , \muxInD[0][6] , \muxInD[0][5] ,
         \muxInD[0][4] , \muxInD[0][3] , \muxInD[0][2] , \muxInD[0][1] ,
         \muxInC[7][31] , \muxInC[7][30] , \muxInC[7][29] , \muxInC[7][28] ,
         \muxInC[7][27] , \muxInC[7][26] , \muxInC[7][25] , \muxInC[7][24] ,
         \muxInC[7][23] , \muxInC[7][22] , \muxInC[7][21] , \muxInC[7][20] ,
         \muxInC[7][19] , \muxInC[7][18] , \muxInC[7][17] , \muxInC[7][16] ,
         \muxInC[7][15] , \muxInC[7][14] , \muxInC[6][31] , \muxInC[6][30] ,
         \muxInC[6][29] , \muxInC[6][28] , \muxInC[6][27] , \muxInC[6][26] ,
         \muxInC[6][25] , \muxInC[6][24] , \muxInC[6][23] , \muxInC[6][22] ,
         \muxInC[6][21] , \muxInC[6][20] , \muxInC[6][19] , \muxInC[6][18] ,
         \muxInC[6][17] , \muxInC[6][16] , \muxInC[6][15] , \muxInC[6][14] ,
         \muxInC[6][13] , \muxInC[6][12] , \muxInC[5][31] , \muxInC[5][30] ,
         \muxInC[5][29] , \muxInC[5][28] , \muxInC[5][27] , \muxInC[5][26] ,
         \muxInC[5][25] , \muxInC[5][24] , \muxInC[5][23] , \muxInC[5][22] ,
         \muxInC[5][21] , \muxInC[5][20] , \muxInC[5][19] , \muxInC[5][18] ,
         \muxInC[5][17] , \muxInC[5][16] , \muxInC[5][15] , \muxInC[5][14] ,
         \muxInC[5][13] , \muxInC[5][12] , \muxInC[5][11] , \muxInC[5][10] ,
         \muxInC[4][31] , \muxInC[4][30] , \muxInC[4][29] , \muxInC[4][28] ,
         \muxInC[4][27] , \muxInC[4][26] , \muxInC[4][25] , \muxInC[4][24] ,
         \muxInC[4][23] , \muxInC[4][22] , \muxInC[4][21] , \muxInC[4][20] ,
         \muxInC[4][19] , \muxInC[4][18] , \muxInC[4][17] , \muxInC[4][16] ,
         \muxInC[4][15] , \muxInC[4][14] , \muxInC[4][13] , \muxInC[4][12] ,
         \muxInC[4][11] , \muxInC[4][10] , \muxInC[4][9] , \muxInC[4][8] ,
         \muxInC[3][31] , \muxInC[3][30] , \muxInC[3][29] , \muxInC[3][28] ,
         \muxInC[3][27] , \muxInC[3][26] , \muxInC[3][25] , \muxInC[3][24] ,
         \muxInC[3][23] , \muxInC[3][22] , \muxInC[3][21] , \muxInC[3][20] ,
         \muxInC[3][19] , \muxInC[3][18] , \muxInC[3][17] , \muxInC[3][16] ,
         \muxInC[3][15] , \muxInC[3][14] , \muxInC[3][13] , \muxInC[3][12] ,
         \muxInC[3][11] , \muxInC[3][10] , \muxInC[3][9] , \muxInC[3][8] ,
         \muxInC[3][7] , \muxInC[3][6] , \muxInC[2][31] , \muxInC[2][30] ,
         \muxInC[2][29] , \muxInC[2][28] , \muxInC[2][27] , \muxInC[2][26] ,
         \muxInC[2][25] , \muxInC[2][24] , \muxInC[2][23] , \muxInC[2][22] ,
         \muxInC[2][21] , \muxInC[2][20] , \muxInC[2][19] , \muxInC[2][18] ,
         \muxInC[2][17] , \muxInC[2][16] , \muxInC[2][15] , \muxInC[2][14] ,
         \muxInC[2][13] , \muxInC[2][12] , \muxInC[2][11] , \muxInC[2][10] ,
         \muxInC[2][9] , \muxInC[2][8] , \muxInC[2][7] , \muxInC[2][6] ,
         \muxInC[2][5] , \muxInC[2][4] , \muxInC[1][31] , \muxInC[1][30] ,
         \muxInC[1][29] , \muxInC[1][28] , \muxInC[1][27] , \muxInC[1][26] ,
         \muxInC[1][25] , \muxInC[1][24] , \muxInC[1][23] , \muxInC[1][22] ,
         \muxInC[1][21] , \muxInC[1][20] , \muxInC[1][18] , \muxInC[1][17] ,
         \muxInC[1][16] , \muxInC[1][15] , \muxInC[1][14] , \muxInC[1][13] ,
         \muxInC[1][12] , \muxInC[1][11] , \muxInC[1][10] , \muxInC[1][9] ,
         \muxInC[1][8] , \muxInC[1][7] , \muxInC[1][6] , \muxInC[1][5] ,
         \muxInC[1][4] , \muxInC[1][3] , \muxInC[1][2] , \muxInC[0][31] ,
         \muxInC[0][30] , \muxInC[0][29] , \muxInC[0][28] , \muxInC[0][27] ,
         \muxInC[0][26] , \muxInC[0][25] , \muxInC[0][24] , \muxInC[0][23] ,
         \muxInC[0][22] , \muxInC[0][21] , \muxInC[0][20] , \muxInC[0][19] ,
         \muxInC[0][18] , \muxInC[0][17] , \muxInC[0][16] , \muxInC[0][15] ,
         \muxInC[0][14] , \muxInC[0][13] , \muxInC[0][12] , \muxInC[0][11] ,
         \muxInC[0][10] , \muxInC[0][9] , \muxInC[0][8] , \muxInC[0][7] ,
         \muxInC[0][6] , \muxInC[0][5] , \muxInC[0][4] , \muxInC[0][3] ,
         \muxInC[0][2] , \muxInC[0][1] , \muxInC[0][0] , \muxInB[7][31] ,
         \muxInB[7][30] , \muxInB[7][29] , \muxInB[7][28] , \muxInB[7][27] ,
         \muxInB[7][26] , \muxInB[7][25] , \muxInB[7][24] , \muxInB[7][23] ,
         \muxInB[7][22] , \muxInB[7][21] , \muxInB[7][20] , \muxInB[7][19] ,
         \muxInB[7][18] , \muxInB[7][17] , \muxInB[7][16] , \muxInB[7][15] ,
         \muxInB[7][14] , \muxInB[6][31] , \muxInB[6][30] , \muxInB[6][29] ,
         \muxInB[6][28] , \muxInB[6][27] , \muxInB[6][26] , \muxInB[6][25] ,
         \muxInB[6][24] , \muxInB[6][23] , \muxInB[6][22] , \muxInB[6][21] ,
         \muxInB[6][20] , \muxInB[6][19] , \muxInB[6][18] , \muxInB[6][17] ,
         \muxInB[6][16] , \muxInB[6][15] , \muxInB[6][14] , \muxInB[6][13] ,
         \muxInB[6][12] , \muxInB[5][31] , \muxInB[5][30] , \muxInB[5][29] ,
         \muxInB[5][28] , \muxInB[5][27] , \muxInB[5][26] , \muxInB[5][25] ,
         \muxInB[5][24] , \muxInB[5][23] , \muxInB[5][22] , \muxInB[5][21] ,
         \muxInB[5][20] , \muxInB[5][19] , \muxInB[5][18] , \muxInB[5][17] ,
         \muxInB[5][16] , \muxInB[5][15] , \muxInB[5][14] , \muxInB[5][13] ,
         \muxInB[5][12] , \muxInB[5][11] , \muxInB[5][10] , \muxInB[4][31] ,
         \muxInB[4][30] , \muxInB[4][29] , \muxInB[4][28] , \muxInB[4][27] ,
         \muxInB[4][26] , \muxInB[4][25] , \muxInB[4][24] , \muxInB[4][23] ,
         \muxInB[4][22] , \muxInB[4][21] , \muxInB[4][20] , \muxInB[4][19] ,
         \muxInB[4][18] , \muxInB[4][17] , \muxInB[4][16] , \muxInB[4][15] ,
         \muxInB[4][14] , \muxInB[4][13] , \muxInB[4][12] , \muxInB[4][11] ,
         \muxInB[4][10] , \muxInB[4][9] , \muxInB[4][8] , \muxInB[3][31] ,
         \muxInB[3][30] , \muxInB[3][29] , \muxInB[3][28] , \muxInB[3][27] ,
         \muxInB[3][26] , \muxInB[3][25] , \muxInB[3][24] , \muxInB[3][23] ,
         \muxInB[3][22] , \muxInB[3][21] , \muxInB[3][20] , \muxInB[3][19] ,
         \muxInB[3][18] , \muxInB[3][17] , \muxInB[3][16] , \muxInB[3][15] ,
         \muxInB[3][14] , \muxInB[3][13] , \muxInB[3][12] , \muxInB[3][11] ,
         \muxInB[3][10] , \muxInB[3][9] , \muxInB[3][8] , \muxInB[3][7] ,
         \muxInB[3][6] , \muxInB[2][31] , \muxInB[2][30] , \muxInB[2][29] ,
         \muxInB[2][28] , \muxInB[2][27] , \muxInB[2][26] , \muxInB[2][25] ,
         \muxInB[2][24] , \muxInB[2][23] , \muxInB[2][22] , \muxInB[2][21] ,
         \muxInB[2][20] , \muxInB[2][19] , \muxInB[2][18] , \muxInB[2][17] ,
         \muxInB[2][16] , \muxInB[2][15] , \muxInB[2][14] , \muxInB[2][13] ,
         \muxInB[2][12] , \muxInB[2][11] , \muxInB[2][10] , \muxInB[2][9] ,
         \muxInB[2][8] , \muxInB[2][7] , \muxInB[2][6] , \muxInB[2][5] ,
         \muxInB[2][4] , \muxInB[1][31] , \muxInB[1][30] , \muxInB[1][29] ,
         \muxInB[1][28] , \muxInB[1][27] , \muxInB[1][26] , \muxInB[1][25] ,
         \muxInB[1][24] , \muxInB[1][23] , \muxInB[1][22] , \muxInB[1][21] ,
         \muxInB[1][20] , \muxInB[1][19] , \muxInB[1][18] , \muxInB[1][17] ,
         \muxInB[1][16] , \muxInB[1][15] , \muxInB[1][14] , \muxInB[1][13] ,
         \muxInB[1][12] , \muxInB[1][11] , \muxInB[1][10] , \muxInB[1][9] ,
         \muxInB[1][8] , \muxInB[1][7] , \muxInB[1][6] , \muxInB[1][5] ,
         \muxInB[1][4] , \muxInB[1][3] , \muxInB[1][2] , \muxInB[0][31] ,
         \muxInB[0][30] , \muxInB[0][29] , \muxInB[0][28] , \muxInB[0][27] ,
         \muxInB[0][26] , \muxInB[0][25] , \muxInB[0][24] , \muxInB[0][23] ,
         \muxInB[0][22] , \muxInB[0][21] , \muxInB[0][20] , \muxInB[0][19] ,
         \muxInB[0][18] , \muxInB[0][17] , \muxInB[0][16] , \muxInB[0][15] ,
         \muxInB[0][14] , \muxInB[0][13] , \muxInB[0][12] , \muxInB[0][11] ,
         \muxInB[0][10] , \muxInB[0][9] , \muxInB[0][8] , \muxInB[0][7] ,
         \muxInB[0][6] , \muxInB[0][5] , \muxInB[0][4] , \muxInB[0][3] ,
         \muxInB[0][2] , \muxInB[0][1] , \muxInB[0][0] , \outmux[7][31] ,
         \outmux[7][30] , \outmux[7][29] , \outmux[7][28] , \outmux[7][27] ,
         \outmux[7][26] , \outmux[7][25] , \outmux[7][24] , \outmux[7][23] ,
         \outmux[7][22] , \outmux[7][21] , \outmux[7][20] , \outmux[7][19] ,
         \outmux[7][18] , \outmux[7][17] , \outmux[7][16] , \outmux[7][15] ,
         \outmux[7][14] , \outmux[7][13] , \outmux[7][12] , \outmux[7][11] ,
         \outmux[7][10] , \outmux[7][9] , \outmux[7][8] , \outmux[7][7] ,
         \outmux[7][6] , \outmux[7][5] , \outmux[7][4] , \outmux[7][3] ,
         \outmux[7][2] , \outmux[7][1] , \outmux[7][0] , \outmux[6][31] ,
         \outmux[6][30] , \outmux[6][29] , \outmux[6][28] , \outmux[6][27] ,
         \outmux[6][26] , \outmux[6][25] , \outmux[6][24] , \outmux[6][23] ,
         \outmux[6][22] , \outmux[6][21] , \outmux[6][20] , \outmux[6][19] ,
         \outmux[6][18] , \outmux[6][17] , \outmux[6][16] , \outmux[6][15] ,
         \outmux[6][14] , \outmux[6][13] , \outmux[6][12] , \outmux[6][11] ,
         \outmux[6][10] , \outmux[6][9] , \outmux[6][8] , \outmux[6][7] ,
         \outmux[6][6] , \outmux[6][5] , \outmux[6][4] , \outmux[6][3] ,
         \outmux[6][2] , \outmux[6][1] , \outmux[6][0] , \outmux[5][31] ,
         \outmux[5][30] , \outmux[5][29] , \outmux[5][28] , \outmux[5][27] ,
         \outmux[5][26] , \outmux[5][25] , \outmux[5][24] , \outmux[5][23] ,
         \outmux[5][22] , \outmux[5][21] , \outmux[5][20] , \outmux[5][19] ,
         \outmux[5][18] , \outmux[5][17] , \outmux[5][16] , \outmux[5][15] ,
         \outmux[5][14] , \outmux[5][13] , \outmux[5][12] , \outmux[5][11] ,
         \outmux[5][10] , \outmux[5][9] , \outmux[5][8] , \outmux[5][7] ,
         \outmux[5][6] , \outmux[5][5] , \outmux[5][4] , \outmux[5][3] ,
         \outmux[5][2] , \outmux[5][1] , \outmux[5][0] , \outmux[4][31] ,
         \outmux[4][30] , \outmux[4][29] , \outmux[4][28] , \outmux[4][27] ,
         \outmux[4][26] , \outmux[4][25] , \outmux[4][24] , \outmux[4][23] ,
         \outmux[4][22] , \outmux[4][21] , \outmux[4][20] , \outmux[4][19] ,
         \outmux[4][18] , \outmux[4][17] , \outmux[4][16] , \outmux[4][15] ,
         \outmux[4][14] , \outmux[4][13] , \outmux[4][12] , \outmux[4][11] ,
         \outmux[4][10] , \outmux[4][9] , \outmux[4][8] , \outmux[4][7] ,
         \outmux[4][6] , \outmux[4][5] , \outmux[4][4] , \outmux[4][3] ,
         \outmux[4][2] , \outmux[4][1] , \outmux[4][0] , \outmux[3][31] ,
         \outmux[3][30] , \outmux[3][29] , \outmux[3][28] , \outmux[3][27] ,
         \outmux[3][26] , \outmux[3][25] , \outmux[3][24] , \outmux[3][23] ,
         \outmux[3][22] , \outmux[3][21] , \outmux[3][20] , \outmux[3][19] ,
         \outmux[3][18] , \outmux[3][17] , \outmux[3][16] , \outmux[3][15] ,
         \outmux[3][14] , \outmux[3][13] , \outmux[3][12] , \outmux[3][11] ,
         \outmux[3][10] , \outmux[3][9] , \outmux[3][8] , \outmux[3][7] ,
         \outmux[3][6] , \outmux[3][5] , \outmux[3][4] , \outmux[3][3] ,
         \outmux[3][2] , \outmux[3][1] , \outmux[3][0] , \outmux[2][31] ,
         \outmux[2][30] , \outmux[2][29] , \outmux[2][28] , \outmux[2][27] ,
         \outmux[2][26] , \outmux[2][25] , \outmux[2][24] , \outmux[2][23] ,
         \outmux[2][22] , \outmux[2][21] , \outmux[2][20] , \outmux[2][19] ,
         \outmux[2][18] , \outmux[2][17] , \outmux[2][16] , \outmux[2][15] ,
         \outmux[2][14] , \outmux[2][13] , \outmux[2][12] , \outmux[2][11] ,
         \outmux[2][10] , \outmux[2][9] , \outmux[2][8] , \outmux[2][7] ,
         \outmux[2][6] , \outmux[2][5] , \outmux[2][4] , \outmux[2][3] ,
         \outmux[2][2] , \outmux[2][1] , \outmux[2][0] , \outmux[1][31] ,
         \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] ,
         \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] ,
         \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] ,
         \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] ,
         \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] ,
         \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] ,
         \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] ,
         \outmux[1][2] , \outmux[1][1] , \outmux[1][0] , \outmux[0][31] ,
         \outmux[0][30] , \outmux[0][29] , \outmux[0][28] , \outmux[0][27] ,
         \outmux[0][26] , \outmux[0][25] , \outmux[0][24] , \outmux[0][23] ,
         \outmux[0][22] , \outmux[0][21] , \outmux[0][20] , \outmux[0][19] ,
         \outmux[0][18] , \outmux[0][17] , \outmux[0][16] , \outmux[0][15] ,
         \outmux[0][14] , \outmux[0][13] , \outmux[0][12] , \outmux[0][11] ,
         \outmux[0][10] , \outmux[0][9] , \outmux[0][8] , \outmux[0][7] ,
         \outmux[0][6] , \outmux[0][5] , \outmux[0][4] , \outmux[0][3] ,
         \outmux[0][2] , \outmux[0][1] , \outmux[0][0] , \cout_array[5][31] ,
         \cout_array[5][30] , \cout_array[5][29] , \cout_array[5][28] ,
         \cout_array[5][27] , \cout_array[5][26] , \cout_array[5][25] ,
         \cout_array[5][24] , \cout_array[5][23] , \cout_array[5][22] ,
         \cout_array[5][21] , \cout_array[5][20] , \cout_array[5][19] ,
         \cout_array[5][18] , \cout_array[5][17] , \cout_array[5][16] ,
         \cout_array[5][15] , \cout_array[5][14] , \cout_array[5][13] ,
         \cout_array[5][12] , \cout_array[5][11] , \cout_array[5][10] ,
         \cout_array[5][9] , \cout_array[5][8] , \cout_array[5][7] ,
         \cout_array[5][6] , \cout_array[5][5] , \cout_array[5][4] ,
         \cout_array[5][3] , \cout_array[5][2] , \cout_array[5][1] ,
         \cout_array[4][31] , \cout_array[4][30] , \cout_array[4][29] ,
         \cout_array[4][28] , \cout_array[4][27] , \cout_array[4][26] ,
         \cout_array[4][25] , \cout_array[4][24] , \cout_array[4][23] ,
         \cout_array[4][22] , \cout_array[4][21] , \cout_array[4][20] ,
         \cout_array[4][19] , \cout_array[4][18] , \cout_array[4][17] ,
         \cout_array[4][16] , \cout_array[4][15] , \cout_array[4][14] ,
         \cout_array[4][13] , \cout_array[4][12] , \cout_array[4][11] ,
         \cout_array[4][10] , \cout_array[4][9] , \cout_array[4][8] ,
         \cout_array[4][7] , \cout_array[4][6] , \cout_array[4][5] ,
         \cout_array[4][4] , \cout_array[4][3] , \cout_array[4][2] ,
         \cout_array[4][1] , \cout_array[3][31] , \cout_array[3][30] ,
         \cout_array[3][29] , \cout_array[3][28] , \cout_array[3][27] ,
         \cout_array[3][26] , \cout_array[3][25] , \cout_array[3][24] ,
         \cout_array[3][23] , \cout_array[3][22] , \cout_array[3][21] ,
         \cout_array[3][20] , \cout_array[3][19] , \cout_array[3][18] ,
         \cout_array[3][17] , \cout_array[3][16] , \cout_array[3][15] ,
         \cout_array[3][14] , \cout_array[3][13] , \cout_array[3][12] ,
         \cout_array[3][11] , \cout_array[3][10] , \cout_array[3][9] ,
         \cout_array[3][8] , \cout_array[3][7] , \cout_array[3][6] ,
         \cout_array[3][5] , \cout_array[3][4] , \cout_array[3][3] ,
         \cout_array[3][2] , \cout_array[3][1] , \cout_array[2][31] ,
         \cout_array[2][30] , \cout_array[2][29] , \cout_array[2][28] ,
         \cout_array[2][27] , \cout_array[2][26] , \cout_array[2][25] ,
         \cout_array[2][24] , \cout_array[2][23] , \cout_array[2][22] ,
         \cout_array[2][21] , \cout_array[2][20] , \cout_array[2][19] ,
         \cout_array[2][18] , \cout_array[2][17] , \cout_array[2][16] ,
         \cout_array[2][15] , \cout_array[2][14] , \cout_array[2][13] ,
         \cout_array[2][12] , \cout_array[2][11] , \cout_array[2][10] ,
         \cout_array[2][9] , \cout_array[2][8] , \cout_array[2][7] ,
         \cout_array[2][6] , \cout_array[2][5] , \cout_array[2][4] ,
         \cout_array[2][3] , \cout_array[2][2] , \cout_array[2][1] ,
         \cout_array[1][31] , \cout_array[1][30] , \cout_array[1][29] ,
         \cout_array[1][28] , \cout_array[1][27] , \cout_array[1][26] ,
         \cout_array[1][25] , \cout_array[1][24] , \cout_array[1][23] ,
         \cout_array[1][22] , \cout_array[1][21] , \cout_array[1][20] ,
         \cout_array[1][19] , \cout_array[1][18] , \cout_array[1][17] ,
         \cout_array[1][16] , \cout_array[1][15] , \cout_array[1][14] ,
         \cout_array[1][13] , \cout_array[1][12] , \cout_array[1][11] ,
         \cout_array[1][10] , \cout_array[1][9] , \cout_array[1][8] ,
         \cout_array[1][7] , \cout_array[1][6] , \cout_array[1][5] ,
         \cout_array[1][4] , \cout_array[1][3] , \cout_array[1][2] ,
         \cout_array[1][1] , \cout_array[0][31] , \cout_array[0][30] ,
         \cout_array[0][29] , \cout_array[0][28] , \cout_array[0][27] ,
         \cout_array[0][26] , \cout_array[0][25] , \cout_array[0][24] ,
         \cout_array[0][23] , \cout_array[0][22] , \cout_array[0][21] ,
         \cout_array[0][20] , \cout_array[0][19] , \cout_array[0][18] ,
         \cout_array[0][17] , \cout_array[0][16] , \cout_array[0][15] ,
         \cout_array[0][14] , \cout_array[0][13] , \cout_array[0][12] ,
         \cout_array[0][11] , \cout_array[0][10] , \cout_array[0][9] ,
         \cout_array[0][8] , \cout_array[0][7] , \cout_array[0][6] ,
         \cout_array[0][5] , \cout_array[0][4] , \cout_array[0][3] ,
         \cout_array[0][2] , \cout_array[0][1] , \sum_array[5][31] ,
         \sum_array[5][30] , \sum_array[5][29] , \sum_array[5][28] ,
         \sum_array[5][27] , \sum_array[5][26] , \sum_array[5][25] ,
         \sum_array[5][24] , \sum_array[5][23] , \sum_array[5][22] ,
         \sum_array[5][21] , \sum_array[5][20] , \sum_array[5][19] ,
         \sum_array[5][18] , \sum_array[5][17] , \sum_array[5][16] ,
         \sum_array[5][15] , \sum_array[5][14] , \sum_array[5][13] ,
         \sum_array[5][12] , \sum_array[5][11] , \sum_array[5][10] ,
         \sum_array[5][9] , \sum_array[5][8] , \sum_array[5][7] ,
         \sum_array[5][6] , \sum_array[5][5] , \sum_array[5][4] ,
         \sum_array[5][3] , \sum_array[5][2] , \sum_array[5][1] ,
         \sum_array[5][0] , \sum_array[4][31] , \sum_array[4][30] ,
         \sum_array[4][29] , \sum_array[4][28] , \sum_array[4][27] ,
         \sum_array[4][26] , \sum_array[4][25] , \sum_array[4][24] ,
         \sum_array[4][23] , \sum_array[4][22] , \sum_array[4][21] ,
         \sum_array[4][20] , \sum_array[4][19] , \sum_array[4][18] ,
         \sum_array[4][17] , \sum_array[4][16] , \sum_array[4][15] ,
         \sum_array[4][14] , \sum_array[4][13] , \sum_array[4][12] ,
         \sum_array[4][11] , \sum_array[4][10] , \sum_array[4][9] ,
         \sum_array[4][8] , \sum_array[4][7] , \sum_array[4][6] ,
         \sum_array[4][5] , \sum_array[4][4] , \sum_array[4][3] ,
         \sum_array[4][2] , \sum_array[4][1] , \sum_array[4][0] ,
         \sum_array[3][31] , \sum_array[3][30] , \sum_array[3][29] ,
         \sum_array[3][28] , \sum_array[3][27] , \sum_array[3][26] ,
         \sum_array[3][25] , \sum_array[3][24] , \sum_array[3][23] ,
         \sum_array[3][22] , \sum_array[3][21] , \sum_array[3][20] ,
         \sum_array[3][19] , \sum_array[3][18] , \sum_array[3][17] ,
         \sum_array[3][16] , \sum_array[3][15] , \sum_array[3][14] ,
         \sum_array[3][13] , \sum_array[3][12] , \sum_array[3][11] ,
         \sum_array[3][10] , \sum_array[3][9] , \sum_array[3][8] ,
         \sum_array[3][7] , \sum_array[3][6] , \sum_array[3][5] ,
         \sum_array[3][4] , \sum_array[3][3] , \sum_array[3][2] ,
         \sum_array[3][1] , \sum_array[3][0] , \sum_array[2][31] ,
         \sum_array[2][30] , \sum_array[2][29] , \sum_array[2][28] ,
         \sum_array[2][27] , \sum_array[2][26] , \sum_array[2][25] ,
         \sum_array[2][24] , \sum_array[2][23] , \sum_array[2][22] ,
         \sum_array[2][21] , \sum_array[2][20] , \sum_array[2][19] ,
         \sum_array[2][18] , \sum_array[2][17] , \sum_array[2][16] ,
         \sum_array[2][15] , \sum_array[2][14] , \sum_array[2][13] ,
         \sum_array[2][12] , \sum_array[2][11] , \sum_array[2][10] ,
         \sum_array[2][9] , \sum_array[2][8] , \sum_array[2][7] ,
         \sum_array[2][6] , \sum_array[2][5] , \sum_array[2][4] ,
         \sum_array[2][3] , \sum_array[2][2] , \sum_array[2][1] ,
         \sum_array[2][0] , \sum_array[1][31] , \sum_array[1][30] ,
         \sum_array[1][29] , \sum_array[1][28] , \sum_array[1][27] ,
         \sum_array[1][26] , \sum_array[1][25] , \sum_array[1][24] ,
         \sum_array[1][23] , \sum_array[1][22] , \sum_array[1][21] ,
         \sum_array[1][20] , \sum_array[1][19] , \sum_array[1][18] ,
         \sum_array[1][17] , \sum_array[1][16] , \sum_array[1][15] ,
         \sum_array[1][14] , \sum_array[1][13] , \sum_array[1][12] ,
         \sum_array[1][11] , \sum_array[1][10] , \sum_array[1][9] ,
         \sum_array[1][8] , \sum_array[1][7] , \sum_array[1][6] ,
         \sum_array[1][5] , \sum_array[1][4] , \sum_array[1][3] ,
         \sum_array[1][2] , \sum_array[1][1] , \sum_array[1][0] ,
         \sum_array[0][31] , \sum_array[0][30] , \sum_array[0][29] ,
         \sum_array[0][28] , \sum_array[0][27] , \sum_array[0][26] ,
         \sum_array[0][25] , \sum_array[0][24] , \sum_array[0][23] ,
         \sum_array[0][22] , \sum_array[0][21] , \sum_array[0][20] ,
         \sum_array[0][19] , \sum_array[0][18] , \sum_array[0][17] ,
         \sum_array[0][16] , \sum_array[0][15] , \sum_array[0][14] ,
         \sum_array[0][13] , \sum_array[0][12] , \sum_array[0][11] ,
         \sum_array[0][10] , \sum_array[0][9] , \sum_array[0][8] ,
         \sum_array[0][7] , \sum_array[0][6] , \sum_array[0][5] ,
         \sum_array[0][4] , \sum_array[0][3] , \sum_array[0][2] ,
         \sum_array[0][1] , \sum_array[0][0] , n4, n5, n6, n7, n8, n9, n12,
         n16, n20, n23, n24, n1, n2, n3, n10, n11, n13, n14, n15, n17, n18,
         n19, n21, n22, n25, n26, n27, n28;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249;
  assign n4 = A[2];
  assign n5 = A[8];
  assign n6 = A[12];
  assign n7 = A[6];
  assign n8 = A[9];
  assign n9 = A[10];
  assign n12 = A[5];
  assign n16 = A[0];
  assign n23 = A[11];
  assign n24 = A[7];
  assign n1 = A[15];

  shift_mul_N16_S0 SHIFTERS_0 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n2}), .B({\muxInB[0][31] , 
        \muxInB[0][30] , \muxInB[0][29] , \muxInB[0][28] , \muxInB[0][27] , 
        \muxInB[0][26] , \muxInB[0][25] , \muxInB[0][24] , \muxInB[0][23] , 
        \muxInB[0][22] , \muxInB[0][21] , \muxInB[0][20] , \muxInB[0][19] , 
        \muxInB[0][18] , \muxInB[0][17] , \muxInB[0][16] , \muxInB[0][15] , 
        \muxInB[0][14] , \muxInB[0][13] , \muxInB[0][12] , \muxInB[0][11] , 
        \muxInB[0][10] , \muxInB[0][9] , \muxInB[0][8] , \muxInB[0][7] , 
        \muxInB[0][6] , \muxInB[0][5] , \muxInB[0][4] , \muxInB[0][3] , 
        \muxInB[0][2] , \muxInB[0][1] , \muxInB[0][0] }), .C({\muxInC[0][31] , 
        \muxInC[0][30] , \muxInC[0][29] , \muxInC[0][28] , \muxInC[0][27] , 
        \muxInC[0][26] , \muxInC[0][25] , \muxInC[0][24] , \muxInC[0][23] , 
        \muxInC[0][22] , \muxInC[0][21] , \muxInC[0][20] , \muxInC[0][19] , 
        \muxInC[0][18] , \muxInC[0][17] , \muxInC[0][16] , \muxInC[0][15] , 
        \muxInC[0][14] , \muxInC[0][13] , \muxInC[0][12] , \muxInC[0][11] , 
        \muxInC[0][10] , \muxInC[0][9] , \muxInC[0][8] , \muxInC[0][7] , 
        \muxInC[0][6] , \muxInC[0][5] , \muxInC[0][4] , \muxInC[0][3] , 
        \muxInC[0][2] , \muxInC[0][1] , \muxInC[0][0] }), .D({\muxInD[0][31] , 
        \muxInD[0][30] , \muxInD[0][29] , \muxInD[0][28] , \muxInD[0][27] , 
        \muxInD[0][26] , \muxInD[0][25] , \muxInD[0][24] , \muxInD[0][23] , 
        \muxInD[0][22] , \muxInD[0][21] , \muxInD[0][20] , \muxInD[0][19] , 
        \muxInD[0][18] , \muxInD[0][17] , \muxInD[0][16] , \muxInD[0][15] , 
        \muxInD[0][14] , \muxInD[0][13] , \muxInD[0][12] , \muxInD[0][11] , 
        \muxInD[0][10] , \muxInD[0][9] , \muxInD[0][8] , \muxInD[0][7] , 
        \muxInD[0][6] , \muxInD[0][5] , \muxInD[0][4] , \muxInD[0][3] , 
        \muxInD[0][2] , \muxInD[0][1] , SYNOPSYS_UNCONNECTED__0}), .E({
        \muxInE[0][31] , \muxInE[0][30] , \muxInE[0][29] , \muxInE[0][28] , 
        \muxInE[0][27] , \muxInE[0][26] , SYNOPSYS_UNCONNECTED__1, 
        \muxInE[0][24] , \muxInE[0][23] , SYNOPSYS_UNCONNECTED__2, 
        \muxInE[0][21] , \muxInE[0][20] , \muxInE[0][19] , \muxInE[0][18] , 
        SYNOPSYS_UNCONNECTED__3, \muxInE[0][16] , \muxInE[0][15] , 
        \muxInE[0][14] , \muxInE[0][13] , \muxInE[0][12] , \muxInE[0][11] , 
        \muxInE[0][10] , \muxInE[0][9] , \muxInE[0][8] , \muxInE[0][7] , 
        \muxInE[0][6] , \muxInE[0][5] , \muxInE[0][4] , \muxInE[0][3] , 
        \muxInE[0][2] , \muxInE[0][1] , SYNOPSYS_UNCONNECTED__4}) );
  shift_mul_N16_S2 SHIFTERS_1 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n2}), .B({\muxInB[1][31] , 
        \muxInB[1][30] , \muxInB[1][29] , \muxInB[1][28] , \muxInB[1][27] , 
        \muxInB[1][26] , \muxInB[1][25] , \muxInB[1][24] , \muxInB[1][23] , 
        \muxInB[1][22] , \muxInB[1][21] , \muxInB[1][20] , \muxInB[1][19] , 
        \muxInB[1][18] , \muxInB[1][17] , \muxInB[1][16] , \muxInB[1][15] , 
        \muxInB[1][14] , \muxInB[1][13] , \muxInB[1][12] , \muxInB[1][11] , 
        \muxInB[1][10] , \muxInB[1][9] , \muxInB[1][8] , \muxInB[1][7] , 
        \muxInB[1][6] , \muxInB[1][5] , \muxInB[1][4] , \muxInB[1][3] , 
        \muxInB[1][2] , SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6}), 
        .C({\muxInC[1][31] , \muxInC[1][30] , \muxInC[1][29] , \muxInC[1][28] , 
        \muxInC[1][27] , \muxInC[1][26] , \muxInC[1][25] , \muxInC[1][24] , 
        \muxInC[1][23] , \muxInC[1][22] , \muxInC[1][21] , \muxInC[1][20] , 
        SYNOPSYS_UNCONNECTED__7, \muxInC[1][18] , \muxInC[1][17] , 
        \muxInC[1][16] , \muxInC[1][15] , \muxInC[1][14] , \muxInC[1][13] , 
        \muxInC[1][12] , \muxInC[1][11] , \muxInC[1][10] , \muxInC[1][9] , 
        \muxInC[1][8] , \muxInC[1][7] , \muxInC[1][6] , \muxInC[1][5] , 
        \muxInC[1][4] , \muxInC[1][3] , \muxInC[1][2] , 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9}), .D({
        \muxInD[1][31] , \muxInD[1][30] , \muxInD[1][29] , \muxInD[1][28] , 
        \muxInD[1][27] , \muxInD[1][26] , \muxInD[1][25] , \muxInD[1][24] , 
        \muxInD[1][23] , \muxInD[1][22] , \muxInD[1][21] , \muxInD[1][20] , 
        \muxInD[1][19] , \muxInD[1][18] , \muxInD[1][17] , \muxInD[1][16] , 
        \muxInD[1][15] , \muxInD[1][14] , \muxInD[1][13] , \muxInD[1][12] , 
        \muxInD[1][11] , \muxInD[1][10] , \muxInD[1][9] , \muxInD[1][8] , 
        \muxInD[1][7] , \muxInD[1][6] , \muxInD[1][5] , \muxInD[1][4] , 
        \muxInD[1][3] , SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12}), .E({\muxInE[1][31] , \muxInE[1][30] , 
        \muxInE[1][29] , \muxInE[1][28] , \muxInE[1][27] , \muxInE[1][26] , 
        \muxInE[1][25] , \muxInE[1][24] , \muxInE[1][23] , \muxInE[1][22] , 
        \muxInE[1][21] , \muxInE[1][20] , \muxInE[1][19] , \muxInE[1][18] , 
        \muxInE[1][17] , \muxInE[1][16] , \muxInE[1][15] , \muxInE[1][14] , 
        \muxInE[1][13] , \muxInE[1][12] , \muxInE[1][11] , \muxInE[1][10] , 
        \muxInE[1][9] , \muxInE[1][8] , \muxInE[1][7] , \muxInE[1][6] , 
        \muxInE[1][5] , \muxInE[1][4] , \muxInE[1][3] , 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15}) );
  shift_mul_N16_S4 SHIFTERS_2 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n2}), .B({\muxInB[2][31] , 
        \muxInB[2][30] , \muxInB[2][29] , \muxInB[2][28] , \muxInB[2][27] , 
        \muxInB[2][26] , \muxInB[2][25] , \muxInB[2][24] , \muxInB[2][23] , 
        \muxInB[2][22] , \muxInB[2][21] , \muxInB[2][20] , \muxInB[2][19] , 
        \muxInB[2][18] , \muxInB[2][17] , \muxInB[2][16] , \muxInB[2][15] , 
        \muxInB[2][14] , \muxInB[2][13] , \muxInB[2][12] , \muxInB[2][11] , 
        \muxInB[2][10] , \muxInB[2][9] , \muxInB[2][8] , \muxInB[2][7] , 
        \muxInB[2][6] , \muxInB[2][5] , \muxInB[2][4] , 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19}), .C({
        \muxInC[2][31] , \muxInC[2][30] , \muxInC[2][29] , \muxInC[2][28] , 
        \muxInC[2][27] , \muxInC[2][26] , \muxInC[2][25] , \muxInC[2][24] , 
        \muxInC[2][23] , \muxInC[2][22] , \muxInC[2][21] , \muxInC[2][20] , 
        \muxInC[2][19] , \muxInC[2][18] , \muxInC[2][17] , \muxInC[2][16] , 
        \muxInC[2][15] , \muxInC[2][14] , \muxInC[2][13] , \muxInC[2][12] , 
        \muxInC[2][11] , \muxInC[2][10] , \muxInC[2][9] , \muxInC[2][8] , 
        \muxInC[2][7] , \muxInC[2][6] , \muxInC[2][5] , \muxInC[2][4] , 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}), .D({
        \muxInD[2][31] , \muxInD[2][30] , \muxInD[2][29] , \muxInD[2][28] , 
        \muxInD[2][27] , \muxInD[2][26] , \muxInD[2][25] , \muxInD[2][24] , 
        \muxInD[2][23] , \muxInD[2][22] , \muxInD[2][21] , \muxInD[2][20] , 
        \muxInD[2][19] , \muxInD[2][18] , \muxInD[2][17] , \muxInD[2][16] , 
        \muxInD[2][15] , \muxInD[2][14] , \muxInD[2][13] , \muxInD[2][12] , 
        \muxInD[2][11] , \muxInD[2][10] , \muxInD[2][9] , \muxInD[2][8] , 
        \muxInD[2][7] , \muxInD[2][6] , \muxInD[2][5] , 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28}), .E({\muxInE[2][31] , \muxInE[2][30] , 
        \muxInE[2][29] , \muxInE[2][28] , \muxInE[2][27] , \muxInE[2][26] , 
        \muxInE[2][25] , \muxInE[2][24] , \muxInE[2][23] , \muxInE[2][22] , 
        \muxInE[2][21] , n20, \muxInE[2][19] , \muxInE[2][18] , 
        \muxInE[2][17] , \muxInE[2][16] , \muxInE[2][15] , \muxInE[2][14] , 
        \muxInE[2][13] , \muxInE[2][12] , \muxInE[2][11] , \muxInE[2][10] , 
        \muxInE[2][9] , \muxInE[2][8] , \muxInE[2][7] , \muxInE[2][6] , 
        \muxInE[2][5] , SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33}) );
  shift_mul_N16_S6 SHIFTERS_3 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n3}), .B({\muxInB[3][31] , 
        \muxInB[3][30] , \muxInB[3][29] , \muxInB[3][28] , \muxInB[3][27] , 
        \muxInB[3][26] , \muxInB[3][25] , \muxInB[3][24] , \muxInB[3][23] , 
        \muxInB[3][22] , \muxInB[3][21] , \muxInB[3][20] , \muxInB[3][19] , 
        \muxInB[3][18] , \muxInB[3][17] , \muxInB[3][16] , \muxInB[3][15] , 
        \muxInB[3][14] , \muxInB[3][13] , \muxInB[3][12] , \muxInB[3][11] , 
        \muxInB[3][10] , \muxInB[3][9] , \muxInB[3][8] , \muxInB[3][7] , 
        \muxInB[3][6] , SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}), .C({
        \muxInC[3][31] , \muxInC[3][30] , \muxInC[3][29] , \muxInC[3][28] , 
        \muxInC[3][27] , \muxInC[3][26] , \muxInC[3][25] , \muxInC[3][24] , 
        \muxInC[3][23] , \muxInC[3][22] , \muxInC[3][21] , \muxInC[3][20] , 
        \muxInC[3][19] , \muxInC[3][18] , \muxInC[3][17] , \muxInC[3][16] , 
        \muxInC[3][15] , \muxInC[3][14] , \muxInC[3][13] , \muxInC[3][12] , 
        \muxInC[3][11] , \muxInC[3][10] , \muxInC[3][9] , \muxInC[3][8] , 
        \muxInC[3][7] , \muxInC[3][6] , SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45}), .D({\muxInD[3][31] , \muxInD[3][30] , 
        \muxInD[3][29] , \muxInD[3][28] , \muxInD[3][27] , \muxInD[3][26] , 
        \muxInD[3][25] , \muxInD[3][24] , \muxInD[3][23] , \muxInD[3][22] , 
        \muxInD[3][21] , \muxInD[3][20] , \muxInD[3][19] , \muxInD[3][18] , 
        \muxInD[3][17] , \muxInD[3][16] , \muxInD[3][15] , \muxInD[3][14] , 
        \muxInD[3][13] , \muxInD[3][12] , \muxInD[3][11] , \muxInD[3][10] , 
        \muxInD[3][9] , \muxInD[3][8] , \muxInD[3][7] , 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52}), .E({\muxInE[3][31] , \muxInE[3][30] , 
        \muxInE[3][29] , \muxInE[3][28] , \muxInE[3][27] , \muxInE[3][26] , 
        \muxInE[3][25] , \muxInE[3][24] , \muxInE[3][23] , \muxInE[3][22] , 
        \muxInE[3][21] , \muxInE[3][20] , \muxInE[3][19] , \muxInE[3][18] , 
        \muxInE[3][17] , \muxInE[3][16] , \muxInE[3][15] , \muxInE[3][14] , 
        \muxInE[3][13] , \muxInE[3][12] , \muxInE[3][11] , \muxInE[3][10] , 
        \muxInE[3][9] , \muxInE[3][8] , \muxInE[3][7] , 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59}) );
  shift_mul_N16_S8 SHIFTERS_4 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n2}), .B({\muxInB[4][31] , 
        \muxInB[4][30] , \muxInB[4][29] , \muxInB[4][28] , \muxInB[4][27] , 
        \muxInB[4][26] , \muxInB[4][25] , \muxInB[4][24] , \muxInB[4][23] , 
        \muxInB[4][22] , \muxInB[4][21] , \muxInB[4][20] , \muxInB[4][19] , 
        \muxInB[4][18] , \muxInB[4][17] , \muxInB[4][16] , \muxInB[4][15] , 
        \muxInB[4][14] , \muxInB[4][13] , \muxInB[4][12] , \muxInB[4][11] , 
        \muxInB[4][10] , \muxInB[4][9] , \muxInB[4][8] , 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67}), .C({
        \muxInC[4][31] , \muxInC[4][30] , \muxInC[4][29] , \muxInC[4][28] , 
        \muxInC[4][27] , \muxInC[4][26] , \muxInC[4][25] , \muxInC[4][24] , 
        \muxInC[4][23] , \muxInC[4][22] , \muxInC[4][21] , \muxInC[4][20] , 
        \muxInC[4][19] , \muxInC[4][18] , \muxInC[4][17] , \muxInC[4][16] , 
        \muxInC[4][15] , \muxInC[4][14] , \muxInC[4][13] , \muxInC[4][12] , 
        \muxInC[4][11] , \muxInC[4][10] , \muxInC[4][9] , \muxInC[4][8] , 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75}), .D({
        \muxInD[4][31] , \muxInD[4][30] , \muxInD[4][29] , \muxInD[4][28] , 
        \muxInD[4][27] , \muxInD[4][26] , \muxInD[4][25] , \muxInD[4][24] , 
        \muxInD[4][23] , \muxInD[4][22] , \muxInD[4][21] , \muxInD[4][20] , 
        \muxInD[4][19] , \muxInD[4][18] , \muxInD[4][17] , \muxInD[4][16] , 
        \muxInD[4][15] , \muxInD[4][14] , \muxInD[4][13] , \muxInD[4][12] , 
        \muxInD[4][11] , \muxInD[4][10] , \muxInD[4][9] , 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84}), .E({\muxInE[4][31] , \muxInE[4][30] , 
        \muxInE[4][29] , \muxInE[4][28] , \muxInE[4][27] , \muxInE[4][26] , 
        \muxInE[4][25] , \muxInE[4][24] , \muxInE[4][23] , \muxInE[4][22] , 
        \muxInE[4][21] , \muxInE[4][20] , \muxInE[4][19] , \muxInE[4][18] , 
        \muxInE[4][17] , \muxInE[4][16] , \muxInE[4][15] , \muxInE[4][14] , 
        \muxInE[4][13] , \muxInE[4][12] , \muxInE[4][11] , \muxInE[4][10] , 
        \muxInE[4][9] , SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93}) );
  shift_mul_N16_S10 SHIFTERS_5 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n3}), .B({\muxInB[5][31] , 
        \muxInB[5][30] , \muxInB[5][29] , \muxInB[5][28] , \muxInB[5][27] , 
        \muxInB[5][26] , \muxInB[5][25] , \muxInB[5][24] , \muxInB[5][23] , 
        \muxInB[5][22] , \muxInB[5][21] , \muxInB[5][20] , \muxInB[5][19] , 
        \muxInB[5][18] , \muxInB[5][17] , \muxInB[5][16] , \muxInB[5][15] , 
        \muxInB[5][14] , \muxInB[5][13] , \muxInB[5][12] , \muxInB[5][11] , 
        \muxInB[5][10] , SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103}), .C({
        \muxInC[5][31] , \muxInC[5][30] , \muxInC[5][29] , \muxInC[5][28] , 
        \muxInC[5][27] , \muxInC[5][26] , \muxInC[5][25] , \muxInC[5][24] , 
        \muxInC[5][23] , \muxInC[5][22] , \muxInC[5][21] , \muxInC[5][20] , 
        \muxInC[5][19] , \muxInC[5][18] , \muxInC[5][17] , \muxInC[5][16] , 
        \muxInC[5][15] , \muxInC[5][14] , \muxInC[5][13] , \muxInC[5][12] , 
        \muxInC[5][11] , \muxInC[5][10] , SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113}), .D({\muxInD[5][31] , \muxInD[5][30] , 
        \muxInD[5][29] , \muxInD[5][28] , \muxInD[5][27] , \muxInD[5][26] , 
        \muxInD[5][25] , \muxInD[5][24] , \muxInD[5][23] , \muxInD[5][22] , 
        \muxInD[5][21] , \muxInD[5][20] , \muxInD[5][19] , \muxInD[5][18] , 
        \muxInD[5][17] , \muxInD[5][16] , \muxInD[5][15] , \muxInD[5][14] , 
        \muxInD[5][13] , \muxInD[5][12] , \muxInD[5][11] , 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124}), .E({\muxInE[5][31] , \muxInE[5][30] , 
        \muxInE[5][29] , \muxInE[5][28] , \muxInE[5][27] , \muxInE[5][26] , 
        \muxInE[5][25] , \muxInE[5][24] , \muxInE[5][23] , \muxInE[5][22] , 
        \muxInE[5][21] , \muxInE[5][20] , \muxInE[5][19] , \muxInE[5][18] , 
        \muxInE[5][17] , \muxInE[5][16] , \muxInE[5][15] , \muxInE[5][14] , 
        \muxInE[5][13] , \muxInE[5][12] , \muxInE[5][11] , 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135}) );
  shift_mul_N16_S12 SHIFTERS_6 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n3}), .B({\muxInB[6][31] , 
        \muxInB[6][30] , \muxInB[6][29] , \muxInB[6][28] , \muxInB[6][27] , 
        \muxInB[6][26] , \muxInB[6][25] , \muxInB[6][24] , \muxInB[6][23] , 
        \muxInB[6][22] , \muxInB[6][21] , \muxInB[6][20] , \muxInB[6][19] , 
        \muxInB[6][18] , \muxInB[6][17] , \muxInB[6][16] , \muxInB[6][15] , 
        \muxInB[6][14] , \muxInB[6][13] , \muxInB[6][12] , 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147}), .C({
        \muxInC[6][31] , \muxInC[6][30] , \muxInC[6][29] , \muxInC[6][28] , 
        \muxInC[6][27] , \muxInC[6][26] , \muxInC[6][25] , \muxInC[6][24] , 
        \muxInC[6][23] , \muxInC[6][22] , \muxInC[6][21] , \muxInC[6][20] , 
        \muxInC[6][19] , \muxInC[6][18] , \muxInC[6][17] , \muxInC[6][16] , 
        \muxInC[6][15] , \muxInC[6][14] , \muxInC[6][13] , \muxInC[6][12] , 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159}), .D({
        \muxInD[6][31] , \muxInD[6][30] , \muxInD[6][29] , \muxInD[6][28] , 
        \muxInD[6][27] , \muxInD[6][26] , \muxInD[6][25] , \muxInD[6][24] , 
        \muxInD[6][23] , \muxInD[6][22] , \muxInD[6][21] , \muxInD[6][20] , 
        \muxInD[6][19] , \muxInD[6][18] , \muxInD[6][17] , \muxInD[6][16] , 
        \muxInD[6][15] , \muxInD[6][14] , \muxInD[6][13] , 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172}), .E({\muxInE[6][31] , \muxInE[6][30] , 
        \muxInE[6][29] , \muxInE[6][28] , \muxInE[6][27] , \muxInE[6][26] , 
        \muxInE[6][25] , \muxInE[6][24] , \muxInE[6][23] , \muxInE[6][22] , 
        \muxInE[6][21] , \muxInE[6][20] , \muxInE[6][19] , \muxInE[6][18] , 
        \muxInE[6][17] , \muxInE[6][16] , \muxInE[6][15] , \muxInE[6][14] , 
        \muxInE[6][13] , SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185}) );
  shift_mul_N16_S14 SHIFTERS_7 ( .A({n28, n27, n26, n25, n22, n21, n19, n18, 
        n17, n15, n14, n13, n11, n4, n10, n2}), .B({\muxInB[7][31] , 
        \muxInB[7][30] , \muxInB[7][29] , \muxInB[7][28] , \muxInB[7][27] , 
        \muxInB[7][26] , \muxInB[7][25] , \muxInB[7][24] , \muxInB[7][23] , 
        \muxInB[7][22] , \muxInB[7][21] , \muxInB[7][20] , \muxInB[7][19] , 
        \muxInB[7][18] , \muxInB[7][17] , \muxInB[7][16] , \muxInB[7][15] , 
        \muxInB[7][14] , SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199}), .C({
        \muxInC[7][31] , \muxInC[7][30] , \muxInC[7][29] , \muxInC[7][28] , 
        \muxInC[7][27] , \muxInC[7][26] , \muxInC[7][25] , \muxInC[7][24] , 
        \muxInC[7][23] , \muxInC[7][22] , \muxInC[7][21] , \muxInC[7][20] , 
        \muxInC[7][19] , \muxInC[7][18] , \muxInC[7][17] , \muxInC[7][16] , 
        \muxInC[7][15] , \muxInC[7][14] , SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, 
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213}), .D({\muxInD[7][31] , \muxInD[7][30] , 
        \muxInD[7][29] , \muxInD[7][28] , \muxInD[7][27] , \muxInD[7][26] , 
        \muxInD[7][25] , \muxInD[7][24] , \muxInD[7][23] , \muxInD[7][22] , 
        \muxInD[7][21] , \muxInD[7][20] , \muxInD[7][19] , \muxInD[7][18] , 
        \muxInD[7][17] , \muxInD[7][16] , \muxInD[7][15] , 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228}), .E({\muxInE[7][31] , \muxInE[7][30] , 
        \muxInE[7][29] , \muxInE[7][28] , \muxInE[7][27] , \muxInE[7][26] , 
        \muxInE[7][25] , \muxInE[7][24] , \muxInE[7][23] , \muxInE[7][22] , 
        \muxInE[7][21] , \muxInE[7][20] , \muxInE[7][19] , \muxInE[7][18] , 
        \muxInE[7][17] , \muxInE[7][16] , \muxInE[7][15] , 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, 
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243}) );
  mux_N32_0 MUXGEN_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[0][31] , \muxInB[0][30] , \muxInB[0][29] , \muxInB[0][28] , 
        \muxInB[0][27] , \muxInB[0][26] , \muxInB[0][25] , \muxInB[0][24] , 
        \muxInB[0][23] , \muxInB[0][22] , \muxInB[0][21] , \muxInB[0][20] , 
        \muxInB[0][19] , \muxInB[0][18] , \muxInB[0][17] , \muxInB[0][16] , 
        \muxInB[0][15] , \muxInB[0][14] , \muxInB[0][13] , \muxInB[0][12] , 
        \muxInB[0][11] , \muxInB[0][10] , \muxInB[0][9] , \muxInB[0][8] , 
        \muxInB[0][7] , \muxInB[0][6] , \muxInB[0][5] , \muxInB[0][4] , 
        \muxInB[0][3] , \muxInB[0][2] , \muxInB[0][1] , \muxInB[0][0] }), .C({
        \muxInC[0][31] , \muxInC[0][30] , \muxInC[0][29] , \muxInC[0][28] , 
        \muxInC[0][20] , \muxInC[0][26] , \muxInC[0][25] , \muxInC[0][24] , 
        \muxInC[0][23] , \muxInC[0][22] , \muxInC[0][21] , \muxInC[0][20] , 
        \muxInC[0][19] , \muxInC[0][18] , \muxInC[0][17] , \muxInC[0][16] , 
        \muxInC[0][15] , \muxInC[0][14] , \muxInC[0][13] , \muxInC[0][12] , 
        \muxInC[0][11] , \muxInC[0][10] , \muxInC[0][9] , \muxInC[0][8] , 
        \muxInC[0][7] , \muxInC[0][6] , \muxInC[0][5] , \muxInC[0][4] , 
        \muxInC[0][3] , \muxInC[0][2] , \muxInC[0][1] , \muxInC[0][0] }), .D({
        \muxInD[0][31] , \muxInD[0][30] , \muxInD[0][29] , \muxInD[0][28] , 
        \muxInD[0][27] , \muxInD[0][26] , \muxInD[0][25] , \muxInD[0][24] , 
        \muxInD[0][23] , \muxInD[0][22] , \muxInD[0][21] , \muxInD[0][20] , 
        \muxInD[0][19] , \muxInD[0][18] , \muxInD[0][17] , \muxInD[0][16] , 
        \muxInD[0][15] , \muxInD[0][14] , \muxInD[0][13] , \muxInD[0][12] , 
        \muxInD[0][11] , \muxInD[0][10] , \muxInD[0][9] , \muxInD[0][8] , 
        \muxInD[0][7] , \muxInD[0][6] , \muxInD[0][5] , \muxInD[0][4] , 
        \muxInD[0][3] , \muxInD[0][2] , \muxInD[0][1] , 1'b0}), .E({
        \muxInE[0][31] , \muxInE[0][30] , \muxInE[0][29] , \muxInE[0][28] , 
        \muxInE[0][27] , \muxInE[0][26] , \muxInC[0][20] , \muxInE[0][24] , 
        \muxInE[0][23] , \muxInC[0][27] , \muxInE[0][21] , \muxInE[0][20] , 
        \muxInE[0][19] , \muxInE[0][18] , \muxInC[0][29] , \muxInE[0][16] , 
        \muxInE[0][15] , \muxInE[0][14] , \muxInE[0][13] , \muxInE[0][12] , 
        \muxInE[0][11] , \muxInE[0][10] , \muxInE[0][9] , \muxInE[0][8] , 
        \muxInE[0][7] , \muxInE[0][6] , \muxInE[0][5] , \muxInE[0][4] , 
        \muxInE[0][3] , \muxInE[0][2] , \muxInE[0][1] , 1'b0}), .Sel({B[1:0], 
        1'b0}), .O({\outmux[0][31] , \outmux[0][30] , \outmux[0][29] , 
        \outmux[0][28] , \outmux[0][27] , \outmux[0][26] , \outmux[0][25] , 
        \outmux[0][24] , \outmux[0][23] , \outmux[0][22] , \outmux[0][21] , 
        \outmux[0][20] , \outmux[0][19] , \outmux[0][18] , \outmux[0][17] , 
        \outmux[0][16] , \outmux[0][15] , \outmux[0][14] , \outmux[0][13] , 
        \outmux[0][12] , \outmux[0][11] , \outmux[0][10] , \outmux[0][9] , 
        \outmux[0][8] , \outmux[0][7] , \outmux[0][6] , \outmux[0][5] , 
        \outmux[0][4] , \outmux[0][3] , \outmux[0][2] , \outmux[0][1] , 
        \outmux[0][0] }) );
  mux_N32_7 MUXGEN_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[1][31] , \muxInB[1][30] , \muxInB[1][29] , \muxInB[1][28] , 
        \muxInB[1][27] , \muxInB[1][26] , \muxInB[1][25] , \muxInB[1][24] , 
        \muxInB[1][23] , \muxInB[1][22] , \muxInB[1][21] , \muxInB[1][20] , 
        \muxInB[1][19] , \muxInB[1][18] , \muxInB[1][17] , \muxInB[1][16] , 
        \muxInB[1][15] , \muxInB[1][14] , \muxInB[1][13] , \muxInB[1][12] , 
        \muxInB[1][11] , \muxInB[1][10] , \muxInB[1][9] , \muxInB[1][8] , 
        \muxInB[1][7] , \muxInB[1][6] , \muxInB[1][5] , \muxInB[1][4] , 
        \muxInB[1][3] , \muxInB[1][2] , 1'b0, 1'b0}), .C({\muxInC[1][31] , 
        \muxInC[1][30] , \muxInC[1][29] , \muxInC[1][28] , \muxInC[1][27] , 
        \muxInC[1][26] , \muxInC[1][25] , \muxInC[1][24] , \muxInE[1][23] , 
        \muxInC[1][22] , \muxInC[1][21] , \muxInC[1][20] , \muxInC[1][23] , 
        \muxInC[1][18] , \muxInC[1][17] , \muxInC[1][16] , \muxInC[1][15] , 
        \muxInC[1][14] , \muxInC[1][13] , \muxInC[1][12] , \muxInC[1][11] , 
        \muxInC[1][10] , \muxInC[1][9] , \muxInC[1][8] , \muxInC[1][7] , 
        \muxInC[1][6] , \muxInC[1][5] , \muxInC[1][4] , \muxInC[1][3] , 
        \muxInC[1][2] , 1'b0, 1'b0}), .D({\muxInD[1][31] , \muxInD[1][30] , 
        \muxInD[1][29] , \muxInD[1][28] , \muxInD[1][27] , \muxInD[1][26] , 
        \muxInD[1][25] , \muxInD[1][24] , \muxInD[1][23] , \muxInD[1][22] , 
        \muxInD[1][21] , \muxInD[1][20] , \muxInD[1][19] , \muxInD[1][18] , 
        \muxInD[1][17] , \muxInD[1][16] , \muxInD[1][15] , \muxInD[1][14] , 
        \muxInD[1][13] , \muxInD[1][12] , \muxInD[1][11] , \muxInD[1][10] , 
        \muxInD[1][9] , \muxInD[1][8] , \muxInD[1][7] , \muxInD[1][6] , 
        \muxInD[1][5] , \muxInD[1][4] , \muxInD[1][3] , 1'b0, 1'b0, 1'b0}), 
        .E({\muxInE[1][31] , \muxInE[1][30] , \muxInE[1][29] , \muxInE[1][28] , 
        \muxInE[1][27] , \muxInE[1][26] , \muxInE[1][25] , \muxInE[1][24] , 
        \muxInE[1][23] , \muxInE[1][22] , \muxInE[1][21] , \muxInE[1][20] , 
        \muxInE[1][19] , \muxInE[1][18] , \muxInE[1][17] , \muxInE[1][16] , 
        \muxInE[1][15] , \muxInE[1][14] , \muxInE[1][13] , \muxInE[1][12] , 
        \muxInE[1][11] , \muxInE[1][10] , \muxInE[1][9] , \muxInE[1][8] , 
        \muxInE[1][7] , \muxInE[1][6] , \muxInE[1][5] , \muxInE[1][4] , 
        \muxInE[1][3] , 1'b0, 1'b0, 1'b0}), .Sel(B[3:1]), .O({\outmux[1][31] , 
        \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , 
        \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , 
        \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , 
        \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , 
        \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , 
        \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , 
        \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }) );
  mux_N32_6 MUXGEN_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[2][31] , \muxInB[2][30] , \muxInB[2][29] , \muxInB[2][28] , 
        \muxInB[2][27] , \muxInB[2][26] , \muxInB[2][25] , \muxInB[2][24] , 
        \muxInB[2][23] , \muxInB[2][22] , \muxInB[2][21] , \muxInB[2][20] , 
        \muxInB[2][19] , \muxInB[2][18] , \muxInB[2][17] , \muxInB[2][16] , 
        \muxInB[2][15] , \muxInB[2][14] , \muxInB[2][13] , \muxInB[2][12] , 
        \muxInB[2][11] , \muxInB[2][10] , \muxInB[2][9] , \muxInB[2][8] , 
        \muxInB[2][7] , \muxInB[2][6] , \muxInB[2][5] , \muxInB[2][4] , 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({\muxInC[2][31] , \muxInC[2][30] , 
        \muxInC[2][29] , \muxInC[2][28] , \muxInC[2][27] , \muxInC[2][26] , 
        \muxInC[2][25] , \muxInC[2][24] , \muxInC[2][23] , \muxInC[2][22] , 
        \muxInC[2][21] , \muxInC[2][20] , n20, \muxInC[2][18] , 
        \muxInC[2][17] , \muxInC[2][16] , \muxInC[2][15] , \muxInC[2][14] , 
        \muxInC[2][13] , \muxInC[2][12] , \muxInC[2][11] , \muxInC[2][10] , 
        \muxInC[2][9] , \muxInC[2][8] , \muxInC[2][7] , \muxInC[2][6] , 
        \muxInC[2][5] , \muxInC[2][4] , 1'b0, 1'b0, 1'b0, 1'b0}), .D({
        \muxInD[2][31] , \muxInD[2][30] , \muxInD[2][29] , \muxInD[2][28] , 
        \muxInD[2][27] , \muxInD[2][26] , \muxInD[2][25] , \muxInD[2][24] , 
        \muxInD[2][23] , \muxInD[2][22] , \muxInD[2][21] , \muxInD[2][20] , 
        \muxInD[2][19] , \muxInD[2][18] , \muxInD[2][17] , \muxInD[2][16] , 
        \muxInD[2][15] , \muxInD[2][14] , \muxInD[2][13] , \muxInD[2][12] , 
        \muxInD[2][11] , \muxInD[2][10] , \muxInD[2][9] , \muxInD[2][8] , 
        \muxInD[2][7] , \muxInD[2][6] , \muxInD[2][5] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\muxInE[2][31] , \muxInE[2][30] , \muxInE[2][29] , 
        \muxInE[2][28] , \muxInE[2][27] , \muxInE[2][26] , \muxInE[2][25] , 
        \muxInE[2][24] , \muxInE[2][23] , \muxInE[2][22] , \muxInE[2][21] , 
        \muxInC[2][19] , \muxInE[2][19] , \muxInE[2][18] , \muxInE[2][17] , 
        \muxInE[2][16] , \muxInE[2][15] , \muxInE[2][14] , \muxInE[2][13] , 
        \muxInE[2][12] , \muxInE[2][11] , \muxInE[2][10] , \muxInE[2][9] , 
        \muxInE[2][8] , \muxInE[2][7] , \muxInE[2][6] , \muxInE[2][5] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .Sel(B[5:3]), .O({\outmux[2][31] , 
        \outmux[2][30] , \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , 
        \outmux[2][26] , \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , 
        \outmux[2][22] , \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , 
        \outmux[2][18] , \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , 
        \outmux[2][14] , \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , 
        \outmux[2][10] , \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , 
        \outmux[2][6] , \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , 
        \outmux[2][2] , \outmux[2][1] , \outmux[2][0] }) );
  mux_N32_5 MUXGEN_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[3][31] , \muxInB[3][30] , \muxInB[3][29] , \muxInB[3][28] , 
        \muxInB[3][27] , \muxInB[3][26] , \muxInB[3][25] , \muxInB[3][24] , 
        \muxInB[3][23] , \muxInB[3][22] , \muxInB[3][21] , \muxInB[3][20] , 
        \muxInB[3][19] , \muxInB[3][18] , \muxInB[3][17] , \muxInB[3][16] , 
        \muxInB[3][15] , \muxInB[3][14] , \muxInB[3][13] , \muxInB[3][12] , 
        \muxInB[3][11] , \muxInB[3][10] , \muxInB[3][9] , \muxInB[3][8] , 
        \muxInB[3][7] , \muxInB[3][6] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .C({\muxInC[3][31] , \muxInC[3][30] , \muxInC[3][29] , \muxInC[3][28] , 
        \muxInC[3][27] , \muxInC[3][26] , \muxInC[3][25] , \muxInC[3][24] , 
        \muxInC[3][23] , \muxInC[3][22] , \muxInC[3][21] , \muxInC[3][20] , 
        \muxInC[3][19] , \muxInC[3][18] , \muxInC[3][17] , \muxInC[3][16] , 
        \muxInC[3][15] , \muxInC[3][14] , \muxInC[3][13] , \muxInC[3][12] , 
        \muxInC[3][11] , \muxInC[3][10] , \muxInC[3][9] , \muxInC[3][8] , 
        \muxInC[3][7] , \muxInC[3][6] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .D({\muxInD[3][31] , \muxInD[3][30] , \muxInD[3][29] , \muxInD[3][28] , 
        \muxInD[3][27] , \muxInD[3][26] , \muxInD[3][25] , \muxInD[3][24] , 
        \muxInD[3][23] , \muxInD[3][22] , \muxInD[3][21] , \muxInD[3][20] , 
        \muxInD[3][19] , \muxInD[3][18] , \muxInD[3][17] , \muxInD[3][16] , 
        \muxInD[3][15] , \muxInD[3][14] , \muxInD[3][13] , \muxInD[3][12] , 
        \muxInD[3][11] , \muxInD[3][10] , \muxInD[3][9] , \muxInD[3][8] , 
        \muxInD[3][7] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({
        \muxInE[3][31] , \muxInE[3][30] , \muxInE[3][29] , \muxInE[3][28] , 
        \muxInE[3][27] , \muxInE[3][26] , \muxInE[3][25] , \muxInE[3][24] , 
        \muxInE[3][23] , \muxInE[3][22] , \muxInE[3][21] , \muxInE[3][20] , 
        \muxInE[3][19] , \muxInE[3][18] , \muxInE[3][17] , \muxInE[3][16] , 
        \muxInE[3][15] , \muxInE[3][14] , \muxInE[3][13] , \muxInE[3][12] , 
        \muxInE[3][11] , \muxInE[3][10] , \muxInE[3][9] , \muxInE[3][8] , 
        \muxInE[3][7] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Sel(
        B[7:5]), .O({\outmux[3][31] , \outmux[3][30] , \outmux[3][29] , 
        \outmux[3][28] , \outmux[3][27] , \outmux[3][26] , \outmux[3][25] , 
        \outmux[3][24] , \outmux[3][23] , \outmux[3][22] , \outmux[3][21] , 
        \outmux[3][20] , \outmux[3][19] , \outmux[3][18] , \outmux[3][17] , 
        \outmux[3][16] , \outmux[3][15] , \outmux[3][14] , \outmux[3][13] , 
        \outmux[3][12] , \outmux[3][11] , \outmux[3][10] , \outmux[3][9] , 
        \outmux[3][8] , \outmux[3][7] , \outmux[3][6] , \outmux[3][5] , 
        \outmux[3][4] , \outmux[3][3] , \outmux[3][2] , \outmux[3][1] , 
        \outmux[3][0] }) );
  mux_N32_4 MUXGEN_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[4][31] , \muxInB[4][30] , \muxInB[4][29] , \muxInB[4][28] , 
        \muxInB[4][27] , \muxInB[4][26] , \muxInB[4][25] , \muxInB[4][24] , 
        \muxInB[4][23] , \muxInB[4][22] , \muxInB[4][21] , \muxInB[4][20] , 
        \muxInB[4][19] , \muxInB[4][18] , \muxInB[4][17] , \muxInB[4][16] , 
        \muxInB[4][15] , \muxInB[4][14] , \muxInB[4][13] , \muxInB[4][12] , 
        \muxInB[4][11] , \muxInB[4][10] , \muxInB[4][9] , \muxInB[4][8] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({\muxInC[4][31] , 
        \muxInC[4][30] , \muxInC[4][29] , \muxInC[4][28] , \muxInC[4][27] , 
        \muxInC[4][26] , \muxInC[4][25] , \muxInC[4][24] , \muxInC[4][23] , 
        \muxInC[4][22] , \muxInC[4][21] , \muxInC[4][20] , \muxInC[4][19] , 
        \muxInC[4][18] , \muxInC[4][17] , \muxInC[4][16] , \muxInC[4][15] , 
        \muxInC[4][14] , \muxInC[4][13] , \muxInC[4][12] , \muxInC[4][11] , 
        \muxInC[4][10] , \muxInC[4][9] , \muxInC[4][8] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({\muxInD[4][31] , \muxInD[4][30] , 
        \muxInD[4][29] , \muxInD[4][28] , \muxInD[4][27] , \muxInD[4][26] , 
        \muxInD[4][25] , \muxInD[4][24] , \muxInD[4][23] , \muxInD[4][22] , 
        \muxInD[4][21] , \muxInD[4][20] , \muxInD[4][19] , \muxInD[4][18] , 
        \muxInD[4][17] , \muxInD[4][16] , \muxInD[4][15] , \muxInD[4][14] , 
        \muxInD[4][13] , \muxInD[4][12] , \muxInD[4][11] , \muxInD[4][10] , 
        \muxInD[4][9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({\muxInE[4][31] , \muxInE[4][30] , \muxInE[4][29] , \muxInE[4][28] , 
        \muxInE[4][27] , \muxInE[4][26] , \muxInE[4][25] , \muxInE[4][24] , 
        \muxInE[4][23] , \muxInE[4][22] , \muxInE[4][21] , \muxInE[4][20] , 
        \muxInE[4][19] , \muxInE[4][18] , \muxInE[4][17] , \muxInE[4][16] , 
        \muxInE[4][15] , \muxInE[4][14] , \muxInE[4][13] , \muxInE[4][12] , 
        \muxInE[4][11] , \muxInE[4][10] , \muxInE[4][9] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Sel(B[9:7]), .O({
        \outmux[4][31] , \outmux[4][30] , \outmux[4][29] , \outmux[4][28] , 
        \outmux[4][27] , \outmux[4][26] , \outmux[4][25] , \outmux[4][24] , 
        \outmux[4][23] , \outmux[4][22] , \outmux[4][21] , \outmux[4][20] , 
        \outmux[4][19] , \outmux[4][18] , \outmux[4][17] , \outmux[4][16] , 
        \outmux[4][15] , \outmux[4][14] , \outmux[4][13] , \outmux[4][12] , 
        \outmux[4][11] , \outmux[4][10] , \outmux[4][9] , \outmux[4][8] , 
        \outmux[4][7] , \outmux[4][6] , \outmux[4][5] , \outmux[4][4] , 
        \outmux[4][3] , \outmux[4][2] , \outmux[4][1] , \outmux[4][0] }) );
  mux_N32_3 MUXGEN_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[5][31] , \muxInB[5][30] , \muxInB[5][29] , \muxInB[5][28] , 
        \muxInB[5][27] , \muxInB[5][26] , \muxInB[5][25] , \muxInB[5][24] , 
        \muxInB[5][23] , \muxInB[5][22] , \muxInB[5][21] , \muxInB[5][20] , 
        \muxInB[5][19] , \muxInB[5][18] , \muxInB[5][17] , \muxInB[5][16] , 
        \muxInB[5][15] , \muxInB[5][14] , \muxInB[5][13] , \muxInB[5][12] , 
        \muxInB[5][11] , \muxInB[5][10] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .C({\muxInC[5][31] , \muxInC[5][30] , 
        \muxInC[5][29] , \muxInC[5][28] , \muxInC[5][27] , \muxInC[5][26] , 
        \muxInC[5][25] , \muxInC[5][24] , \muxInC[5][23] , \muxInC[5][22] , 
        \muxInC[5][21] , \muxInC[5][20] , \muxInC[5][19] , \muxInC[5][18] , 
        \muxInC[5][17] , \muxInC[5][16] , \muxInC[5][15] , \muxInC[5][14] , 
        \muxInC[5][13] , \muxInC[5][12] , \muxInC[5][11] , \muxInC[5][10] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({
        \muxInD[5][31] , \muxInD[5][30] , \muxInD[5][29] , \muxInD[5][28] , 
        \muxInD[5][27] , \muxInD[5][26] , \muxInD[5][25] , \muxInD[5][24] , 
        \muxInD[5][23] , \muxInD[5][22] , \muxInD[5][21] , \muxInD[5][20] , 
        \muxInD[5][19] , \muxInD[5][18] , \muxInD[5][17] , \muxInD[5][16] , 
        \muxInD[5][15] , \muxInD[5][14] , \muxInD[5][13] , \muxInD[5][12] , 
        \muxInD[5][11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .E({\muxInE[5][31] , \muxInE[5][30] , \muxInE[5][29] , 
        \muxInE[5][28] , \muxInE[5][27] , \muxInE[5][26] , \muxInE[5][25] , 
        \muxInE[5][24] , \muxInE[5][23] , \muxInE[5][22] , \muxInE[5][21] , 
        \muxInE[5][20] , \muxInE[5][19] , \muxInE[5][18] , \muxInE[5][17] , 
        \muxInE[5][16] , \muxInE[5][15] , \muxInE[5][14] , \muxInE[5][13] , 
        \muxInE[5][12] , \muxInE[5][11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Sel(B[11:9]), .O({\outmux[5][31] , 
        \outmux[5][30] , \outmux[5][29] , \outmux[5][28] , \outmux[5][27] , 
        \outmux[5][26] , \outmux[5][25] , \outmux[5][24] , \outmux[5][23] , 
        \outmux[5][22] , \outmux[5][21] , \outmux[5][20] , \outmux[5][19] , 
        \outmux[5][18] , \outmux[5][17] , \outmux[5][16] , \outmux[5][15] , 
        \outmux[5][14] , \outmux[5][13] , \outmux[5][12] , \outmux[5][11] , 
        \outmux[5][10] , \outmux[5][9] , \outmux[5][8] , \outmux[5][7] , 
        \outmux[5][6] , \outmux[5][5] , \outmux[5][4] , \outmux[5][3] , 
        \outmux[5][2] , \outmux[5][1] , \outmux[5][0] }) );
  mux_N32_2 MUXGEN_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[6][31] , \muxInB[6][30] , \muxInB[6][29] , \muxInB[6][28] , 
        \muxInB[6][27] , \muxInB[6][26] , \muxInB[6][25] , \muxInB[6][24] , 
        \muxInB[6][23] , \muxInB[6][22] , \muxInB[6][21] , \muxInB[6][20] , 
        \muxInB[6][19] , \muxInB[6][18] , \muxInB[6][17] , \muxInB[6][16] , 
        \muxInB[6][15] , \muxInB[6][14] , \muxInB[6][13] , \muxInB[6][12] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({\muxInC[6][31] , \muxInC[6][30] , \muxInC[6][29] , \muxInC[6][28] , 
        \muxInC[6][27] , \muxInC[6][26] , \muxInC[6][25] , \muxInC[6][24] , 
        \muxInC[6][23] , \muxInC[6][22] , \muxInC[6][21] , \muxInC[6][20] , 
        \muxInC[6][19] , \muxInC[6][18] , \muxInC[6][17] , \muxInC[6][16] , 
        \muxInC[6][15] , \muxInC[6][14] , \muxInC[6][13] , \muxInC[6][12] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({\muxInD[6][31] , \muxInD[6][30] , \muxInD[6][29] , \muxInD[6][28] , 
        \muxInD[6][27] , \muxInD[6][26] , \muxInD[6][25] , \muxInD[6][24] , 
        \muxInD[6][23] , \muxInD[6][22] , \muxInD[6][21] , \muxInD[6][20] , 
        \muxInD[6][19] , \muxInD[6][18] , \muxInD[6][17] , \muxInD[6][16] , 
        \muxInD[6][15] , \muxInD[6][14] , \muxInD[6][13] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({
        \muxInE[6][31] , \muxInE[6][30] , \muxInE[6][29] , \muxInE[6][28] , 
        \muxInE[6][27] , \muxInE[6][26] , \muxInE[6][25] , \muxInE[6][24] , 
        \muxInE[6][23] , \muxInE[6][22] , \muxInE[6][21] , \muxInE[6][20] , 
        \muxInE[6][19] , \muxInE[6][18] , \muxInE[6][17] , \muxInE[6][16] , 
        \muxInE[6][15] , \muxInE[6][14] , \muxInE[6][13] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Sel(
        B[13:11]), .O({\outmux[6][31] , \outmux[6][30] , \outmux[6][29] , 
        \outmux[6][28] , \outmux[6][27] , \outmux[6][26] , \outmux[6][25] , 
        \outmux[6][24] , \outmux[6][23] , \outmux[6][22] , \outmux[6][21] , 
        \outmux[6][20] , \outmux[6][19] , \outmux[6][18] , \outmux[6][17] , 
        \outmux[6][16] , \outmux[6][15] , \outmux[6][14] , \outmux[6][13] , 
        \outmux[6][12] , \outmux[6][11] , \outmux[6][10] , \outmux[6][9] , 
        \outmux[6][8] , \outmux[6][7] , \outmux[6][6] , \outmux[6][5] , 
        \outmux[6][4] , \outmux[6][3] , \outmux[6][2] , \outmux[6][1] , 
        \outmux[6][0] }) );
  mux_N32_1 MUXGEN_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\muxInB[7][31] , \muxInB[7][30] , \muxInB[7][29] , \muxInB[7][28] , 
        \muxInB[7][27] , \muxInB[7][26] , \muxInB[7][25] , \muxInB[7][24] , 
        \muxInB[7][23] , \muxInB[7][22] , \muxInB[7][21] , \muxInB[7][20] , 
        \muxInB[7][19] , \muxInB[7][18] , \muxInB[7][17] , \muxInB[7][16] , 
        \muxInB[7][15] , \muxInB[7][14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({\muxInC[7][31] , 
        \muxInC[7][30] , \muxInC[7][29] , \muxInC[7][28] , \muxInC[7][27] , 
        \muxInC[7][26] , \muxInC[7][25] , \muxInC[7][24] , \muxInC[7][23] , 
        \muxInC[7][22] , \muxInC[7][21] , \muxInC[7][20] , \muxInC[7][19] , 
        \muxInC[7][18] , \muxInC[7][17] , \muxInC[7][16] , \muxInC[7][15] , 
        \muxInC[7][14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({\muxInD[7][31] , \muxInD[7][30] , 
        \muxInD[7][29] , \muxInD[7][28] , \muxInD[7][27] , \muxInD[7][26] , 
        \muxInD[7][25] , \muxInD[7][24] , \muxInD[7][23] , \muxInD[7][22] , 
        \muxInD[7][21] , \muxInD[7][20] , \muxInD[7][19] , \muxInD[7][18] , 
        \muxInD[7][17] , \muxInD[7][16] , \muxInD[7][15] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({\muxInE[7][31] , \muxInE[7][30] , \muxInE[7][29] , \muxInE[7][28] , 
        \muxInE[7][27] , \muxInE[7][26] , \muxInE[7][25] , \muxInE[7][24] , 
        \muxInE[7][23] , \muxInE[7][22] , \muxInE[7][21] , \muxInE[7][20] , 
        \muxInE[7][19] , \muxInE[7][18] , \muxInE[7][17] , \muxInE[7][16] , 
        \muxInE[7][15] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Sel(B[15:13]), .O({
        \outmux[7][31] , \outmux[7][30] , \outmux[7][29] , \outmux[7][28] , 
        \outmux[7][27] , \outmux[7][26] , \outmux[7][25] , \outmux[7][24] , 
        \outmux[7][23] , \outmux[7][22] , \outmux[7][21] , \outmux[7][20] , 
        \outmux[7][19] , \outmux[7][18] , \outmux[7][17] , \outmux[7][16] , 
        \outmux[7][15] , \outmux[7][14] , \outmux[7][13] , \outmux[7][12] , 
        \outmux[7][11] , \outmux[7][10] , \outmux[7][9] , \outmux[7][8] , 
        \outmux[7][7] , \outmux[7][6] , \outmux[7][5] , \outmux[7][4] , 
        \outmux[7][3] , \outmux[7][2] , \outmux[7][1] , \outmux[7][0] }) );
  CSA_Nbits32_0 Add1IL ( .A({\outmux[0][31] , \outmux[0][30] , \outmux[0][29] , 
        \outmux[0][28] , \outmux[0][27] , \outmux[0][26] , \outmux[0][25] , 
        \outmux[0][24] , \outmux[0][23] , \outmux[0][22] , \outmux[0][21] , 
        \outmux[0][20] , \outmux[0][19] , \outmux[0][18] , \outmux[0][17] , 
        \outmux[0][16] , \outmux[0][15] , \outmux[0][14] , \outmux[0][13] , 
        \outmux[0][12] , \outmux[0][11] , \outmux[0][10] , \outmux[0][9] , 
        \outmux[0][8] , \outmux[0][7] , \outmux[0][6] , \outmux[0][5] , 
        \outmux[0][4] , \outmux[0][3] , \outmux[0][2] , \outmux[0][1] , 
        \outmux[0][0] }), .B({\outmux[1][31] , \outmux[1][30] , 
        \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , \outmux[1][26] , 
        \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , \outmux[1][22] , 
        \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , \outmux[1][18] , 
        \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , \outmux[1][14] , 
        \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , \outmux[1][10] , 
        \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , \outmux[1][6] , 
        \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , \outmux[1][2] , 
        \outmux[1][1] , \outmux[1][0] }), .C({\outmux[2][31] , \outmux[2][30] , 
        \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , \outmux[2][26] , 
        \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , \outmux[2][22] , 
        \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , \outmux[2][18] , 
        \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , \outmux[2][14] , 
        \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , \outmux[2][10] , 
        \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , \outmux[2][6] , 
        \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , \outmux[2][2] , 
        \outmux[2][1] , \outmux[2][0] }), .S({\sum_array[0][31] , 
        \sum_array[0][30] , \sum_array[0][29] , \sum_array[0][28] , 
        \sum_array[0][27] , \sum_array[0][26] , \sum_array[0][25] , 
        \sum_array[0][24] , \sum_array[0][23] , \sum_array[0][22] , 
        \sum_array[0][21] , \sum_array[0][20] , \sum_array[0][19] , 
        \sum_array[0][18] , \sum_array[0][17] , \sum_array[0][16] , 
        \sum_array[0][15] , \sum_array[0][14] , \sum_array[0][13] , 
        \sum_array[0][12] , \sum_array[0][11] , \sum_array[0][10] , 
        \sum_array[0][9] , \sum_array[0][8] , \sum_array[0][7] , 
        \sum_array[0][6] , \sum_array[0][5] , \sum_array[0][4] , 
        \sum_array[0][3] , \sum_array[0][2] , \sum_array[0][1] , 
        \sum_array[0][0] }), .Cout({\cout_array[0][31] , \cout_array[0][30] , 
        \cout_array[0][29] , \cout_array[0][28] , \cout_array[0][27] , 
        \cout_array[0][26] , \cout_array[0][25] , \cout_array[0][24] , 
        \cout_array[0][23] , \cout_array[0][22] , \cout_array[0][21] , 
        \cout_array[0][20] , \cout_array[0][19] , \cout_array[0][18] , 
        \cout_array[0][17] , \cout_array[0][16] , \cout_array[0][15] , 
        \cout_array[0][14] , \cout_array[0][13] , \cout_array[0][12] , 
        \cout_array[0][11] , \cout_array[0][10] , \cout_array[0][9] , 
        \cout_array[0][8] , \cout_array[0][7] , \cout_array[0][6] , 
        \cout_array[0][5] , \cout_array[0][4] , \cout_array[0][3] , 
        \cout_array[0][2] , \cout_array[0][1] , SYNOPSYS_UNCONNECTED__244}) );
  CSA_Nbits32_5 Add2IL ( .A({\outmux[3][31] , \outmux[3][30] , \outmux[3][29] , 
        \outmux[3][28] , \outmux[3][27] , \outmux[3][26] , \outmux[3][25] , 
        \outmux[3][24] , \outmux[3][23] , \outmux[3][22] , \outmux[3][21] , 
        \outmux[3][20] , \outmux[3][19] , \outmux[3][18] , \outmux[3][17] , 
        \outmux[3][16] , \outmux[3][15] , \outmux[3][14] , \outmux[3][13] , 
        \outmux[3][12] , \outmux[3][11] , \outmux[3][10] , \outmux[3][9] , 
        \outmux[3][8] , \outmux[3][7] , \outmux[3][6] , \outmux[3][5] , 
        \outmux[3][4] , \outmux[3][3] , \outmux[3][2] , \outmux[3][1] , 
        \outmux[3][0] }), .B({\outmux[4][31] , \outmux[4][30] , 
        \outmux[4][29] , \outmux[4][28] , \outmux[4][27] , \outmux[4][26] , 
        \outmux[4][25] , \outmux[4][24] , \outmux[4][23] , \outmux[4][22] , 
        \outmux[4][21] , \outmux[4][20] , \outmux[4][19] , \outmux[4][18] , 
        \outmux[4][17] , \outmux[4][16] , \outmux[4][15] , \outmux[4][14] , 
        \outmux[4][13] , \outmux[4][12] , \outmux[4][11] , \outmux[4][10] , 
        \outmux[4][9] , \outmux[4][8] , \outmux[4][7] , \outmux[4][6] , 
        \outmux[4][5] , \outmux[4][4] , \outmux[4][3] , \outmux[4][2] , 
        \outmux[4][1] , \outmux[4][0] }), .C({\outmux[5][31] , \outmux[5][30] , 
        \outmux[5][29] , \outmux[5][28] , \outmux[5][27] , \outmux[5][26] , 
        \outmux[5][25] , \outmux[5][24] , \outmux[5][23] , \outmux[5][22] , 
        \outmux[5][21] , \outmux[5][20] , \outmux[5][19] , \outmux[5][18] , 
        \outmux[5][17] , \outmux[5][16] , \outmux[5][15] , \outmux[5][14] , 
        \outmux[5][13] , \outmux[5][12] , \outmux[5][11] , \outmux[5][10] , 
        \outmux[5][9] , \outmux[5][8] , \outmux[5][7] , \outmux[5][6] , 
        \outmux[5][5] , \outmux[5][4] , \outmux[5][3] , \outmux[5][2] , 
        \outmux[5][1] , \outmux[5][0] }), .S({\sum_array[1][31] , 
        \sum_array[1][30] , \sum_array[1][29] , \sum_array[1][28] , 
        \sum_array[1][27] , \sum_array[1][26] , \sum_array[1][25] , 
        \sum_array[1][24] , \sum_array[1][23] , \sum_array[1][22] , 
        \sum_array[1][21] , \sum_array[1][20] , \sum_array[1][19] , 
        \sum_array[1][18] , \sum_array[1][17] , \sum_array[1][16] , 
        \sum_array[1][15] , \sum_array[1][14] , \sum_array[1][13] , 
        \sum_array[1][12] , \sum_array[1][11] , \sum_array[1][10] , 
        \sum_array[1][9] , \sum_array[1][8] , \sum_array[1][7] , 
        \sum_array[1][6] , \sum_array[1][5] , \sum_array[1][4] , 
        \sum_array[1][3] , \sum_array[1][2] , \sum_array[1][1] , 
        \sum_array[1][0] }), .Cout({\cout_array[1][31] , \cout_array[1][30] , 
        \cout_array[1][29] , \cout_array[1][28] , \cout_array[1][27] , 
        \cout_array[1][26] , \cout_array[1][25] , \cout_array[1][24] , 
        \cout_array[1][23] , \cout_array[1][22] , \cout_array[1][21] , 
        \cout_array[1][20] , \cout_array[1][19] , \cout_array[1][18] , 
        \cout_array[1][17] , \cout_array[1][16] , \cout_array[1][15] , 
        \cout_array[1][14] , \cout_array[1][13] , \cout_array[1][12] , 
        \cout_array[1][11] , \cout_array[1][10] , \cout_array[1][9] , 
        \cout_array[1][8] , \cout_array[1][7] , \cout_array[1][6] , 
        \cout_array[1][5] , \cout_array[1][4] , \cout_array[1][3] , 
        \cout_array[1][2] , \cout_array[1][1] , SYNOPSYS_UNCONNECTED__245}) );
  CSA_Nbits32_4 Add1IIL ( .A({\sum_array[0][31] , \sum_array[0][30] , 
        \sum_array[0][29] , \sum_array[0][28] , \sum_array[0][27] , 
        \sum_array[0][26] , \sum_array[0][25] , \sum_array[0][24] , 
        \sum_array[0][23] , \sum_array[0][22] , \sum_array[0][21] , 
        \sum_array[0][20] , \sum_array[0][19] , \sum_array[0][18] , 
        \sum_array[0][17] , \sum_array[0][16] , \sum_array[0][15] , 
        \sum_array[0][14] , \sum_array[0][13] , \sum_array[0][12] , 
        \sum_array[0][11] , \sum_array[0][10] , \sum_array[0][9] , 
        \sum_array[0][8] , \sum_array[0][7] , \sum_array[0][6] , 
        \sum_array[0][5] , \sum_array[0][4] , \sum_array[0][3] , 
        \sum_array[0][2] , \sum_array[0][1] , \sum_array[0][0] }), .B({
        \cout_array[0][31] , \cout_array[0][30] , \cout_array[0][29] , 
        \cout_array[0][28] , \cout_array[0][27] , \cout_array[0][26] , 
        \cout_array[0][25] , \cout_array[0][24] , \cout_array[0][23] , 
        \cout_array[0][22] , \cout_array[0][21] , \cout_array[0][20] , 
        \cout_array[0][19] , \cout_array[0][18] , \cout_array[0][17] , 
        \cout_array[0][16] , \cout_array[0][15] , \cout_array[0][14] , 
        \cout_array[0][13] , \cout_array[0][12] , \cout_array[0][11] , 
        \cout_array[0][10] , \cout_array[0][9] , \cout_array[0][8] , 
        \cout_array[0][7] , \cout_array[0][6] , \cout_array[0][5] , 
        \cout_array[0][4] , \cout_array[0][3] , \cout_array[0][2] , 
        \cout_array[0][1] , 1'b0}), .C({\sum_array[1][31] , \sum_array[1][30] , 
        \sum_array[1][29] , \sum_array[1][28] , \sum_array[1][27] , 
        \sum_array[1][26] , \sum_array[1][25] , \sum_array[1][24] , 
        \sum_array[1][23] , \sum_array[1][22] , \sum_array[1][21] , 
        \sum_array[1][20] , \sum_array[1][19] , \sum_array[1][18] , 
        \sum_array[1][17] , \sum_array[1][16] , \sum_array[1][15] , 
        \sum_array[1][14] , \sum_array[1][13] , \sum_array[1][12] , 
        \sum_array[1][11] , \sum_array[1][10] , \sum_array[1][9] , 
        \sum_array[1][8] , \sum_array[1][7] , \sum_array[1][6] , 
        \sum_array[1][5] , \sum_array[1][4] , \sum_array[1][3] , 
        \sum_array[1][2] , \sum_array[1][1] , \sum_array[1][0] }), .S({
        \sum_array[2][31] , \sum_array[2][30] , \sum_array[2][29] , 
        \sum_array[2][28] , \sum_array[2][27] , \sum_array[2][26] , 
        \sum_array[2][25] , \sum_array[2][24] , \sum_array[2][23] , 
        \sum_array[2][22] , \sum_array[2][21] , \sum_array[2][20] , 
        \sum_array[2][19] , \sum_array[2][18] , \sum_array[2][17] , 
        \sum_array[2][16] , \sum_array[2][15] , \sum_array[2][14] , 
        \sum_array[2][13] , \sum_array[2][12] , \sum_array[2][11] , 
        \sum_array[2][10] , \sum_array[2][9] , \sum_array[2][8] , 
        \sum_array[2][7] , \sum_array[2][6] , \sum_array[2][5] , 
        \sum_array[2][4] , \sum_array[2][3] , \sum_array[2][2] , 
        \sum_array[2][1] , \sum_array[2][0] }), .Cout({\cout_array[2][31] , 
        \cout_array[2][30] , \cout_array[2][29] , \cout_array[2][28] , 
        \cout_array[2][27] , \cout_array[2][26] , \cout_array[2][25] , 
        \cout_array[2][24] , \cout_array[2][23] , \cout_array[2][22] , 
        \cout_array[2][21] , \cout_array[2][20] , \cout_array[2][19] , 
        \cout_array[2][18] , \cout_array[2][17] , \cout_array[2][16] , 
        \cout_array[2][15] , \cout_array[2][14] , \cout_array[2][13] , 
        \cout_array[2][12] , \cout_array[2][11] , \cout_array[2][10] , 
        \cout_array[2][9] , \cout_array[2][8] , \cout_array[2][7] , 
        \cout_array[2][6] , \cout_array[2][5] , \cout_array[2][4] , 
        \cout_array[2][3] , \cout_array[2][2] , \cout_array[2][1] , 
        SYNOPSYS_UNCONNECTED__246}) );
  CSA_Nbits32_3 Add2IIL ( .A({\cout_array[1][31] , \cout_array[1][30] , 
        \cout_array[1][29] , \cout_array[1][28] , \cout_array[1][27] , 
        \cout_array[1][26] , \cout_array[1][25] , \cout_array[1][24] , 
        \cout_array[1][23] , \cout_array[1][22] , \cout_array[1][21] , 
        \cout_array[1][20] , \cout_array[1][19] , \cout_array[1][18] , 
        \cout_array[1][17] , \cout_array[1][16] , \cout_array[1][15] , 
        \cout_array[1][14] , \cout_array[1][13] , \cout_array[1][12] , 
        \cout_array[1][11] , \cout_array[1][10] , \cout_array[1][9] , 
        \cout_array[1][8] , \cout_array[1][7] , \cout_array[1][6] , 
        \cout_array[1][5] , \cout_array[1][4] , \cout_array[1][3] , 
        \cout_array[1][2] , \cout_array[1][1] , 1'b0}), .B({\outmux[6][31] , 
        \outmux[6][30] , \outmux[6][29] , \outmux[6][28] , \outmux[6][27] , 
        \outmux[6][26] , \outmux[6][25] , \outmux[6][24] , \outmux[6][23] , 
        \outmux[6][22] , \outmux[6][21] , \outmux[6][20] , \outmux[6][19] , 
        \outmux[6][18] , \outmux[6][17] , \outmux[6][16] , \outmux[6][15] , 
        \outmux[6][14] , \outmux[6][13] , \outmux[6][12] , \outmux[6][11] , 
        \outmux[6][10] , \outmux[6][9] , \outmux[6][8] , \outmux[6][7] , 
        \outmux[6][6] , \outmux[6][5] , \outmux[6][4] , \outmux[6][3] , 
        \outmux[6][2] , \outmux[6][1] , \outmux[6][0] }), .C({\outmux[7][31] , 
        \outmux[7][30] , \outmux[7][29] , \outmux[7][28] , \outmux[7][27] , 
        \outmux[7][26] , \outmux[7][25] , \outmux[7][24] , \outmux[7][23] , 
        \outmux[7][22] , \outmux[7][21] , \outmux[7][20] , \outmux[7][19] , 
        \outmux[7][18] , \outmux[7][17] , \outmux[7][16] , \outmux[7][15] , 
        \outmux[7][14] , \outmux[7][13] , \outmux[7][12] , \outmux[7][11] , 
        \outmux[7][10] , \outmux[7][9] , \outmux[7][8] , \outmux[7][7] , 
        \outmux[7][6] , \outmux[7][5] , \outmux[7][4] , \outmux[7][3] , 
        \outmux[7][2] , \outmux[7][1] , \outmux[7][0] }), .S({
        \sum_array[3][31] , \sum_array[3][30] , \sum_array[3][29] , 
        \sum_array[3][28] , \sum_array[3][27] , \sum_array[3][26] , 
        \sum_array[3][25] , \sum_array[3][24] , \sum_array[3][23] , 
        \sum_array[3][22] , \sum_array[3][21] , \sum_array[3][20] , 
        \sum_array[3][19] , \sum_array[3][18] , \sum_array[3][17] , 
        \sum_array[3][16] , \sum_array[3][15] , \sum_array[3][14] , 
        \sum_array[3][13] , \sum_array[3][12] , \sum_array[3][11] , 
        \sum_array[3][10] , \sum_array[3][9] , \sum_array[3][8] , 
        \sum_array[3][7] , \sum_array[3][6] , \sum_array[3][5] , 
        \sum_array[3][4] , \sum_array[3][3] , \sum_array[3][2] , 
        \sum_array[3][1] , \sum_array[3][0] }), .Cout({\cout_array[3][31] , 
        \cout_array[3][30] , \cout_array[3][29] , \cout_array[3][28] , 
        \cout_array[3][27] , \cout_array[3][26] , \cout_array[3][25] , 
        \cout_array[3][24] , \cout_array[3][23] , \cout_array[3][22] , 
        \cout_array[3][21] , \cout_array[3][20] , \cout_array[3][19] , 
        \cout_array[3][18] , \cout_array[3][17] , \cout_array[3][16] , 
        \cout_array[3][15] , \cout_array[3][14] , \cout_array[3][13] , 
        \cout_array[3][12] , \cout_array[3][11] , \cout_array[3][10] , 
        \cout_array[3][9] , \cout_array[3][8] , \cout_array[3][7] , 
        \cout_array[3][6] , \cout_array[3][5] , \cout_array[3][4] , 
        \cout_array[3][3] , \cout_array[3][2] , \cout_array[3][1] , 
        SYNOPSYS_UNCONNECTED__247}) );
  CSA_Nbits32_2 Add1IIIL ( .A({\sum_array[2][31] , \sum_array[2][30] , 
        \sum_array[2][29] , \sum_array[2][28] , \sum_array[2][27] , 
        \sum_array[2][26] , \sum_array[2][25] , \sum_array[2][24] , 
        \sum_array[2][23] , \sum_array[2][22] , \sum_array[2][21] , 
        \sum_array[2][20] , \sum_array[2][19] , \sum_array[2][18] , 
        \sum_array[2][17] , \sum_array[2][16] , \sum_array[2][15] , 
        \sum_array[2][14] , \sum_array[2][13] , \sum_array[2][12] , 
        \sum_array[2][11] , \sum_array[2][10] , \sum_array[2][9] , 
        \sum_array[2][8] , \sum_array[2][7] , \sum_array[2][6] , 
        \sum_array[2][5] , \sum_array[2][4] , \sum_array[2][3] , 
        \sum_array[2][2] , \sum_array[2][1] , \sum_array[2][0] }), .B({
        \cout_array[2][31] , \cout_array[2][30] , \cout_array[2][29] , 
        \cout_array[2][28] , \cout_array[2][27] , \cout_array[2][26] , 
        \cout_array[2][25] , \cout_array[2][24] , \cout_array[2][23] , 
        \cout_array[2][22] , \cout_array[2][21] , \cout_array[2][20] , 
        \cout_array[2][19] , \cout_array[2][18] , \cout_array[2][17] , 
        \cout_array[2][16] , \cout_array[2][15] , \cout_array[2][14] , 
        \cout_array[2][13] , \cout_array[2][12] , \cout_array[2][11] , 
        \cout_array[2][10] , \cout_array[2][9] , \cout_array[2][8] , 
        \cout_array[2][7] , \cout_array[2][6] , \cout_array[2][5] , 
        \cout_array[2][4] , \cout_array[2][3] , \cout_array[2][2] , 
        \cout_array[2][1] , 1'b0}), .C({\sum_array[3][31] , \sum_array[3][30] , 
        \sum_array[3][29] , \sum_array[3][28] , \sum_array[3][27] , 
        \sum_array[3][26] , \sum_array[3][25] , \sum_array[3][24] , 
        \sum_array[3][23] , \sum_array[3][22] , \sum_array[3][21] , 
        \sum_array[3][20] , \sum_array[3][19] , \sum_array[3][18] , 
        \sum_array[3][17] , \sum_array[3][16] , \sum_array[3][15] , 
        \sum_array[3][14] , \sum_array[3][13] , \sum_array[3][12] , 
        \sum_array[3][11] , \sum_array[3][10] , \sum_array[3][9] , 
        \sum_array[3][8] , \sum_array[3][7] , \sum_array[3][6] , 
        \sum_array[3][5] , \sum_array[3][4] , \sum_array[3][3] , 
        \sum_array[3][2] , \sum_array[3][1] , \sum_array[3][0] }), .S({
        \sum_array[4][31] , \sum_array[4][30] , \sum_array[4][29] , 
        \sum_array[4][28] , \sum_array[4][27] , \sum_array[4][26] , 
        \sum_array[4][25] , \sum_array[4][24] , \sum_array[4][23] , 
        \sum_array[4][22] , \sum_array[4][21] , \sum_array[4][20] , 
        \sum_array[4][19] , \sum_array[4][18] , \sum_array[4][17] , 
        \sum_array[4][16] , \sum_array[4][15] , \sum_array[4][14] , 
        \sum_array[4][13] , \sum_array[4][12] , \sum_array[4][11] , 
        \sum_array[4][10] , \sum_array[4][9] , \sum_array[4][8] , 
        \sum_array[4][7] , \sum_array[4][6] , \sum_array[4][5] , 
        \sum_array[4][4] , \sum_array[4][3] , \sum_array[4][2] , 
        \sum_array[4][1] , \sum_array[4][0] }), .Cout({\cout_array[4][31] , 
        \cout_array[4][30] , \cout_array[4][29] , \cout_array[4][28] , 
        \cout_array[4][27] , \cout_array[4][26] , \cout_array[4][25] , 
        \cout_array[4][24] , \cout_array[4][23] , \cout_array[4][22] , 
        \cout_array[4][21] , \cout_array[4][20] , \cout_array[4][19] , 
        \cout_array[4][18] , \cout_array[4][17] , \cout_array[4][16] , 
        \cout_array[4][15] , \cout_array[4][14] , \cout_array[4][13] , 
        \cout_array[4][12] , \cout_array[4][11] , \cout_array[4][10] , 
        \cout_array[4][9] , \cout_array[4][8] , \cout_array[4][7] , 
        \cout_array[4][6] , \cout_array[4][5] , \cout_array[4][4] , 
        \cout_array[4][3] , \cout_array[4][2] , \cout_array[4][1] , 
        SYNOPSYS_UNCONNECTED__248}) );
  CSA_Nbits32_1 AddRCA ( .A({\sum_array[4][31] , \sum_array[4][30] , 
        \sum_array[4][29] , \sum_array[4][28] , \sum_array[4][27] , 
        \sum_array[4][26] , \sum_array[4][25] , \sum_array[4][24] , 
        \sum_array[4][23] , \sum_array[4][22] , \sum_array[4][21] , 
        \sum_array[4][20] , \sum_array[4][19] , \sum_array[4][18] , 
        \sum_array[4][17] , \sum_array[4][16] , \sum_array[4][15] , 
        \sum_array[4][14] , \sum_array[4][13] , \sum_array[4][12] , 
        \sum_array[4][11] , \sum_array[4][10] , \sum_array[4][9] , 
        \sum_array[4][8] , \sum_array[4][7] , \sum_array[4][6] , 
        \sum_array[4][5] , \sum_array[4][4] , \sum_array[4][3] , 
        \sum_array[4][2] , \sum_array[4][1] , \sum_array[4][0] }), .B({
        \cout_array[4][31] , \cout_array[4][30] , \cout_array[4][29] , 
        \cout_array[4][28] , \cout_array[4][27] , \cout_array[4][26] , 
        \cout_array[4][25] , \cout_array[4][24] , \cout_array[4][23] , 
        \cout_array[4][22] , \cout_array[4][21] , \cout_array[4][20] , 
        \cout_array[4][19] , \cout_array[4][18] , \cout_array[4][17] , 
        \cout_array[4][16] , \cout_array[4][15] , \cout_array[4][14] , 
        \cout_array[4][13] , \cout_array[4][12] , \cout_array[4][11] , 
        \cout_array[4][10] , \cout_array[4][9] , \cout_array[4][8] , 
        \cout_array[4][7] , \cout_array[4][6] , \cout_array[4][5] , 
        \cout_array[4][4] , \cout_array[4][3] , \cout_array[4][2] , 
        \cout_array[4][1] , 1'b0}), .C({\cout_array[3][31] , 
        \cout_array[3][30] , \cout_array[3][29] , \cout_array[3][28] , 
        \cout_array[3][27] , \cout_array[3][26] , \cout_array[3][25] , 
        \cout_array[3][24] , \cout_array[3][23] , \cout_array[3][22] , 
        \cout_array[3][21] , \cout_array[3][20] , \cout_array[3][19] , 
        \cout_array[3][18] , \cout_array[3][17] , \cout_array[3][16] , 
        \cout_array[3][15] , \cout_array[3][14] , \cout_array[3][13] , 
        \cout_array[3][12] , \cout_array[3][11] , \cout_array[3][10] , 
        \cout_array[3][9] , \cout_array[3][8] , \cout_array[3][7] , 
        \cout_array[3][6] , \cout_array[3][5] , \cout_array[3][4] , 
        \cout_array[3][3] , \cout_array[3][2] , \cout_array[3][1] , 1'b0}), 
        .S({\sum_array[5][31] , \sum_array[5][30] , \sum_array[5][29] , 
        \sum_array[5][28] , \sum_array[5][27] , \sum_array[5][26] , 
        \sum_array[5][25] , \sum_array[5][24] , \sum_array[5][23] , 
        \sum_array[5][22] , \sum_array[5][21] , \sum_array[5][20] , 
        \sum_array[5][19] , \sum_array[5][18] , \sum_array[5][17] , 
        \sum_array[5][16] , \sum_array[5][15] , \sum_array[5][14] , 
        \sum_array[5][13] , \sum_array[5][12] , \sum_array[5][11] , 
        \sum_array[5][10] , \sum_array[5][9] , \sum_array[5][8] , 
        \sum_array[5][7] , \sum_array[5][6] , \sum_array[5][5] , 
        \sum_array[5][4] , \sum_array[5][3] , \sum_array[5][2] , 
        \sum_array[5][1] , \sum_array[5][0] }), .Cout({\cout_array[5][31] , 
        \cout_array[5][30] , \cout_array[5][29] , \cout_array[5][28] , 
        \cout_array[5][27] , \cout_array[5][26] , \cout_array[5][25] , 
        \cout_array[5][24] , \cout_array[5][23] , \cout_array[5][22] , 
        \cout_array[5][21] , \cout_array[5][20] , \cout_array[5][19] , 
        \cout_array[5][18] , \cout_array[5][17] , \cout_array[5][16] , 
        \cout_array[5][15] , \cout_array[5][14] , \cout_array[5][13] , 
        \cout_array[5][12] , \cout_array[5][11] , \cout_array[5][10] , 
        \cout_array[5][9] , \cout_array[5][8] , \cout_array[5][7] , 
        \cout_array[5][6] , \cout_array[5][5] , \cout_array[5][4] , 
        \cout_array[5][3] , \cout_array[5][2] , \cout_array[5][1] , 
        SYNOPSYS_UNCONNECTED__249}) );
  cla_adder_N32_1 P4adder ( .A({\sum_array[5][31] , \sum_array[5][30] , 
        \sum_array[5][29] , \sum_array[5][28] , \sum_array[5][27] , 
        \sum_array[5][26] , \sum_array[5][25] , \sum_array[5][24] , 
        \sum_array[5][23] , \sum_array[5][22] , \sum_array[5][21] , 
        \sum_array[5][20] , \sum_array[5][19] , \sum_array[5][18] , 
        \sum_array[5][17] , \sum_array[5][16] , \sum_array[5][15] , 
        \sum_array[5][14] , \sum_array[5][13] , \sum_array[5][12] , 
        \sum_array[5][11] , \sum_array[5][10] , \sum_array[5][9] , 
        \sum_array[5][8] , \sum_array[5][7] , \sum_array[5][6] , 
        \sum_array[5][5] , \sum_array[5][4] , \sum_array[5][3] , 
        \sum_array[5][2] , \sum_array[5][1] , \sum_array[5][0] }), .B({
        \cout_array[5][31] , \cout_array[5][30] , \cout_array[5][29] , 
        \cout_array[5][28] , \cout_array[5][27] , \cout_array[5][26] , 
        \cout_array[5][25] , \cout_array[5][24] , \cout_array[5][23] , 
        \cout_array[5][22] , \cout_array[5][21] , \cout_array[5][20] , 
        \cout_array[5][19] , \cout_array[5][18] , \cout_array[5][17] , 
        \cout_array[5][16] , \cout_array[5][15] , \cout_array[5][14] , 
        \cout_array[5][13] , \cout_array[5][12] , \cout_array[5][11] , 
        \cout_array[5][10] , \cout_array[5][9] , \cout_array[5][8] , 
        \cout_array[5][7] , \cout_array[5][6] , \cout_array[5][5] , 
        \cout_array[5][4] , \cout_array[5][3] , \cout_array[5][2] , 
        \cout_array[5][1] , 1'b0}), .Ci(1'b0), .Sum(Y) );
  BUF_X1 U248 ( .A(n6), .Z(n25) );
  BUF_X1 U249 ( .A(n5), .Z(n18) );
  BUF_X1 U250 ( .A(n23), .Z(n22) );
  BUF_X1 U251 ( .A(A[14]), .Z(n27) );
  BUF_X1 U252 ( .A(n9), .Z(n21) );
  BUF_X2 U253 ( .A(A[13]), .Z(n26) );
  BUF_X2 U254 ( .A(n8), .Z(n19) );
  BUF_X2 U255 ( .A(A[3]), .Z(n11) );
  BUF_X2 U256 ( .A(n24), .Z(n17) );
  BUF_X2 U257 ( .A(A[1]), .Z(n10) );
  BUF_X2 U258 ( .A(n16), .Z(n2) );
  BUF_X2 U259 ( .A(n12), .Z(n14) );
  BUF_X1 U260 ( .A(n7), .Z(n15) );
  BUF_X1 U261 ( .A(n16), .Z(n3) );
  BUF_X1 U262 ( .A(A[4]), .Z(n13) );
  BUF_X1 U263 ( .A(n1), .Z(n28) );
endmodule


module adder_sub_N32 ( A, B, Ci, Cout, Sum );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Ci;
  output Cout;

  wire   [31:0] B_in;

  generic_xor_N32 xor_g ( .A(B), .B(Ci), .Y(B_in) );
  cla_adder_N32_0 add ( .A(A), .B(B_in), .Ci(Ci), .Cout(Cout), .Sum(Sum) );
endmodule


module mux_fwd_1 ( OP, alu_out, alu_wb_in, lmd_out, OPF, sel );
  input [31:0] OP;
  input [31:0] alu_out;
  input [31:0] alu_wb_in;
  input [31:0] lmd_out;
  output [31:0] OPF;
  input [2:0] sel;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164;

  BUF_X1 U1 ( .A(n5), .Z(n160) );
  BUF_X1 U2 ( .A(n5), .Z(n159) );
  BUF_X1 U3 ( .A(n7), .Z(n154) );
  BUF_X1 U4 ( .A(n7), .Z(n153) );
  BUF_X1 U5 ( .A(n6), .Z(n157) );
  BUF_X1 U6 ( .A(n6), .Z(n156) );
  BUF_X1 U7 ( .A(n5), .Z(n161) );
  BUF_X1 U8 ( .A(n7), .Z(n155) );
  BUF_X1 U9 ( .A(n6), .Z(n158) );
  NOR3_X1 U10 ( .A1(sel[1]), .A2(n164), .A3(n70), .ZN(n5) );
  INV_X1 U11 ( .A(sel[0]), .ZN(n70) );
  NOR3_X1 U12 ( .A1(sel[1]), .A2(n164), .A3(sel[0]), .ZN(n6) );
  BUF_X1 U13 ( .A(sel[2]), .Z(n164) );
  NOR2_X1 U14 ( .A1(n71), .A2(n164), .ZN(n7) );
  INV_X1 U15 ( .A(sel[1]), .ZN(n71) );
  BUF_X1 U16 ( .A(sel[2]), .Z(n163) );
  BUF_X1 U17 ( .A(sel[2]), .Z(n162) );
  NAND2_X1 U18 ( .A1(n10), .A2(n11), .ZN(OPF[7]) );
  AOI22_X1 U19 ( .A1(alu_wb_in[7]), .A2(n155), .B1(alu_out[7]), .B2(n162), 
        .ZN(n10) );
  AOI22_X1 U20 ( .A1(lmd_out[7]), .A2(n161), .B1(OP[7]), .B2(n158), .ZN(n11)
         );
  NAND2_X1 U21 ( .A1(n68), .A2(n69), .ZN(OPF[0]) );
  AOI22_X1 U22 ( .A1(alu_wb_in[0]), .A2(n153), .B1(alu_out[0]), .B2(n164), 
        .ZN(n68) );
  AOI22_X1 U23 ( .A1(lmd_out[0]), .A2(n159), .B1(OP[0]), .B2(n156), .ZN(n69)
         );
  NAND2_X1 U24 ( .A1(n46), .A2(n47), .ZN(OPF[1]) );
  AOI22_X1 U25 ( .A1(alu_wb_in[1]), .A2(n153), .B1(alu_out[1]), .B2(n163), 
        .ZN(n46) );
  AOI22_X1 U26 ( .A1(lmd_out[1]), .A2(n159), .B1(OP[1]), .B2(n156), .ZN(n47)
         );
  NAND2_X1 U27 ( .A1(n24), .A2(n25), .ZN(OPF[2]) );
  AOI22_X1 U28 ( .A1(alu_wb_in[2]), .A2(n154), .B1(alu_out[2]), .B2(n162), 
        .ZN(n24) );
  AOI22_X1 U29 ( .A1(lmd_out[2]), .A2(n160), .B1(OP[2]), .B2(n157), .ZN(n25)
         );
  NAND2_X1 U30 ( .A1(n18), .A2(n19), .ZN(OPF[3]) );
  AOI22_X1 U31 ( .A1(alu_wb_in[3]), .A2(n155), .B1(alu_out[3]), .B2(n162), 
        .ZN(n18) );
  AOI22_X1 U32 ( .A1(lmd_out[3]), .A2(n161), .B1(OP[3]), .B2(n158), .ZN(n19)
         );
  NAND2_X1 U33 ( .A1(n16), .A2(n17), .ZN(OPF[4]) );
  AOI22_X1 U34 ( .A1(alu_wb_in[4]), .A2(n155), .B1(alu_out[4]), .B2(n162), 
        .ZN(n16) );
  AOI22_X1 U35 ( .A1(lmd_out[4]), .A2(n161), .B1(OP[4]), .B2(n158), .ZN(n17)
         );
  NAND2_X1 U36 ( .A1(n14), .A2(n15), .ZN(OPF[5]) );
  AOI22_X1 U37 ( .A1(alu_wb_in[5]), .A2(n155), .B1(alu_out[5]), .B2(n162), 
        .ZN(n14) );
  AOI22_X1 U38 ( .A1(lmd_out[5]), .A2(n161), .B1(OP[5]), .B2(n158), .ZN(n15)
         );
  NAND2_X1 U39 ( .A1(n12), .A2(n13), .ZN(OPF[6]) );
  AOI22_X1 U40 ( .A1(alu_wb_in[6]), .A2(n155), .B1(alu_out[6]), .B2(n162), 
        .ZN(n12) );
  AOI22_X1 U41 ( .A1(lmd_out[6]), .A2(n161), .B1(OP[6]), .B2(n158), .ZN(n13)
         );
  NAND2_X1 U42 ( .A1(n8), .A2(n9), .ZN(OPF[8]) );
  AOI22_X1 U43 ( .A1(alu_wb_in[8]), .A2(n155), .B1(alu_out[8]), .B2(n162), 
        .ZN(n8) );
  AOI22_X1 U44 ( .A1(lmd_out[8]), .A2(n161), .B1(OP[8]), .B2(n158), .ZN(n9) );
  NAND2_X1 U45 ( .A1(n3), .A2(n4), .ZN(OPF[9]) );
  AOI22_X1 U46 ( .A1(alu_wb_in[9]), .A2(n155), .B1(n164), .B2(alu_out[9]), 
        .ZN(n3) );
  AOI22_X1 U47 ( .A1(lmd_out[9]), .A2(n161), .B1(OP[9]), .B2(n158), .ZN(n4) );
  NAND2_X1 U48 ( .A1(n66), .A2(n67), .ZN(OPF[10]) );
  AOI22_X1 U49 ( .A1(alu_wb_in[10]), .A2(n153), .B1(alu_out[10]), .B2(n164), 
        .ZN(n66) );
  AOI22_X1 U50 ( .A1(lmd_out[10]), .A2(n159), .B1(OP[10]), .B2(n156), .ZN(n67)
         );
  NAND2_X1 U51 ( .A1(n64), .A2(n65), .ZN(OPF[11]) );
  AOI22_X1 U52 ( .A1(alu_wb_in[11]), .A2(n153), .B1(alu_out[11]), .B2(n164), 
        .ZN(n64) );
  AOI22_X1 U53 ( .A1(lmd_out[11]), .A2(n159), .B1(OP[11]), .B2(n156), .ZN(n65)
         );
  NAND2_X1 U54 ( .A1(n62), .A2(n63), .ZN(OPF[12]) );
  AOI22_X1 U55 ( .A1(alu_wb_in[12]), .A2(n153), .B1(alu_out[12]), .B2(n164), 
        .ZN(n62) );
  AOI22_X1 U56 ( .A1(lmd_out[12]), .A2(n159), .B1(OP[12]), .B2(n156), .ZN(n63)
         );
  NAND2_X1 U57 ( .A1(n60), .A2(n61), .ZN(OPF[13]) );
  AOI22_X1 U58 ( .A1(alu_wb_in[13]), .A2(n153), .B1(alu_out[13]), .B2(n164), 
        .ZN(n60) );
  AOI22_X1 U59 ( .A1(lmd_out[13]), .A2(n159), .B1(OP[13]), .B2(n156), .ZN(n61)
         );
  NAND2_X1 U60 ( .A1(n58), .A2(n59), .ZN(OPF[14]) );
  AOI22_X1 U61 ( .A1(alu_wb_in[14]), .A2(n153), .B1(alu_out[14]), .B2(n164), 
        .ZN(n58) );
  AOI22_X1 U62 ( .A1(lmd_out[14]), .A2(n159), .B1(OP[14]), .B2(n156), .ZN(n59)
         );
  NAND2_X1 U63 ( .A1(n56), .A2(n57), .ZN(OPF[15]) );
  AOI22_X1 U64 ( .A1(alu_wb_in[15]), .A2(n153), .B1(alu_out[15]), .B2(n164), 
        .ZN(n56) );
  AOI22_X1 U65 ( .A1(lmd_out[15]), .A2(n159), .B1(OP[15]), .B2(n156), .ZN(n57)
         );
  NAND2_X1 U66 ( .A1(n20), .A2(n21), .ZN(OPF[31]) );
  AOI22_X1 U67 ( .A1(alu_wb_in[31]), .A2(n155), .B1(alu_out[31]), .B2(n162), 
        .ZN(n20) );
  AOI22_X1 U68 ( .A1(lmd_out[31]), .A2(n161), .B1(OP[31]), .B2(n158), .ZN(n21)
         );
  NAND2_X1 U69 ( .A1(n54), .A2(n55), .ZN(OPF[16]) );
  AOI22_X1 U70 ( .A1(alu_wb_in[16]), .A2(n153), .B1(alu_out[16]), .B2(n163), 
        .ZN(n54) );
  AOI22_X1 U71 ( .A1(lmd_out[16]), .A2(n159), .B1(OP[16]), .B2(n156), .ZN(n55)
         );
  NAND2_X1 U72 ( .A1(n52), .A2(n53), .ZN(OPF[17]) );
  AOI22_X1 U73 ( .A1(alu_wb_in[17]), .A2(n153), .B1(alu_out[17]), .B2(n163), 
        .ZN(n52) );
  AOI22_X1 U74 ( .A1(lmd_out[17]), .A2(n159), .B1(OP[17]), .B2(n156), .ZN(n53)
         );
  NAND2_X1 U75 ( .A1(n50), .A2(n51), .ZN(OPF[18]) );
  AOI22_X1 U76 ( .A1(alu_wb_in[18]), .A2(n153), .B1(alu_out[18]), .B2(n163), 
        .ZN(n50) );
  AOI22_X1 U77 ( .A1(lmd_out[18]), .A2(n159), .B1(OP[18]), .B2(n156), .ZN(n51)
         );
  NAND2_X1 U78 ( .A1(n48), .A2(n49), .ZN(OPF[19]) );
  AOI22_X1 U79 ( .A1(alu_wb_in[19]), .A2(n153), .B1(alu_out[19]), .B2(n163), 
        .ZN(n48) );
  AOI22_X1 U80 ( .A1(lmd_out[19]), .A2(n159), .B1(OP[19]), .B2(n156), .ZN(n49)
         );
  NAND2_X1 U81 ( .A1(n44), .A2(n45), .ZN(OPF[20]) );
  AOI22_X1 U82 ( .A1(alu_wb_in[20]), .A2(n154), .B1(alu_out[20]), .B2(n163), 
        .ZN(n44) );
  AOI22_X1 U83 ( .A1(lmd_out[20]), .A2(n160), .B1(OP[20]), .B2(n157), .ZN(n45)
         );
  NAND2_X1 U84 ( .A1(n42), .A2(n43), .ZN(OPF[21]) );
  AOI22_X1 U85 ( .A1(alu_wb_in[21]), .A2(n154), .B1(alu_out[21]), .B2(n163), 
        .ZN(n42) );
  AOI22_X1 U86 ( .A1(lmd_out[21]), .A2(n160), .B1(OP[21]), .B2(n157), .ZN(n43)
         );
  NAND2_X1 U87 ( .A1(n40), .A2(n41), .ZN(OPF[22]) );
  AOI22_X1 U88 ( .A1(alu_wb_in[22]), .A2(n154), .B1(alu_out[22]), .B2(n163), 
        .ZN(n40) );
  AOI22_X1 U89 ( .A1(lmd_out[22]), .A2(n160), .B1(OP[22]), .B2(n157), .ZN(n41)
         );
  NAND2_X1 U90 ( .A1(n38), .A2(n39), .ZN(OPF[23]) );
  AOI22_X1 U91 ( .A1(alu_wb_in[23]), .A2(n154), .B1(alu_out[23]), .B2(n163), 
        .ZN(n38) );
  AOI22_X1 U92 ( .A1(lmd_out[23]), .A2(n160), .B1(OP[23]), .B2(n157), .ZN(n39)
         );
  NAND2_X1 U93 ( .A1(n36), .A2(n37), .ZN(OPF[24]) );
  AOI22_X1 U94 ( .A1(alu_wb_in[24]), .A2(n154), .B1(alu_out[24]), .B2(n163), 
        .ZN(n36) );
  AOI22_X1 U95 ( .A1(lmd_out[24]), .A2(n160), .B1(OP[24]), .B2(n157), .ZN(n37)
         );
  NAND2_X1 U96 ( .A1(n34), .A2(n35), .ZN(OPF[25]) );
  AOI22_X1 U97 ( .A1(alu_wb_in[25]), .A2(n154), .B1(alu_out[25]), .B2(n163), 
        .ZN(n34) );
  AOI22_X1 U98 ( .A1(lmd_out[25]), .A2(n160), .B1(OP[25]), .B2(n157), .ZN(n35)
         );
  NAND2_X1 U99 ( .A1(n32), .A2(n33), .ZN(OPF[26]) );
  AOI22_X1 U100 ( .A1(alu_wb_in[26]), .A2(n154), .B1(alu_out[26]), .B2(n162), 
        .ZN(n32) );
  AOI22_X1 U101 ( .A1(lmd_out[26]), .A2(n160), .B1(OP[26]), .B2(n157), .ZN(n33) );
  NAND2_X1 U102 ( .A1(n30), .A2(n31), .ZN(OPF[27]) );
  AOI22_X1 U103 ( .A1(alu_wb_in[27]), .A2(n154), .B1(alu_out[27]), .B2(n162), 
        .ZN(n30) );
  AOI22_X1 U104 ( .A1(lmd_out[27]), .A2(n160), .B1(OP[27]), .B2(n157), .ZN(n31) );
  NAND2_X1 U105 ( .A1(n28), .A2(n29), .ZN(OPF[28]) );
  AOI22_X1 U106 ( .A1(alu_wb_in[28]), .A2(n154), .B1(alu_out[28]), .B2(n162), 
        .ZN(n28) );
  AOI22_X1 U107 ( .A1(lmd_out[28]), .A2(n160), .B1(OP[28]), .B2(n157), .ZN(n29) );
  NAND2_X1 U108 ( .A1(n26), .A2(n27), .ZN(OPF[29]) );
  AOI22_X1 U109 ( .A1(alu_wb_in[29]), .A2(n154), .B1(alu_out[29]), .B2(n162), 
        .ZN(n26) );
  AOI22_X1 U110 ( .A1(lmd_out[29]), .A2(n160), .B1(OP[29]), .B2(n157), .ZN(n27) );
  NAND2_X1 U111 ( .A1(n22), .A2(n23), .ZN(OPF[30]) );
  AOI22_X1 U112 ( .A1(alu_wb_in[30]), .A2(n154), .B1(alu_out[30]), .B2(n163), 
        .ZN(n22) );
  AOI22_X1 U113 ( .A1(lmd_out[30]), .A2(n160), .B1(OP[30]), .B2(n157), .ZN(n23) );
endmodule


module mux_fwd_0 ( OP, alu_out, alu_wb_in, lmd_out, OPF, sel );
  input [31:0] OP;
  input [31:0] alu_out;
  input [31:0] alu_wb_in;
  input [31:0] lmd_out;
  output [31:0] OPF;
  input [2:0] sel;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94;

  BUF_X1 U1 ( .A(n5), .Z(n89) );
  BUF_X1 U2 ( .A(n5), .Z(n90) );
  BUF_X1 U3 ( .A(n7), .Z(n83) );
  BUF_X1 U4 ( .A(n7), .Z(n84) );
  BUF_X1 U5 ( .A(n6), .Z(n86) );
  BUF_X1 U6 ( .A(n6), .Z(n87) );
  BUF_X1 U7 ( .A(n5), .Z(n91) );
  BUF_X1 U8 ( .A(n7), .Z(n85) );
  BUF_X1 U9 ( .A(n6), .Z(n88) );
  NOR3_X1 U10 ( .A1(sel[1]), .A2(n94), .A3(n70), .ZN(n5) );
  INV_X1 U11 ( .A(sel[0]), .ZN(n70) );
  NOR3_X1 U12 ( .A1(sel[1]), .A2(n94), .A3(sel[0]), .ZN(n6) );
  BUF_X1 U13 ( .A(sel[2]), .Z(n94) );
  NOR2_X1 U14 ( .A1(n71), .A2(n94), .ZN(n7) );
  INV_X1 U15 ( .A(sel[1]), .ZN(n71) );
  BUF_X1 U16 ( .A(sel[2]), .Z(n93) );
  BUF_X1 U17 ( .A(sel[2]), .Z(n92) );
  NAND2_X1 U18 ( .A1(n20), .A2(n21), .ZN(OPF[31]) );
  AOI22_X1 U19 ( .A1(alu_wb_in[31]), .A2(n85), .B1(alu_out[31]), .B2(n92), 
        .ZN(n20) );
  AOI22_X1 U20 ( .A1(lmd_out[31]), .A2(n91), .B1(OP[31]), .B2(n88), .ZN(n21)
         );
  NAND2_X1 U21 ( .A1(n10), .A2(n11), .ZN(OPF[7]) );
  AOI22_X1 U22 ( .A1(alu_wb_in[7]), .A2(n85), .B1(alu_out[7]), .B2(n92), .ZN(
        n10) );
  AOI22_X1 U23 ( .A1(lmd_out[7]), .A2(n91), .B1(OP[7]), .B2(n88), .ZN(n11) );
  NAND2_X1 U24 ( .A1(n68), .A2(n69), .ZN(OPF[0]) );
  AOI22_X1 U25 ( .A1(alu_wb_in[0]), .A2(n83), .B1(alu_out[0]), .B2(n94), .ZN(
        n68) );
  AOI22_X1 U26 ( .A1(lmd_out[0]), .A2(n89), .B1(OP[0]), .B2(n86), .ZN(n69) );
  NAND2_X1 U27 ( .A1(n46), .A2(n47), .ZN(OPF[1]) );
  AOI22_X1 U28 ( .A1(alu_wb_in[1]), .A2(n83), .B1(alu_out[1]), .B2(n93), .ZN(
        n46) );
  AOI22_X1 U29 ( .A1(lmd_out[1]), .A2(n89), .B1(OP[1]), .B2(n86), .ZN(n47) );
  NAND2_X1 U30 ( .A1(n24), .A2(n25), .ZN(OPF[2]) );
  AOI22_X1 U31 ( .A1(alu_wb_in[2]), .A2(n84), .B1(alu_out[2]), .B2(n92), .ZN(
        n24) );
  AOI22_X1 U32 ( .A1(lmd_out[2]), .A2(n90), .B1(OP[2]), .B2(n87), .ZN(n25) );
  NAND2_X1 U33 ( .A1(n18), .A2(n19), .ZN(OPF[3]) );
  AOI22_X1 U34 ( .A1(alu_wb_in[3]), .A2(n85), .B1(alu_out[3]), .B2(n92), .ZN(
        n18) );
  AOI22_X1 U35 ( .A1(lmd_out[3]), .A2(n91), .B1(OP[3]), .B2(n88), .ZN(n19) );
  NAND2_X1 U36 ( .A1(n16), .A2(n17), .ZN(OPF[4]) );
  AOI22_X1 U37 ( .A1(alu_wb_in[4]), .A2(n85), .B1(alu_out[4]), .B2(n92), .ZN(
        n16) );
  AOI22_X1 U38 ( .A1(lmd_out[4]), .A2(n91), .B1(OP[4]), .B2(n88), .ZN(n17) );
  NAND2_X1 U39 ( .A1(n14), .A2(n15), .ZN(OPF[5]) );
  AOI22_X1 U40 ( .A1(alu_wb_in[5]), .A2(n85), .B1(alu_out[5]), .B2(n92), .ZN(
        n14) );
  AOI22_X1 U41 ( .A1(lmd_out[5]), .A2(n91), .B1(OP[5]), .B2(n88), .ZN(n15) );
  NAND2_X1 U42 ( .A1(n12), .A2(n13), .ZN(OPF[6]) );
  AOI22_X1 U43 ( .A1(alu_wb_in[6]), .A2(n85), .B1(alu_out[6]), .B2(n92), .ZN(
        n12) );
  AOI22_X1 U44 ( .A1(lmd_out[6]), .A2(n91), .B1(OP[6]), .B2(n88), .ZN(n13) );
  NAND2_X1 U45 ( .A1(n8), .A2(n9), .ZN(OPF[8]) );
  AOI22_X1 U46 ( .A1(alu_wb_in[8]), .A2(n85), .B1(alu_out[8]), .B2(n92), .ZN(
        n8) );
  AOI22_X1 U47 ( .A1(lmd_out[8]), .A2(n91), .B1(OP[8]), .B2(n88), .ZN(n9) );
  NAND2_X1 U48 ( .A1(n3), .A2(n4), .ZN(OPF[9]) );
  AOI22_X1 U49 ( .A1(alu_wb_in[9]), .A2(n85), .B1(n94), .B2(alu_out[9]), .ZN(
        n3) );
  AOI22_X1 U50 ( .A1(lmd_out[9]), .A2(n91), .B1(OP[9]), .B2(n88), .ZN(n4) );
  NAND2_X1 U51 ( .A1(n66), .A2(n67), .ZN(OPF[10]) );
  AOI22_X1 U52 ( .A1(alu_wb_in[10]), .A2(n83), .B1(alu_out[10]), .B2(n94), 
        .ZN(n66) );
  AOI22_X1 U53 ( .A1(lmd_out[10]), .A2(n89), .B1(OP[10]), .B2(n86), .ZN(n67)
         );
  NAND2_X1 U54 ( .A1(n64), .A2(n65), .ZN(OPF[11]) );
  AOI22_X1 U55 ( .A1(alu_wb_in[11]), .A2(n83), .B1(alu_out[11]), .B2(n94), 
        .ZN(n64) );
  AOI22_X1 U56 ( .A1(lmd_out[11]), .A2(n89), .B1(OP[11]), .B2(n86), .ZN(n65)
         );
  NAND2_X1 U57 ( .A1(n62), .A2(n63), .ZN(OPF[12]) );
  AOI22_X1 U58 ( .A1(alu_wb_in[12]), .A2(n83), .B1(alu_out[12]), .B2(n94), 
        .ZN(n62) );
  AOI22_X1 U59 ( .A1(lmd_out[12]), .A2(n89), .B1(OP[12]), .B2(n86), .ZN(n63)
         );
  NAND2_X1 U60 ( .A1(n60), .A2(n61), .ZN(OPF[13]) );
  AOI22_X1 U61 ( .A1(alu_wb_in[13]), .A2(n83), .B1(alu_out[13]), .B2(n94), 
        .ZN(n60) );
  AOI22_X1 U62 ( .A1(lmd_out[13]), .A2(n89), .B1(OP[13]), .B2(n86), .ZN(n61)
         );
  NAND2_X1 U63 ( .A1(n58), .A2(n59), .ZN(OPF[14]) );
  AOI22_X1 U64 ( .A1(alu_wb_in[14]), .A2(n83), .B1(alu_out[14]), .B2(n94), 
        .ZN(n58) );
  AOI22_X1 U65 ( .A1(lmd_out[14]), .A2(n89), .B1(OP[14]), .B2(n86), .ZN(n59)
         );
  NAND2_X1 U66 ( .A1(n56), .A2(n57), .ZN(OPF[15]) );
  AOI22_X1 U67 ( .A1(alu_wb_in[15]), .A2(n83), .B1(alu_out[15]), .B2(n94), 
        .ZN(n56) );
  AOI22_X1 U68 ( .A1(lmd_out[15]), .A2(n89), .B1(OP[15]), .B2(n86), .ZN(n57)
         );
  NAND2_X1 U69 ( .A1(n54), .A2(n55), .ZN(OPF[16]) );
  AOI22_X1 U70 ( .A1(alu_wb_in[16]), .A2(n83), .B1(alu_out[16]), .B2(n93), 
        .ZN(n54) );
  AOI22_X1 U71 ( .A1(lmd_out[16]), .A2(n89), .B1(OP[16]), .B2(n86), .ZN(n55)
         );
  NAND2_X1 U72 ( .A1(n52), .A2(n53), .ZN(OPF[17]) );
  AOI22_X1 U73 ( .A1(alu_wb_in[17]), .A2(n83), .B1(alu_out[17]), .B2(n93), 
        .ZN(n52) );
  AOI22_X1 U74 ( .A1(lmd_out[17]), .A2(n89), .B1(OP[17]), .B2(n86), .ZN(n53)
         );
  NAND2_X1 U75 ( .A1(n50), .A2(n51), .ZN(OPF[18]) );
  AOI22_X1 U76 ( .A1(alu_wb_in[18]), .A2(n83), .B1(alu_out[18]), .B2(n93), 
        .ZN(n50) );
  AOI22_X1 U77 ( .A1(lmd_out[18]), .A2(n89), .B1(OP[18]), .B2(n86), .ZN(n51)
         );
  NAND2_X1 U78 ( .A1(n48), .A2(n49), .ZN(OPF[19]) );
  AOI22_X1 U79 ( .A1(alu_wb_in[19]), .A2(n83), .B1(alu_out[19]), .B2(n93), 
        .ZN(n48) );
  AOI22_X1 U80 ( .A1(lmd_out[19]), .A2(n89), .B1(OP[19]), .B2(n86), .ZN(n49)
         );
  NAND2_X1 U81 ( .A1(n44), .A2(n45), .ZN(OPF[20]) );
  AOI22_X1 U82 ( .A1(alu_wb_in[20]), .A2(n84), .B1(alu_out[20]), .B2(n93), 
        .ZN(n44) );
  AOI22_X1 U83 ( .A1(lmd_out[20]), .A2(n90), .B1(OP[20]), .B2(n87), .ZN(n45)
         );
  NAND2_X1 U84 ( .A1(n42), .A2(n43), .ZN(OPF[21]) );
  AOI22_X1 U85 ( .A1(alu_wb_in[21]), .A2(n84), .B1(alu_out[21]), .B2(n93), 
        .ZN(n42) );
  AOI22_X1 U86 ( .A1(lmd_out[21]), .A2(n90), .B1(OP[21]), .B2(n87), .ZN(n43)
         );
  NAND2_X1 U87 ( .A1(n40), .A2(n41), .ZN(OPF[22]) );
  AOI22_X1 U88 ( .A1(alu_wb_in[22]), .A2(n84), .B1(alu_out[22]), .B2(n93), 
        .ZN(n40) );
  AOI22_X1 U89 ( .A1(lmd_out[22]), .A2(n90), .B1(OP[22]), .B2(n87), .ZN(n41)
         );
  NAND2_X1 U90 ( .A1(n38), .A2(n39), .ZN(OPF[23]) );
  AOI22_X1 U91 ( .A1(alu_wb_in[23]), .A2(n84), .B1(alu_out[23]), .B2(n93), 
        .ZN(n38) );
  AOI22_X1 U92 ( .A1(lmd_out[23]), .A2(n90), .B1(OP[23]), .B2(n87), .ZN(n39)
         );
  NAND2_X1 U93 ( .A1(n36), .A2(n37), .ZN(OPF[24]) );
  AOI22_X1 U94 ( .A1(alu_wb_in[24]), .A2(n84), .B1(alu_out[24]), .B2(n93), 
        .ZN(n36) );
  AOI22_X1 U95 ( .A1(lmd_out[24]), .A2(n90), .B1(OP[24]), .B2(n87), .ZN(n37)
         );
  NAND2_X1 U96 ( .A1(n34), .A2(n35), .ZN(OPF[25]) );
  AOI22_X1 U97 ( .A1(alu_wb_in[25]), .A2(n84), .B1(alu_out[25]), .B2(n93), 
        .ZN(n34) );
  AOI22_X1 U98 ( .A1(lmd_out[25]), .A2(n90), .B1(OP[25]), .B2(n87), .ZN(n35)
         );
  NAND2_X1 U99 ( .A1(n32), .A2(n33), .ZN(OPF[26]) );
  AOI22_X1 U100 ( .A1(alu_wb_in[26]), .A2(n84), .B1(alu_out[26]), .B2(n92), 
        .ZN(n32) );
  AOI22_X1 U101 ( .A1(lmd_out[26]), .A2(n90), .B1(OP[26]), .B2(n87), .ZN(n33)
         );
  NAND2_X1 U102 ( .A1(n30), .A2(n31), .ZN(OPF[27]) );
  AOI22_X1 U103 ( .A1(alu_wb_in[27]), .A2(n84), .B1(alu_out[27]), .B2(n92), 
        .ZN(n30) );
  AOI22_X1 U104 ( .A1(lmd_out[27]), .A2(n90), .B1(OP[27]), .B2(n87), .ZN(n31)
         );
  NAND2_X1 U105 ( .A1(n28), .A2(n29), .ZN(OPF[28]) );
  AOI22_X1 U106 ( .A1(alu_wb_in[28]), .A2(n84), .B1(alu_out[28]), .B2(n92), 
        .ZN(n28) );
  AOI22_X1 U107 ( .A1(lmd_out[28]), .A2(n90), .B1(OP[28]), .B2(n87), .ZN(n29)
         );
  NAND2_X1 U108 ( .A1(n26), .A2(n27), .ZN(OPF[29]) );
  AOI22_X1 U109 ( .A1(alu_wb_in[29]), .A2(n84), .B1(alu_out[29]), .B2(n92), 
        .ZN(n26) );
  AOI22_X1 U110 ( .A1(lmd_out[29]), .A2(n90), .B1(OP[29]), .B2(n87), .ZN(n27)
         );
  NAND2_X1 U111 ( .A1(n22), .A2(n23), .ZN(OPF[30]) );
  AOI22_X1 U112 ( .A1(alu_wb_in[30]), .A2(n84), .B1(alu_out[30]), .B2(n93), 
        .ZN(n22) );
  AOI22_X1 U113 ( .A1(lmd_out[30]), .A2(n90), .B1(OP[30]), .B2(n87), .ZN(n23)
         );
endmodule


module counter ( clk, rst, tc );
  input clk, rst;
  output tc;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N125, N127, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n68, net227481,
         net227482, net227483, net227484, net227485, net227486, net227487,
         net227488, net227489, net227490, net227491, net227492, net227493,
         net227494, net227495, net227496, net227505, net227506, net227507,
         net227508, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n119, n120, n121, n122, n123;
  wire   [30:0] i;
  assign n68 = rst;

  DFFR_X1 \i_reg[0]  ( .D(n118), .CK(clk), .RN(n121), .Q(i[0]) );
  DFFR_X1 \i_reg[30]  ( .D(n117), .CK(clk), .RN(n122), .Q(i[30]) );
  DFFR_X1 \i_reg[28]  ( .D(n116), .CK(clk), .RN(n122), .Q(i[28]) );
  DFFR_X1 \i_reg[26]  ( .D(n115), .CK(clk), .RN(n122), .Q(i[26]), .QN(
        net227508) );
  DFFR_X1 \i_reg[24]  ( .D(n114), .CK(clk), .RN(n122), .Q(i[24]), .QN(
        net227507) );
  DFFR_X1 \i_reg[22]  ( .D(n113), .CK(clk), .RN(n122), .Q(i[22]), .QN(
        net227506) );
  DFFR_X1 \i_reg[20]  ( .D(n112), .CK(clk), .RN(n122), .Q(i[20]), .QN(
        net227505) );
  DFFR_X1 \i_reg[18]  ( .D(n111), .CK(clk), .RN(n121), .Q(i[18]) );
  DFFR_X1 \i_reg[16]  ( .D(n110), .CK(clk), .RN(n121), .Q(i[16]) );
  DFFR_X1 \i_reg[14]  ( .D(n109), .CK(clk), .RN(n121), .Q(i[14]) );
  DFFR_X1 \i_reg[12]  ( .D(n108), .CK(clk), .RN(n121), .Q(i[12]) );
  DFFR_X1 \i_reg[10]  ( .D(n107), .CK(clk), .RN(n121), .Q(i[10]) );
  DFFR_X1 \i_reg[8]  ( .D(n106), .CK(clk), .RN(n122), .Q(i[8]) );
  DFFR_X1 \i_reg[6]  ( .D(n105), .CK(clk), .RN(n123), .Q(i[6]) );
  DFFR_X1 \i_reg[4]  ( .D(n104), .CK(clk), .RN(n123), .Q(i[4]) );
  DFFR_X1 \i_reg[2]  ( .D(n103), .CK(clk), .RN(n122), .Q(i[2]), .QN(net227496)
         );
  DFFS_X1 \i_reg[1]  ( .D(n102), .CK(clk), .SN(n123), .Q(i[1]), .QN(net227495)
         );
  DFFR_X1 \i_reg[3]  ( .D(n101), .CK(clk), .RN(n123), .Q(i[3]), .QN(net227494)
         );
  DFFR_X1 \i_reg[5]  ( .D(n100), .CK(clk), .RN(n123), .Q(i[5]), .QN(net227493)
         );
  DFFR_X1 \i_reg[7]  ( .D(n99), .CK(clk), .RN(n123), .Q(i[7]), .QN(net227492)
         );
  DFFR_X1 \i_reg[9]  ( .D(n98), .CK(clk), .RN(n123), .Q(i[9]), .QN(net227491)
         );
  DFFR_X1 \i_reg[11]  ( .D(n97), .CK(clk), .RN(n122), .Q(i[11]), .QN(net227490) );
  DFFR_X1 \i_reg[13]  ( .D(n96), .CK(clk), .RN(n122), .Q(i[13]), .QN(net227489) );
  DFFR_X1 \i_reg[15]  ( .D(n95), .CK(clk), .RN(n122), .Q(i[15]), .QN(net227488) );
  DFFR_X1 \i_reg[17]  ( .D(n94), .CK(clk), .RN(n121), .Q(i[17]), .QN(net227487) );
  DFFR_X1 \i_reg[19]  ( .D(n93), .CK(clk), .RN(n122), .Q(i[19]), .QN(net227486) );
  DFFR_X1 \i_reg[21]  ( .D(n92), .CK(clk), .RN(n121), .Q(i[21]), .QN(net227485) );
  DFFR_X1 \i_reg[23]  ( .D(n91), .CK(clk), .RN(n121), .Q(i[23]), .QN(net227484) );
  DFFR_X1 \i_reg[25]  ( .D(n90), .CK(clk), .RN(n121), .Q(i[25]), .QN(net227483) );
  DFFR_X1 \i_reg[27]  ( .D(n89), .CK(clk), .RN(n121), .Q(i[27]), .QN(net227482) );
  DFFR_X1 \i_reg[29]  ( .D(n88), .CK(clk), .RN(n121), .Q(i[29]), .QN(net227481) );
  DFFS_X1 tc_reg ( .D(N125), .CK(clk), .SN(n123), .Q(tc) );
  counter_DW01_dec_0 sub_19 ( .A(i), .SUM({N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N127, N4}) );
  OR3_X1 U3 ( .A1(n77), .A2(n78), .A3(n76), .ZN(n84) );
  NOR2_X1 U4 ( .A1(n120), .A2(n39), .ZN(n93) );
  NOR2_X1 U5 ( .A1(n120), .A2(n37), .ZN(n95) );
  NOR2_X1 U6 ( .A1(n119), .A2(n47), .ZN(n116) );
  INV_X1 U7 ( .A(N31), .ZN(n47) );
  NOR2_X1 U8 ( .A1(n119), .A2(n41), .ZN(n91) );
  INV_X1 U9 ( .A(N26), .ZN(n41) );
  NOR2_X1 U10 ( .A1(n119), .A2(n52), .ZN(n111) );
  NOR2_X1 U11 ( .A1(n119), .A2(n51), .ZN(n112) );
  NOR2_X1 U12 ( .A1(n119), .A2(n50), .ZN(n113) );
  INV_X1 U13 ( .A(N25), .ZN(n50) );
  NOR2_X1 U14 ( .A1(n119), .A2(n48), .ZN(n115) );
  INV_X1 U15 ( .A(N29), .ZN(n48) );
  NOR2_X1 U16 ( .A1(n86), .A2(n57), .ZN(n106) );
  NOR2_X1 U17 ( .A1(n86), .A2(n56), .ZN(n107) );
  INV_X1 U18 ( .A(N13), .ZN(n56) );
  NOR4_X1 U19 ( .A1(N15), .A2(N14), .A3(N13), .A4(N127), .ZN(n79) );
  NOR4_X1 U20 ( .A1(N9), .A2(N8), .A3(N7), .A4(N6), .ZN(n83) );
  NOR4_X1 U21 ( .A1(N31), .A2(N30), .A3(N29), .A4(N28), .ZN(n81) );
  NOR4_X1 U22 ( .A1(N27), .A2(N26), .A3(N25), .A4(N24), .ZN(n80) );
  OR2_X1 U23 ( .A1(N5), .A2(N4), .ZN(n85) );
  INV_X1 U24 ( .A(N21), .ZN(n52) );
  NOR2_X1 U25 ( .A1(n120), .A2(n40), .ZN(n92) );
  INV_X1 U26 ( .A(N24), .ZN(n40) );
  NOR2_X1 U27 ( .A1(n120), .A2(n38), .ZN(n94) );
  NOR2_X1 U28 ( .A1(n120), .A2(n36), .ZN(n96) );
  NOR2_X1 U29 ( .A1(n120), .A2(n35), .ZN(n97) );
  INV_X1 U30 ( .A(N14), .ZN(n35) );
  NOR2_X1 U31 ( .A1(n120), .A2(n34), .ZN(n98) );
  NOR2_X1 U32 ( .A1(n120), .A2(n33), .ZN(n99) );
  NOR2_X1 U33 ( .A1(n119), .A2(n44), .ZN(n88) );
  INV_X1 U34 ( .A(N32), .ZN(n44) );
  NOR2_X1 U35 ( .A1(n119), .A2(n43), .ZN(n89) );
  INV_X1 U36 ( .A(N30), .ZN(n43) );
  NOR2_X1 U37 ( .A1(n119), .A2(n46), .ZN(n117) );
  NOR2_X1 U38 ( .A1(n119), .A2(n42), .ZN(n90) );
  INV_X1 U39 ( .A(N28), .ZN(n42) );
  NOR2_X1 U40 ( .A1(n119), .A2(n49), .ZN(n114) );
  INV_X1 U41 ( .A(N27), .ZN(n49) );
  NOR2_X1 U42 ( .A1(n86), .A2(n55), .ZN(n108) );
  INV_X1 U43 ( .A(N15), .ZN(n55) );
  NOR2_X1 U44 ( .A1(n86), .A2(n54), .ZN(n109) );
  NOR2_X1 U45 ( .A1(n86), .A2(n53), .ZN(n110) );
  INV_X1 U46 ( .A(N18), .ZN(n37) );
  INV_X1 U47 ( .A(N22), .ZN(n39) );
  INV_X1 U48 ( .A(N11), .ZN(n57) );
  INV_X1 U49 ( .A(N23), .ZN(n51) );
  BUF_X1 U50 ( .A(n32), .Z(n119) );
  BUF_X1 U51 ( .A(n32), .Z(n86) );
  BUF_X1 U52 ( .A(n32), .Z(n120) );
  NOR2_X1 U53 ( .A1(n86), .A2(n61), .ZN(n102) );
  INV_X1 U54 ( .A(N127), .ZN(n61) );
  NOR2_X1 U55 ( .A1(n119), .A2(n45), .ZN(n118) );
  INV_X1 U56 ( .A(N4), .ZN(n45) );
  NOR2_X1 U57 ( .A1(n86), .A2(n63), .ZN(n100) );
  INV_X1 U58 ( .A(N8), .ZN(n63) );
  NOR2_X1 U59 ( .A1(n86), .A2(n62), .ZN(n101) );
  INV_X1 U60 ( .A(N6), .ZN(n62) );
  NOR2_X1 U61 ( .A1(n86), .A2(n60), .ZN(n103) );
  INV_X1 U62 ( .A(N5), .ZN(n60) );
  NOR2_X1 U63 ( .A1(n86), .A2(n59), .ZN(n104) );
  INV_X1 U64 ( .A(N7), .ZN(n59) );
  NOR2_X1 U65 ( .A1(n86), .A2(n58), .ZN(n105) );
  INV_X1 U66 ( .A(N9), .ZN(n58) );
  BUF_X1 U67 ( .A(n68), .Z(n122) );
  BUF_X1 U68 ( .A(n68), .Z(n121) );
  BUF_X1 U69 ( .A(n68), .Z(n123) );
  INV_X1 U70 ( .A(N19), .ZN(n53) );
  INV_X1 U71 ( .A(N20), .ZN(n38) );
  INV_X1 U72 ( .A(N17), .ZN(n54) );
  INV_X1 U73 ( .A(N10), .ZN(n33) );
  INV_X1 U74 ( .A(N12), .ZN(n34) );
  INV_X1 U75 ( .A(N16), .ZN(n36) );
  NOR4_X1 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(n69) );
  NAND4_X1 U77 ( .A1(net227484), .A2(net227483), .A3(net227482), .A4(net227481), .ZN(n70) );
  NAND4_X1 U78 ( .A1(net227488), .A2(net227487), .A3(net227486), .A4(net227485), .ZN(n71) );
  NAND4_X1 U79 ( .A1(net227492), .A2(net227491), .A3(net227490), .A4(net227489), .ZN(n72) );
  NAND4_X1 U80 ( .A1(net227496), .A2(net227495), .A3(net227494), .A4(net227493), .ZN(n73) );
  NAND4_X1 U81 ( .A1(net227508), .A2(net227507), .A3(net227506), .A4(net227505), .ZN(n74) );
  AND4_X1 U82 ( .A1(n65), .A2(n66), .A3(n67), .A4(n69), .ZN(n32) );
  NOR4_X1 U83 ( .A1(i[12]), .A2(i[14]), .A3(i[16]), .A4(i[18]), .ZN(n65) );
  NOR4_X1 U84 ( .A1(i[4]), .A2(i[6]), .A3(i[8]), .A4(i[10]), .ZN(n66) );
  NOR3_X1 U85 ( .A1(N33), .A2(N32), .A3(n85), .ZN(n82) );
  NOR2_X1 U86 ( .A1(n75), .A2(n84), .ZN(n64) );
  NAND4_X1 U87 ( .A1(n57), .A2(n34), .A3(n33), .A4(n79), .ZN(n76) );
  NAND4_X1 U88 ( .A1(n38), .A2(n52), .A3(n39), .A4(n51), .ZN(n77) );
  NAND4_X1 U89 ( .A1(n36), .A2(n54), .A3(n37), .A4(n53), .ZN(n78) );
  NOR2_X1 U90 ( .A1(n64), .A2(n86), .ZN(N125) );
  NOR4_X1 U91 ( .A1(n74), .A2(i[0]), .A3(i[28]), .A4(i[30]), .ZN(n67) );
  INV_X1 U92 ( .A(N33), .ZN(n46) );
  NAND4_X1 U93 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(n75) );
endmodule


module reg_N2_0 ( clk, rst, d_in, d_out );
  input [1:0] d_in;
  output [1:0] d_out;
  input clk, rst;
  wire   N2, N3;

  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U4 ( .A1(rst), .A2(d_in[1]), .ZN(N3) );
endmodule


module mux_pc ( A, B, C, D, E, F, sel, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [2:0] sel;
  output [31:0] Y;
  wire   n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n23, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169;
  tri   [31:0] Y;

  TBUF_X1 \Y_tri[12]  ( .A(n126), .EN(n169), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n125), .EN(n169), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n124), .EN(n169), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n123), .EN(n169), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n122), .EN(n169), .Z(Y[16]) );
  TBUF_X1 \Y_tri[18]  ( .A(n120), .EN(n169), .Z(Y[18]) );
  TBUF_X1 \Y_tri[21]  ( .A(n117), .EN(n169), .Z(Y[21]) );
  TBUF_X1 \Y_tri[23]  ( .A(n115), .EN(n169), .Z(Y[23]) );
  TBUF_X1 \Y_tri[3]  ( .A(n136), .EN(n167), .Z(Y[3]) );
  TBUF_X1 \Y_tri[5]  ( .A(n134), .EN(n167), .Z(Y[5]) );
  TBUF_X1 \Y_tri[7]  ( .A(n132), .EN(n167), .Z(Y[7]) );
  TBUF_X1 \Y_tri[9]  ( .A(n129), .EN(n167), .Z(Y[9]) );
  TBUF_X1 \Y_tri[25]  ( .A(n113), .EN(n167), .Z(Y[25]) );
  TBUF_X1 \Y_tri[27]  ( .A(n111), .EN(n167), .Z(Y[27]) );
  TBUF_X1 \Y_tri[2]  ( .A(n137), .EN(n167), .Z(Y[2]) );
  TBUF_X1 \Y_tri[4]  ( .A(n135), .EN(n167), .Z(Y[4]) );
  TBUF_X1 \Y_tri[6]  ( .A(n133), .EN(n167), .Z(Y[6]) );
  TBUF_X1 \Y_tri[8]  ( .A(n131), .EN(n168), .Z(Y[8]) );
  TBUF_X1 \Y_tri[17]  ( .A(n121), .EN(n168), .Z(Y[17]) );
  TBUF_X1 \Y_tri[19]  ( .A(n119), .EN(n168), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n118), .EN(n168), .Z(Y[20]) );
  TBUF_X1 \Y_tri[22]  ( .A(n116), .EN(n168), .Z(Y[22]) );
  TBUF_X1 \Y_tri[24]  ( .A(n114), .EN(n168), .Z(Y[24]) );
  TBUF_X1 \Y_tri[26]  ( .A(n112), .EN(n168), .Z(Y[26]) );
  TBUF_X1 \Y_tri[28]  ( .A(n110), .EN(n168), .Z(Y[28]) );
  TBUF_X1 \Y_tri[0]  ( .A(n139), .EN(n168), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n138), .EN(n168), .Z(Y[1]) );
  TBUF_X1 \Y_tri[10]  ( .A(n128), .EN(n168), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n127), .EN(n168), .Z(Y[11]) );
  TBUF_X1 \Y_tri[31]  ( .A(n107), .EN(n167), .Z(Y[31]) );
  TBUF_X1 \Y_tri[29]  ( .A(n109), .EN(n167), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n108), .EN(n167), .Z(Y[30]) );
  BUF_X1 U1 ( .A(n23), .Z(n168) );
  BUF_X1 U2 ( .A(n23), .Z(n167) );
  BUF_X1 U3 ( .A(n9), .Z(n162) );
  BUF_X1 U4 ( .A(n9), .Z(n161) );
  BUF_X1 U5 ( .A(n10), .Z(n159) );
  BUF_X1 U6 ( .A(n10), .Z(n158) );
  BUF_X1 U7 ( .A(n9), .Z(n163) );
  BUF_X1 U8 ( .A(n10), .Z(n160) );
  BUF_X1 U9 ( .A(n23), .Z(n169) );
  BUF_X1 U10 ( .A(n12), .Z(n153) );
  BUF_X1 U11 ( .A(n12), .Z(n152) );
  NOR2_X1 U12 ( .A1(n77), .A2(n4), .ZN(n10) );
  NOR2_X1 U13 ( .A1(n77), .A2(n5), .ZN(n9) );
  BUF_X1 U14 ( .A(n13), .Z(n150) );
  BUF_X1 U15 ( .A(n13), .Z(n149) );
  BUF_X1 U16 ( .A(n11), .Z(n156) );
  BUF_X1 U17 ( .A(n8), .Z(n165) );
  BUF_X1 U18 ( .A(n11), .Z(n155) );
  BUF_X1 U19 ( .A(n8), .Z(n164) );
  BUF_X1 U20 ( .A(n12), .Z(n154) );
  BUF_X1 U21 ( .A(n13), .Z(n151) );
  BUF_X1 U22 ( .A(n11), .Z(n157) );
  BUF_X1 U23 ( .A(n8), .Z(n166) );
  NOR2_X1 U24 ( .A1(n4), .A2(n5), .ZN(n23) );
  NOR3_X1 U25 ( .A1(sel[1]), .A2(sel[2]), .A3(n77), .ZN(n13) );
  NOR3_X1 U26 ( .A1(sel[1]), .A2(sel[2]), .A3(sel[0]), .ZN(n12) );
  NOR2_X1 U27 ( .A1(n5), .A2(sel[0]), .ZN(n11) );
  NOR2_X1 U28 ( .A1(n4), .A2(sel[0]), .ZN(n8) );
  INV_X1 U29 ( .A(sel[1]), .ZN(n5) );
  INV_X1 U30 ( .A(sel[0]), .ZN(n77) );
  INV_X1 U31 ( .A(sel[2]), .ZN(n4) );
  NAND2_X1 U32 ( .A1(n73), .A2(n74), .ZN(n108) );
  AOI222_X1 U33 ( .A1(E[30]), .A2(n164), .B1(D[30]), .B2(n161), .C1(F[30]), 
        .C2(n158), .ZN(n74) );
  AOI222_X1 U34 ( .A1(C[30]), .A2(n155), .B1(A[30]), .B2(n152), .C1(B[30]), 
        .C2(n149), .ZN(n73) );
  NAND2_X1 U35 ( .A1(n71), .A2(n72), .ZN(n109) );
  AOI222_X1 U36 ( .A1(E[29]), .A2(n164), .B1(D[29]), .B2(n161), .C1(F[29]), 
        .C2(n158), .ZN(n72) );
  AOI222_X1 U37 ( .A1(C[29]), .A2(n155), .B1(A[29]), .B2(n152), .C1(B[29]), 
        .C2(n149), .ZN(n71) );
  NAND2_X1 U38 ( .A1(n59), .A2(n60), .ZN(n115) );
  AOI222_X1 U39 ( .A1(E[23]), .A2(n164), .B1(D[23]), .B2(n161), .C1(F[23]), 
        .C2(n158), .ZN(n60) );
  AOI222_X1 U40 ( .A1(C[23]), .A2(n155), .B1(A[23]), .B2(n152), .C1(B[23]), 
        .C2(n149), .ZN(n59) );
  NAND2_X1 U41 ( .A1(n69), .A2(n70), .ZN(n110) );
  AOI222_X1 U42 ( .A1(E[28]), .A2(n164), .B1(D[28]), .B2(n161), .C1(F[28]), 
        .C2(n158), .ZN(n70) );
  AOI222_X1 U43 ( .A1(C[28]), .A2(n155), .B1(A[28]), .B2(n152), .C1(B[28]), 
        .C2(n149), .ZN(n69) );
  NAND2_X1 U44 ( .A1(n65), .A2(n66), .ZN(n112) );
  AOI222_X1 U45 ( .A1(E[26]), .A2(n164), .B1(D[26]), .B2(n161), .C1(F[26]), 
        .C2(n158), .ZN(n66) );
  AOI222_X1 U46 ( .A1(C[26]), .A2(n155), .B1(A[26]), .B2(n152), .C1(B[26]), 
        .C2(n149), .ZN(n65) );
  NAND2_X1 U47 ( .A1(n61), .A2(n62), .ZN(n114) );
  AOI222_X1 U48 ( .A1(E[24]), .A2(n164), .B1(D[24]), .B2(n161), .C1(F[24]), 
        .C2(n158), .ZN(n62) );
  AOI222_X1 U49 ( .A1(C[24]), .A2(n155), .B1(A[24]), .B2(n152), .C1(B[24]), 
        .C2(n149), .ZN(n61) );
  NAND2_X1 U50 ( .A1(n67), .A2(n68), .ZN(n111) );
  AOI222_X1 U51 ( .A1(E[27]), .A2(n164), .B1(D[27]), .B2(n161), .C1(F[27]), 
        .C2(n158), .ZN(n68) );
  AOI222_X1 U52 ( .A1(C[27]), .A2(n155), .B1(A[27]), .B2(n152), .C1(B[27]), 
        .C2(n149), .ZN(n67) );
  NAND2_X1 U53 ( .A1(n63), .A2(n64), .ZN(n113) );
  AOI222_X1 U54 ( .A1(E[25]), .A2(n164), .B1(D[25]), .B2(n161), .C1(F[25]), 
        .C2(n158), .ZN(n64) );
  AOI222_X1 U55 ( .A1(C[25]), .A2(n155), .B1(A[25]), .B2(n152), .C1(B[25]), 
        .C2(n149), .ZN(n63) );
  NAND2_X1 U56 ( .A1(n14), .A2(n15), .ZN(n138) );
  AOI222_X1 U57 ( .A1(E[1]), .A2(n166), .B1(D[1]), .B2(n163), .C1(F[1]), .C2(
        n160), .ZN(n15) );
  AOI222_X1 U58 ( .A1(C[1]), .A2(n157), .B1(A[1]), .B2(n154), .C1(B[1]), .C2(
        n151), .ZN(n14) );
  NAND2_X1 U59 ( .A1(n6), .A2(n7), .ZN(n139) );
  AOI222_X1 U60 ( .A1(E[0]), .A2(n166), .B1(D[0]), .B2(n163), .C1(F[0]), .C2(
        n160), .ZN(n7) );
  AOI222_X1 U61 ( .A1(C[0]), .A2(n157), .B1(A[0]), .B2(n154), .C1(B[0]), .C2(
        n151), .ZN(n6) );
  NAND2_X1 U62 ( .A1(n25), .A2(n26), .ZN(n133) );
  AOI222_X1 U63 ( .A1(E[6]), .A2(n166), .B1(D[6]), .B2(n163), .C1(F[6]), .C2(
        n160), .ZN(n26) );
  AOI222_X1 U64 ( .A1(C[6]), .A2(n157), .B1(A[6]), .B2(n154), .C1(B[6]), .C2(
        n151), .ZN(n25) );
  NAND2_X1 U65 ( .A1(n20), .A2(n21), .ZN(n135) );
  AOI222_X1 U66 ( .A1(E[4]), .A2(n166), .B1(D[4]), .B2(n163), .C1(F[4]), .C2(
        n160), .ZN(n21) );
  AOI222_X1 U67 ( .A1(C[4]), .A2(n157), .B1(A[4]), .B2(n154), .C1(B[4]), .C2(
        n151), .ZN(n20) );
  NAND2_X1 U68 ( .A1(n16), .A2(n17), .ZN(n137) );
  AOI222_X1 U69 ( .A1(E[2]), .A2(n166), .B1(D[2]), .B2(n163), .C1(F[2]), .C2(
        n160), .ZN(n17) );
  AOI222_X1 U70 ( .A1(C[2]), .A2(n157), .B1(A[2]), .B2(n154), .C1(B[2]), .C2(
        n151), .ZN(n16) );
  NAND2_X1 U71 ( .A1(n27), .A2(n28), .ZN(n132) );
  AOI222_X1 U72 ( .A1(E[7]), .A2(n166), .B1(D[7]), .B2(n163), .C1(F[7]), .C2(
        n160), .ZN(n28) );
  AOI222_X1 U73 ( .A1(C[7]), .A2(n157), .B1(A[7]), .B2(n154), .C1(B[7]), .C2(
        n151), .ZN(n27) );
  NAND2_X1 U74 ( .A1(n22), .A2(n24), .ZN(n134) );
  AOI222_X1 U75 ( .A1(E[5]), .A2(n166), .B1(D[5]), .B2(n163), .C1(F[5]), .C2(
        n160), .ZN(n24) );
  AOI222_X1 U76 ( .A1(C[5]), .A2(n157), .B1(A[5]), .B2(n154), .C1(B[5]), .C2(
        n151), .ZN(n22) );
  NAND2_X1 U77 ( .A1(n18), .A2(n19), .ZN(n136) );
  AOI222_X1 U78 ( .A1(E[3]), .A2(n166), .B1(D[3]), .B2(n163), .C1(F[3]), .C2(
        n160), .ZN(n19) );
  AOI222_X1 U79 ( .A1(C[3]), .A2(n157), .B1(A[3]), .B2(n154), .C1(B[3]), .C2(
        n151), .ZN(n18) );
  NAND2_X1 U80 ( .A1(n75), .A2(n76), .ZN(n107) );
  AOI222_X1 U81 ( .A1(E[31]), .A2(n164), .B1(D[31]), .B2(n161), .C1(F[31]), 
        .C2(n158), .ZN(n76) );
  AOI222_X1 U82 ( .A1(C[31]), .A2(n155), .B1(A[31]), .B2(n152), .C1(B[31]), 
        .C2(n149), .ZN(n75) );
  NAND2_X1 U83 ( .A1(n55), .A2(n56), .ZN(n117) );
  AOI222_X1 U84 ( .A1(E[21]), .A2(n164), .B1(D[21]), .B2(n161), .C1(F[21]), 
        .C2(n158), .ZN(n56) );
  AOI222_X1 U85 ( .A1(C[21]), .A2(n155), .B1(A[21]), .B2(n152), .C1(B[21]), 
        .C2(n149), .ZN(n55) );
  NAND2_X1 U86 ( .A1(n49), .A2(n50), .ZN(n120) );
  AOI222_X1 U87 ( .A1(E[18]), .A2(n165), .B1(D[18]), .B2(n162), .C1(F[18]), 
        .C2(n159), .ZN(n50) );
  AOI222_X1 U88 ( .A1(C[18]), .A2(n156), .B1(A[18]), .B2(n153), .C1(B[18]), 
        .C2(n150), .ZN(n49) );
  NAND2_X1 U89 ( .A1(n45), .A2(n46), .ZN(n122) );
  AOI222_X1 U90 ( .A1(E[16]), .A2(n165), .B1(D[16]), .B2(n162), .C1(F[16]), 
        .C2(n159), .ZN(n46) );
  AOI222_X1 U91 ( .A1(C[16]), .A2(n156), .B1(A[16]), .B2(n153), .C1(B[16]), 
        .C2(n150), .ZN(n45) );
  NAND2_X1 U92 ( .A1(n43), .A2(n44), .ZN(n123) );
  AOI222_X1 U93 ( .A1(E[15]), .A2(n165), .B1(D[15]), .B2(n162), .C1(F[15]), 
        .C2(n159), .ZN(n44) );
  AOI222_X1 U94 ( .A1(C[15]), .A2(n156), .B1(A[15]), .B2(n153), .C1(B[15]), 
        .C2(n150), .ZN(n43) );
  NAND2_X1 U95 ( .A1(n41), .A2(n42), .ZN(n124) );
  AOI222_X1 U96 ( .A1(E[14]), .A2(n165), .B1(D[14]), .B2(n162), .C1(F[14]), 
        .C2(n159), .ZN(n42) );
  AOI222_X1 U97 ( .A1(C[14]), .A2(n156), .B1(A[14]), .B2(n153), .C1(B[14]), 
        .C2(n150), .ZN(n41) );
  NAND2_X1 U98 ( .A1(n39), .A2(n40), .ZN(n125) );
  AOI222_X1 U99 ( .A1(E[13]), .A2(n165), .B1(D[13]), .B2(n162), .C1(F[13]), 
        .C2(n159), .ZN(n40) );
  AOI222_X1 U100 ( .A1(C[13]), .A2(n156), .B1(A[13]), .B2(n153), .C1(B[13]), 
        .C2(n150), .ZN(n39) );
  NAND2_X1 U101 ( .A1(n37), .A2(n38), .ZN(n126) );
  AOI222_X1 U102 ( .A1(E[12]), .A2(n165), .B1(D[12]), .B2(n162), .C1(F[12]), 
        .C2(n159), .ZN(n38) );
  AOI222_X1 U103 ( .A1(C[12]), .A2(n156), .B1(A[12]), .B2(n153), .C1(B[12]), 
        .C2(n150), .ZN(n37) );
  NAND2_X1 U104 ( .A1(n35), .A2(n36), .ZN(n127) );
  AOI222_X1 U105 ( .A1(E[11]), .A2(n165), .B1(D[11]), .B2(n162), .C1(F[11]), 
        .C2(n159), .ZN(n36) );
  AOI222_X1 U106 ( .A1(C[11]), .A2(n156), .B1(A[11]), .B2(n153), .C1(B[11]), 
        .C2(n150), .ZN(n35) );
  NAND2_X1 U107 ( .A1(n33), .A2(n34), .ZN(n128) );
  AOI222_X1 U108 ( .A1(E[10]), .A2(n165), .B1(D[10]), .B2(n162), .C1(F[10]), 
        .C2(n159), .ZN(n34) );
  AOI222_X1 U109 ( .A1(C[10]), .A2(n156), .B1(A[10]), .B2(n153), .C1(B[10]), 
        .C2(n150), .ZN(n33) );
  NAND2_X1 U110 ( .A1(n57), .A2(n58), .ZN(n116) );
  AOI222_X1 U111 ( .A1(E[22]), .A2(n164), .B1(D[22]), .B2(n161), .C1(F[22]), 
        .C2(n158), .ZN(n58) );
  AOI222_X1 U112 ( .A1(C[22]), .A2(n155), .B1(A[22]), .B2(n152), .C1(B[22]), 
        .C2(n149), .ZN(n57) );
  NAND2_X1 U113 ( .A1(n53), .A2(n54), .ZN(n118) );
  AOI222_X1 U114 ( .A1(E[20]), .A2(n164), .B1(D[20]), .B2(n161), .C1(F[20]), 
        .C2(n158), .ZN(n54) );
  AOI222_X1 U115 ( .A1(C[20]), .A2(n155), .B1(A[20]), .B2(n152), .C1(B[20]), 
        .C2(n149), .ZN(n53) );
  NAND2_X1 U116 ( .A1(n51), .A2(n52), .ZN(n119) );
  AOI222_X1 U117 ( .A1(E[19]), .A2(n165), .B1(D[19]), .B2(n162), .C1(F[19]), 
        .C2(n159), .ZN(n52) );
  AOI222_X1 U118 ( .A1(C[19]), .A2(n156), .B1(A[19]), .B2(n153), .C1(B[19]), 
        .C2(n150), .ZN(n51) );
  NAND2_X1 U119 ( .A1(n47), .A2(n48), .ZN(n121) );
  AOI222_X1 U120 ( .A1(E[17]), .A2(n165), .B1(D[17]), .B2(n162), .C1(F[17]), 
        .C2(n159), .ZN(n48) );
  AOI222_X1 U121 ( .A1(C[17]), .A2(n156), .B1(A[17]), .B2(n153), .C1(B[17]), 
        .C2(n150), .ZN(n47) );
  NAND2_X1 U122 ( .A1(n29), .A2(n30), .ZN(n131) );
  AOI222_X1 U123 ( .A1(E[8]), .A2(n165), .B1(D[8]), .B2(n162), .C1(F[8]), .C2(
        n159), .ZN(n30) );
  AOI222_X1 U124 ( .A1(C[8]), .A2(n156), .B1(A[8]), .B2(n153), .C1(B[8]), .C2(
        n150), .ZN(n29) );
  NAND2_X1 U125 ( .A1(n31), .A2(n32), .ZN(n129) );
  AOI222_X1 U126 ( .A1(E[9]), .A2(n165), .B1(D[9]), .B2(n162), .C1(F[9]), .C2(
        n159), .ZN(n32) );
  AOI222_X1 U127 ( .A1(C[9]), .A2(n156), .B1(A[9]), .B2(n153), .C1(B[9]), .C2(
        n150), .ZN(n31) );
endmodule


module ff_0 ( clk, rst, d_in, d_out );
  input clk, rst, d_in;
  output d_out;
  wire   N2;

  DFF_X1 d_out_reg ( .D(N2), .CK(clk), .Q(d_out) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in), .ZN(N2) );
endmodule


module reg_N32_4 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U4 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U5 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U6 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U7 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U8 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U9 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U10 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U11 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U12 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U13 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U14 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U15 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U16 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U17 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U18 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U19 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  BUF_X1 U20 ( .A(rst), .Z(n68) );
  BUF_X1 U21 ( .A(rst), .Z(n69) );
  BUF_X1 U22 ( .A(rst), .Z(n70) );
  AND2_X1 U23 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U24 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U25 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U26 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U27 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U28 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U29 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U30 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U31 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U32 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U33 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U34 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U35 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U36 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U37 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
endmodule


module PC_incr ( PC, NPC );
  input [31:0] PC;
  output [31:0] NPC;


  PC_incr_DW01_add_1 add_14 ( .A(PC), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM(NPC) );
endmodule


module reg_en_N32 ( clk, rst, en, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst, en;
  wire   n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, net227477, net227478, net227479, n34, n35,
         n36, n66, n67, n68, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135;
  tri   [31:0] d_in;

  DFF_X1 \d_out_reg[31]  ( .D(n100), .CK(clk), .Q(d_out[31]), .QN(net227479)
         );
  DFF_X1 \d_out_reg[30]  ( .D(n99), .CK(clk), .Q(d_out[30]), .QN(net227478) );
  DFF_X1 \d_out_reg[29]  ( .D(n98), .CK(clk), .Q(d_out[29]), .QN(net227477) );
  DFF_X1 \d_out_reg[28]  ( .D(n97), .CK(clk), .Q(d_out[28]), .QN(n65) );
  DFF_X1 \d_out_reg[27]  ( .D(n96), .CK(clk), .Q(d_out[27]), .QN(n64) );
  DFF_X1 \d_out_reg[26]  ( .D(n95), .CK(clk), .Q(d_out[26]), .QN(n63) );
  DFF_X1 \d_out_reg[25]  ( .D(n94), .CK(clk), .Q(d_out[25]), .QN(n62) );
  DFF_X1 \d_out_reg[24]  ( .D(n93), .CK(clk), .Q(d_out[24]), .QN(n61) );
  DFF_X1 \d_out_reg[23]  ( .D(n92), .CK(clk), .Q(d_out[23]), .QN(n60) );
  DFF_X1 \d_out_reg[22]  ( .D(n91), .CK(clk), .Q(d_out[22]), .QN(n59) );
  DFF_X1 \d_out_reg[21]  ( .D(n90), .CK(clk), .Q(d_out[21]), .QN(n58) );
  DFF_X1 \d_out_reg[20]  ( .D(n89), .CK(clk), .Q(d_out[20]), .QN(n57) );
  DFF_X1 \d_out_reg[19]  ( .D(n88), .CK(clk), .Q(d_out[19]), .QN(n56) );
  DFF_X1 \d_out_reg[18]  ( .D(n87), .CK(clk), .Q(d_out[18]), .QN(n55) );
  DFF_X1 \d_out_reg[17]  ( .D(n86), .CK(clk), .Q(d_out[17]), .QN(n54) );
  DFF_X1 \d_out_reg[16]  ( .D(n85), .CK(clk), .Q(d_out[16]), .QN(n53) );
  DFF_X1 \d_out_reg[15]  ( .D(n84), .CK(clk), .Q(d_out[15]), .QN(n52) );
  DFF_X1 \d_out_reg[14]  ( .D(n83), .CK(clk), .Q(d_out[14]), .QN(n51) );
  DFF_X1 \d_out_reg[13]  ( .D(n82), .CK(clk), .Q(d_out[13]), .QN(n50) );
  DFF_X1 \d_out_reg[12]  ( .D(n81), .CK(clk), .Q(d_out[12]), .QN(n49) );
  DFF_X1 \d_out_reg[11]  ( .D(n80), .CK(clk), .Q(d_out[11]), .QN(n48) );
  DFF_X1 \d_out_reg[10]  ( .D(n79), .CK(clk), .Q(d_out[10]), .QN(n47) );
  DFF_X1 \d_out_reg[9]  ( .D(n78), .CK(clk), .Q(d_out[9]), .QN(n46) );
  DFF_X1 \d_out_reg[8]  ( .D(n77), .CK(clk), .Q(d_out[8]), .QN(n45) );
  DFF_X1 \d_out_reg[7]  ( .D(n76), .CK(clk), .Q(d_out[7]), .QN(n44) );
  DFF_X1 \d_out_reg[6]  ( .D(n75), .CK(clk), .Q(d_out[6]), .QN(n43) );
  DFF_X1 \d_out_reg[5]  ( .D(n74), .CK(clk), .Q(d_out[5]), .QN(n42) );
  DFF_X1 \d_out_reg[4]  ( .D(n73), .CK(clk), .Q(d_out[4]), .QN(n41) );
  DFF_X1 \d_out_reg[3]  ( .D(n72), .CK(clk), .Q(d_out[3]), .QN(n40) );
  DFF_X1 \d_out_reg[2]  ( .D(n71), .CK(clk), .Q(d_out[2]), .QN(n39) );
  DFF_X1 \d_out_reg[1]  ( .D(n70), .CK(clk), .Q(d_out[1]), .QN(n38) );
  DFF_X1 \d_out_reg[0]  ( .D(n69), .CK(clk), .Q(d_out[0]), .QN(n37) );
  BUF_X1 U3 ( .A(n35), .Z(n131) );
  BUF_X1 U4 ( .A(n35), .Z(n130) );
  BUF_X1 U5 ( .A(n35), .Z(n132) );
  BUF_X1 U6 ( .A(n34), .Z(n135) );
  BUF_X1 U7 ( .A(n34), .Z(n133) );
  BUF_X1 U8 ( .A(n34), .Z(n134) );
  NAND2_X1 U9 ( .A1(rst), .A2(n133), .ZN(n35) );
  OAI22_X1 U10 ( .A1(net227477), .A2(n135), .B1(n132), .B2(n66), .ZN(n98) );
  INV_X1 U11 ( .A(d_in[29]), .ZN(n66) );
  OAI22_X1 U12 ( .A1(net227478), .A2(n135), .B1(n132), .B2(n36), .ZN(n99) );
  INV_X1 U13 ( .A(d_in[30]), .ZN(n36) );
  OAI22_X1 U14 ( .A1(n60), .A2(n135), .B1(n132), .B2(n104), .ZN(n92) );
  INV_X1 U15 ( .A(d_in[23]), .ZN(n104) );
  OAI22_X1 U16 ( .A1(n61), .A2(n135), .B1(n132), .B2(n103), .ZN(n93) );
  INV_X1 U17 ( .A(d_in[24]), .ZN(n103) );
  OAI22_X1 U18 ( .A1(n62), .A2(n135), .B1(n132), .B2(n102), .ZN(n94) );
  INV_X1 U19 ( .A(d_in[25]), .ZN(n102) );
  OAI22_X1 U20 ( .A1(n63), .A2(n135), .B1(n132), .B2(n101), .ZN(n95) );
  INV_X1 U21 ( .A(d_in[26]), .ZN(n101) );
  OAI22_X1 U22 ( .A1(n64), .A2(n135), .B1(n132), .B2(n68), .ZN(n96) );
  INV_X1 U23 ( .A(d_in[27]), .ZN(n68) );
  OAI22_X1 U24 ( .A1(n65), .A2(n135), .B1(n132), .B2(n67), .ZN(n97) );
  INV_X1 U25 ( .A(d_in[28]), .ZN(n67) );
  OAI22_X1 U26 ( .A1(net227479), .A2(n133), .B1(n130), .B2(n128), .ZN(n100) );
  INV_X1 U27 ( .A(d_in[31]), .ZN(n128) );
  OAI22_X1 U28 ( .A1(n37), .A2(n133), .B1(n130), .B2(n127), .ZN(n69) );
  INV_X1 U29 ( .A(d_in[0]), .ZN(n127) );
  OAI22_X1 U30 ( .A1(n38), .A2(n133), .B1(n130), .B2(n126), .ZN(n70) );
  INV_X1 U31 ( .A(d_in[1]), .ZN(n126) );
  OAI22_X1 U32 ( .A1(n39), .A2(n133), .B1(n130), .B2(n125), .ZN(n71) );
  INV_X1 U33 ( .A(d_in[2]), .ZN(n125) );
  OAI22_X1 U34 ( .A1(n40), .A2(n133), .B1(n130), .B2(n124), .ZN(n72) );
  INV_X1 U35 ( .A(d_in[3]), .ZN(n124) );
  OAI22_X1 U36 ( .A1(n41), .A2(n133), .B1(n130), .B2(n123), .ZN(n73) );
  INV_X1 U37 ( .A(d_in[4]), .ZN(n123) );
  OAI22_X1 U38 ( .A1(n42), .A2(n133), .B1(n130), .B2(n122), .ZN(n74) );
  INV_X1 U39 ( .A(d_in[5]), .ZN(n122) );
  OAI22_X1 U40 ( .A1(n43), .A2(n133), .B1(n130), .B2(n121), .ZN(n75) );
  INV_X1 U41 ( .A(d_in[6]), .ZN(n121) );
  OAI22_X1 U42 ( .A1(n44), .A2(n133), .B1(n130), .B2(n120), .ZN(n76) );
  INV_X1 U43 ( .A(d_in[7]), .ZN(n120) );
  OAI22_X1 U44 ( .A1(n45), .A2(n133), .B1(n130), .B2(n119), .ZN(n77) );
  INV_X1 U45 ( .A(d_in[8]), .ZN(n119) );
  OAI22_X1 U46 ( .A1(n46), .A2(n133), .B1(n130), .B2(n118), .ZN(n78) );
  INV_X1 U47 ( .A(d_in[9]), .ZN(n118) );
  OAI22_X1 U48 ( .A1(n47), .A2(n134), .B1(n130), .B2(n117), .ZN(n79) );
  INV_X1 U49 ( .A(d_in[10]), .ZN(n117) );
  OAI22_X1 U50 ( .A1(n48), .A2(n134), .B1(n131), .B2(n116), .ZN(n80) );
  INV_X1 U51 ( .A(d_in[11]), .ZN(n116) );
  OAI22_X1 U52 ( .A1(n49), .A2(n134), .B1(n131), .B2(n115), .ZN(n81) );
  INV_X1 U53 ( .A(d_in[12]), .ZN(n115) );
  OAI22_X1 U54 ( .A1(n50), .A2(n134), .B1(n131), .B2(n114), .ZN(n82) );
  INV_X1 U55 ( .A(d_in[13]), .ZN(n114) );
  OAI22_X1 U56 ( .A1(n51), .A2(n134), .B1(n131), .B2(n113), .ZN(n83) );
  INV_X1 U57 ( .A(d_in[14]), .ZN(n113) );
  OAI22_X1 U58 ( .A1(n52), .A2(n134), .B1(n131), .B2(n112), .ZN(n84) );
  INV_X1 U59 ( .A(d_in[15]), .ZN(n112) );
  OAI22_X1 U60 ( .A1(n53), .A2(n134), .B1(n131), .B2(n111), .ZN(n85) );
  INV_X1 U61 ( .A(d_in[16]), .ZN(n111) );
  OAI22_X1 U62 ( .A1(n54), .A2(n134), .B1(n131), .B2(n110), .ZN(n86) );
  INV_X1 U63 ( .A(d_in[17]), .ZN(n110) );
  OAI22_X1 U64 ( .A1(n55), .A2(n134), .B1(n131), .B2(n109), .ZN(n87) );
  INV_X1 U65 ( .A(d_in[18]), .ZN(n109) );
  OAI22_X1 U66 ( .A1(n56), .A2(n134), .B1(n131), .B2(n108), .ZN(n88) );
  INV_X1 U67 ( .A(d_in[19]), .ZN(n108) );
  OAI22_X1 U68 ( .A1(n57), .A2(n134), .B1(n131), .B2(n107), .ZN(n89) );
  INV_X1 U69 ( .A(d_in[20]), .ZN(n107) );
  OAI22_X1 U70 ( .A1(n58), .A2(n134), .B1(n131), .B2(n106), .ZN(n90) );
  INV_X1 U71 ( .A(d_in[21]), .ZN(n106) );
  OAI22_X1 U72 ( .A1(n59), .A2(n135), .B1(n131), .B2(n105), .ZN(n91) );
  INV_X1 U73 ( .A(d_in[22]), .ZN(n105) );
  NAND2_X1 U74 ( .A1(n129), .A2(rst), .ZN(n34) );
  INV_X1 U75 ( .A(en), .ZN(n129) );
endmodule


module MUX21_GENERIC_N32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n3, n4, n5, n6;
  assign n3 = SEL;

  MUX21_90 M_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_89 M_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_88 M_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_87 M_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_86 M_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_85 M_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_84 M_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_83 M_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_82 M_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_81 M_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_80 M_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_79 M_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_78 M_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_77 M_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_76 M_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_75 M_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_74 M_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_73 M_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_72 M_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_71 M_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_70 M_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_69 M_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_68 M_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_67 M_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_66 M_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_65 M_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_64 M_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_63 M_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_62 M_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_61 M_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_31 M_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_30 M_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n4) );
  BUF_X1 U2 ( .A(n3), .Z(n5) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module reg_N32_5 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U7 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U8 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U9 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U10 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U11 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U12 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U13 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U14 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  AND2_X1 U15 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U16 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U17 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U20 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U21 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U22 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U23 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U24 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U25 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U26 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U27 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U28 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U29 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U30 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U31 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U32 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U33 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U34 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U35 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
endmodule


module reg_N32_6 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U10 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U11 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U14 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U15 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U16 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U17 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U18 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U19 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U20 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U21 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U22 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  AND2_X1 U23 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U24 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U25 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U26 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U27 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U28 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U29 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U30 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U31 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U32 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U33 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U34 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U35 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U36 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U37 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
endmodule


module reg_N32_10 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U4 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U5 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U6 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U7 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U8 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U9 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U10 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U11 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U12 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U13 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U14 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U15 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U16 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U17 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U18 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U19 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U20 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U21 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U22 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U23 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U24 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U25 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U26 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U27 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U28 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U29 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U30 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U31 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U32 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U33 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U34 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
  BUF_X1 U35 ( .A(rst), .Z(n68) );
  BUF_X1 U36 ( .A(rst), .Z(n69) );
  BUF_X1 U37 ( .A(rst), .Z(n70) );
endmodule


module MUX21_GENERIC_N32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_0 M_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_217 M_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_216 M_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_215 M_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_214 M_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_213 M_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_212 M_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_211 M_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_210 M_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_209 M_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_208 M_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_207 M_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_206 M_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_205 M_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_204 M_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_203 M_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_202 M_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_201 M_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_200 M_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_199 M_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_198 M_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_197 M_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_196 M_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_195 M_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_194 M_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_193 M_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_192 M_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_191 M_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_190 M_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_189 M_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_188 M_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_187 M_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module sign_ext_Nstart26_Nend32 ( Ain, Aout );
  input [25:0] Ain;
  output [31:0] Aout;
  wire   Aout_31;
  assign Aout[31] = Aout_31;
  assign Aout[30] = Aout_31;
  assign Aout[29] = Aout_31;
  assign Aout[28] = Aout_31;
  assign Aout[27] = Aout_31;
  assign Aout[26] = Aout_31;
  assign Aout[25] = Aout_31;
  assign Aout_31 = Ain[25];
  assign Aout[24] = Ain[24];
  assign Aout[23] = Ain[23];
  assign Aout[22] = Ain[22];
  assign Aout[21] = Ain[21];
  assign Aout[20] = Ain[20];
  assign Aout[19] = Ain[19];
  assign Aout[18] = Ain[18];
  assign Aout[17] = Ain[17];
  assign Aout[16] = Ain[16];
  assign Aout[15] = Ain[15];
  assign Aout[14] = Ain[14];
  assign Aout[13] = Ain[13];
  assign Aout[12] = Ain[12];
  assign Aout[11] = Ain[11];
  assign Aout[10] = Ain[10];
  assign Aout[9] = Ain[9];
  assign Aout[8] = Ain[8];
  assign Aout[7] = Ain[7];
  assign Aout[6] = Ain[6];
  assign Aout[5] = Ain[5];
  assign Aout[4] = Ain[4];
  assign Aout[3] = Ain[3];
  assign Aout[2] = Ain[2];
  assign Aout[1] = Ain[1];
  assign Aout[0] = Ain[0];

endmodule


module sign_ext_Nstart16_Nend32 ( Ain, Aout );
  input [15:0] Ain;
  output [31:0] Aout;
  wire   Aout_31;
  assign Aout[31] = Aout_31;
  assign Aout[30] = Aout_31;
  assign Aout[29] = Aout_31;
  assign Aout[28] = Aout_31;
  assign Aout[27] = Aout_31;
  assign Aout[26] = Aout_31;
  assign Aout[25] = Aout_31;
  assign Aout[24] = Aout_31;
  assign Aout[23] = Aout_31;
  assign Aout[22] = Aout_31;
  assign Aout[21] = Aout_31;
  assign Aout[20] = Aout_31;
  assign Aout[19] = Aout_31;
  assign Aout[18] = Aout_31;
  assign Aout[17] = Aout_31;
  assign Aout[16] = Aout_31;
  assign Aout[15] = Aout_31;
  assign Aout_31 = Ain[15];
  assign Aout[14] = Ain[14];
  assign Aout[13] = Ain[13];
  assign Aout[12] = Ain[12];
  assign Aout[11] = Ain[11];
  assign Aout[10] = Ain[10];
  assign Aout[9] = Ain[9];
  assign Aout[8] = Ain[8];
  assign Aout[7] = Ain[7];
  assign Aout[6] = Ain[6];
  assign Aout[5] = Ain[5];
  assign Aout[4] = Ain[4];
  assign Aout[3] = Ain[3];
  assign Aout[2] = Ain[2];
  assign Aout[1] = Ain[1];
  assign Aout[0] = Ain[0];

endmodule


module reg_N32_13 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module w_reg_file_M8_N8_F4_Nbit32 ( clk, reset, enable, rd1, rd2, wr, add_wr, 
        add_rd1, add_rd2, datain, out1, out2, call, ret, spill, fill, to_mem, 
        from_mem );
  input [4:0] add_wr;
  input [4:0] add_rd1;
  input [4:0] add_rd2;
  input [31:0] datain;
  output [31:0] out1;
  output [31:0] out2;
  output [31:0] to_mem;
  input [31:0] from_mem;
  input clk, reset, enable, rd1, rd2, wr, call, ret;
  output spill, fill;
  wire   \registers[0][31] , \registers[0][30] , \registers[0][29] ,
         \registers[0][28] , \registers[0][27] , \registers[0][26] ,
         \registers[0][25] , \registers[0][24] , \registers[0][23] ,
         \registers[0][22] , \registers[0][21] , \registers[0][20] ,
         \registers[0][19] , \registers[0][18] , \registers[0][17] ,
         \registers[0][16] , \registers[0][15] , \registers[0][14] ,
         \registers[0][13] , \registers[0][12] , \registers[0][11] ,
         \registers[0][10] , \registers[0][9] , \registers[0][8] ,
         \registers[0][7] , \registers[0][6] , \registers[0][5] ,
         \registers[0][4] , \registers[0][3] , \registers[0][2] ,
         \registers[0][1] , \registers[0][0] , \registers[1][31] ,
         \registers[1][30] , \registers[1][29] , \registers[1][28] ,
         \registers[1][27] , \registers[1][26] , \registers[1][25] ,
         \registers[1][24] , \registers[1][23] , \registers[1][22] ,
         \registers[1][21] , \registers[1][20] , \registers[1][19] ,
         \registers[1][18] , \registers[1][17] , \registers[1][16] ,
         \registers[1][15] , \registers[1][14] , \registers[1][13] ,
         \registers[1][12] , \registers[1][11] , \registers[1][10] ,
         \registers[1][9] , \registers[1][8] , \registers[1][7] ,
         \registers[1][6] , \registers[1][5] , \registers[1][4] ,
         \registers[1][3] , \registers[1][2] , \registers[1][1] ,
         \registers[1][0] , \registers[2][31] , \registers[2][30] ,
         \registers[2][29] , \registers[2][28] , \registers[2][27] ,
         \registers[2][26] , \registers[2][25] , \registers[2][24] ,
         \registers[2][23] , \registers[2][22] , \registers[2][21] ,
         \registers[2][20] , \registers[2][19] , \registers[2][18] ,
         \registers[2][17] , \registers[2][16] , \registers[2][15] ,
         \registers[2][14] , \registers[2][13] , \registers[2][12] ,
         \registers[2][11] , \registers[2][10] , \registers[2][9] ,
         \registers[2][8] , \registers[2][7] , \registers[2][6] ,
         \registers[2][5] , \registers[2][4] , \registers[2][3] ,
         \registers[2][2] , \registers[2][1] , \registers[2][0] ,
         \registers[4][31] , \registers[4][30] , \registers[4][29] ,
         \registers[4][28] , \registers[4][27] , \registers[4][26] ,
         \registers[4][25] , \registers[4][24] , \registers[4][23] ,
         \registers[4][22] , \registers[4][21] , \registers[4][20] ,
         \registers[4][19] , \registers[4][18] , \registers[4][17] ,
         \registers[4][16] , \registers[4][15] , \registers[4][14] ,
         \registers[4][13] , \registers[4][12] , \registers[4][11] ,
         \registers[4][10] , \registers[4][9] , \registers[4][8] ,
         \registers[4][7] , \registers[4][6] , \registers[4][5] ,
         \registers[4][4] , \registers[4][3] , \registers[4][2] ,
         \registers[4][1] , \registers[4][0] , \registers[5][31] ,
         \registers[5][30] , \registers[5][29] , \registers[5][28] ,
         \registers[5][27] , \registers[5][26] , \registers[5][25] ,
         \registers[5][24] , \registers[5][23] , \registers[5][22] ,
         \registers[5][21] , \registers[5][20] , \registers[5][19] ,
         \registers[5][18] , \registers[5][17] , \registers[5][16] ,
         \registers[5][15] , \registers[5][14] , \registers[5][13] ,
         \registers[5][12] , \registers[5][11] , \registers[5][10] ,
         \registers[5][9] , \registers[5][8] , \registers[5][7] ,
         \registers[5][6] , \registers[5][5] , \registers[5][4] ,
         \registers[5][3] , \registers[5][2] , \registers[5][1] ,
         \registers[5][0] , \registers[7][31] , \registers[7][30] ,
         \registers[7][29] , \registers[7][28] , \registers[7][27] ,
         \registers[7][26] , \registers[7][25] , \registers[7][24] ,
         \registers[7][23] , \registers[7][22] , \registers[7][21] ,
         \registers[7][20] , \registers[7][19] , \registers[7][18] ,
         \registers[7][17] , \registers[7][16] , \registers[7][15] ,
         \registers[7][14] , \registers[7][13] , \registers[7][12] ,
         \registers[7][11] , \registers[7][10] , \registers[7][9] ,
         \registers[7][8] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[9][31] , \registers[9][30] , \registers[9][29] ,
         \registers[9][28] , \registers[9][27] , \registers[9][26] ,
         \registers[9][25] , \registers[9][24] , \registers[9][23] ,
         \registers[9][22] , \registers[9][21] , \registers[9][20] ,
         \registers[9][19] , \registers[9][18] , \registers[9][17] ,
         \registers[9][16] , \registers[9][15] , \registers[9][14] ,
         \registers[9][13] , \registers[9][12] , \registers[9][11] ,
         \registers[9][10] , \registers[9][9] , \registers[9][8] ,
         \registers[9][7] , \registers[9][6] , \registers[9][5] ,
         \registers[9][4] , \registers[9][3] , \registers[9][2] ,
         \registers[9][1] , \registers[9][0] , \registers[10][31] ,
         \registers[10][30] , \registers[10][29] , \registers[10][28] ,
         \registers[10][27] , \registers[10][26] , \registers[10][25] ,
         \registers[10][24] , \registers[10][23] , \registers[10][22] ,
         \registers[10][21] , \registers[10][20] , \registers[10][19] ,
         \registers[10][18] , \registers[10][17] , \registers[10][16] ,
         \registers[10][15] , \registers[10][14] , \registers[10][13] ,
         \registers[10][12] , \registers[10][11] , \registers[10][10] ,
         \registers[10][9] , \registers[10][8] , \registers[10][7] ,
         \registers[10][6] , \registers[10][5] , \registers[10][4] ,
         \registers[10][3] , \registers[10][2] , \registers[10][1] ,
         \registers[10][0] , \registers[11][31] , \registers[11][30] ,
         \registers[11][29] , \registers[11][28] , \registers[11][27] ,
         \registers[11][26] , \registers[11][25] , \registers[11][24] ,
         \registers[11][23] , \registers[11][22] , \registers[11][21] ,
         \registers[11][20] , \registers[11][19] , \registers[11][18] ,
         \registers[11][17] , \registers[11][16] , \registers[11][15] ,
         \registers[11][14] , \registers[11][13] , \registers[11][12] ,
         \registers[11][11] , \registers[11][10] , \registers[11][9] ,
         \registers[11][8] , \registers[11][7] , \registers[11][6] ,
         \registers[11][5] , \registers[11][4] , \registers[11][3] ,
         \registers[11][2] , \registers[11][1] , \registers[11][0] ,
         \registers[12][31] , \registers[12][30] , \registers[12][29] ,
         \registers[12][28] , \registers[12][27] , \registers[12][26] ,
         \registers[12][25] , \registers[12][24] , \registers[12][23] ,
         \registers[12][22] , \registers[12][21] , \registers[12][20] ,
         \registers[12][19] , \registers[12][18] , \registers[12][17] ,
         \registers[12][16] , \registers[12][15] , \registers[12][14] ,
         \registers[12][13] , \registers[12][12] , \registers[12][11] ,
         \registers[12][10] , \registers[12][9] , \registers[12][8] ,
         \registers[12][7] , \registers[12][6] , \registers[12][5] ,
         \registers[12][4] , \registers[12][3] , \registers[12][2] ,
         \registers[12][1] , \registers[12][0] , \registers[15][31] ,
         \registers[15][30] , \registers[15][29] , \registers[15][28] ,
         \registers[15][27] , \registers[15][26] , \registers[15][25] ,
         \registers[15][24] , \registers[15][23] , \registers[15][22] ,
         \registers[15][21] , \registers[15][20] , \registers[15][19] ,
         \registers[15][18] , \registers[15][17] , \registers[15][16] ,
         \registers[15][15] , \registers[15][14] , \registers[15][13] ,
         \registers[15][12] , \registers[15][11] , \registers[15][10] ,
         \registers[15][9] , \registers[15][8] , \registers[15][7] ,
         \registers[15][6] , \registers[15][5] , \registers[15][4] ,
         \registers[15][3] , \registers[15][2] , \registers[15][1] ,
         \registers[15][0] , \registers[16][31] , \registers[16][30] ,
         \registers[16][29] , \registers[16][28] , \registers[16][27] ,
         \registers[16][26] , \registers[16][25] , \registers[16][24] ,
         \registers[16][23] , \registers[16][22] , \registers[16][21] ,
         \registers[16][20] , \registers[16][19] , \registers[16][18] ,
         \registers[16][17] , \registers[16][16] , \registers[16][15] ,
         \registers[16][14] , \registers[16][13] , \registers[16][12] ,
         \registers[16][11] , \registers[16][10] , \registers[16][9] ,
         \registers[16][8] , \registers[16][7] , \registers[16][6] ,
         \registers[16][5] , \registers[16][4] , \registers[16][3] ,
         \registers[16][2] , \registers[16][1] , \registers[16][0] ,
         \registers[17][31] , \registers[17][30] , \registers[17][29] ,
         \registers[17][28] , \registers[17][27] , \registers[17][26] ,
         \registers[17][25] , \registers[17][24] , \registers[17][23] ,
         \registers[17][22] , \registers[17][21] , \registers[17][20] ,
         \registers[17][19] , \registers[17][18] , \registers[17][17] ,
         \registers[17][16] , \registers[17][15] , \registers[17][14] ,
         \registers[17][13] , \registers[17][12] , \registers[17][11] ,
         \registers[17][10] , \registers[17][9] , \registers[17][8] ,
         \registers[17][7] , \registers[17][6] , \registers[17][5] ,
         \registers[17][4] , \registers[17][3] , \registers[17][2] ,
         \registers[17][1] , \registers[17][0] , \registers[18][31] ,
         \registers[18][30] , \registers[18][29] , \registers[18][28] ,
         \registers[18][27] , \registers[18][26] , \registers[18][25] ,
         \registers[18][24] , \registers[18][23] , \registers[18][22] ,
         \registers[18][21] , \registers[18][20] , \registers[18][19] ,
         \registers[18][18] , \registers[18][17] , \registers[18][16] ,
         \registers[18][15] , \registers[18][14] , \registers[18][13] ,
         \registers[18][12] , \registers[18][11] , \registers[18][10] ,
         \registers[18][9] , \registers[18][8] , \registers[18][7] ,
         \registers[18][6] , \registers[18][5] , \registers[18][4] ,
         \registers[18][3] , \registers[18][2] , \registers[18][1] ,
         \registers[18][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[25][31] , \registers[25][30] ,
         \registers[25][29] , \registers[25][28] , \registers[25][27] ,
         \registers[25][26] , \registers[25][25] , \registers[25][24] ,
         \registers[25][23] , \registers[25][22] , \registers[25][21] ,
         \registers[25][20] , \registers[25][19] , \registers[25][18] ,
         \registers[25][17] , \registers[25][16] , \registers[25][15] ,
         \registers[25][14] , \registers[25][13] , \registers[25][12] ,
         \registers[25][11] , \registers[25][10] , \registers[25][9] ,
         \registers[25][8] , \registers[25][7] , \registers[25][6] ,
         \registers[25][5] , \registers[25][4] , \registers[25][3] ,
         \registers[25][2] , \registers[25][1] , \registers[25][0] ,
         \registers[29][31] , \registers[29][30] , \registers[29][29] ,
         \registers[29][28] , \registers[29][27] , \registers[29][26] ,
         \registers[29][25] , \registers[29][24] , \registers[29][23] ,
         \registers[29][22] , \registers[29][21] , \registers[29][20] ,
         \registers[29][19] , \registers[29][18] , \registers[29][17] ,
         \registers[29][16] , \registers[29][15] , \registers[29][14] ,
         \registers[29][13] , \registers[29][12] , \registers[29][11] ,
         \registers[29][10] , \registers[29][9] , \registers[29][8] ,
         \registers[29][7] , \registers[29][6] , \registers[29][5] ,
         \registers[29][4] , \registers[29][3] , \registers[29][2] ,
         \registers[29][1] , \registers[29][0] , \registers[30][31] ,
         \registers[30][30] , \registers[30][29] , \registers[30][28] ,
         \registers[30][27] , \registers[30][26] , \registers[30][25] ,
         \registers[30][24] , \registers[30][23] , \registers[30][22] ,
         \registers[30][21] , \registers[30][20] , \registers[30][19] ,
         \registers[30][18] , \registers[30][17] , \registers[30][16] ,
         \registers[30][15] , \registers[30][14] , \registers[30][13] ,
         \registers[30][12] , \registers[30][11] , \registers[30][10] ,
         \registers[30][9] , \registers[30][8] , \registers[30][7] ,
         \registers[30][6] , \registers[30][5] , \registers[30][4] ,
         \registers[30][3] , \registers[30][2] , \registers[30][1] ,
         \registers[30][0] , \registers[34][31] , \registers[34][30] ,
         \registers[34][29] , \registers[34][28] , \registers[34][27] ,
         \registers[34][26] , \registers[34][25] , \registers[34][24] ,
         \registers[34][23] , \registers[34][22] , \registers[34][21] ,
         \registers[34][20] , \registers[34][19] , \registers[34][18] ,
         \registers[34][17] , \registers[34][16] , \registers[34][15] ,
         \registers[34][14] , \registers[34][13] , \registers[34][12] ,
         \registers[34][11] , \registers[34][10] , \registers[34][9] ,
         \registers[34][8] , \registers[34][7] , \registers[34][6] ,
         \registers[34][5] , \registers[34][4] , \registers[34][3] ,
         \registers[34][2] , \registers[34][1] , \registers[34][0] ,
         \registers[36][31] , \registers[36][30] , \registers[36][29] ,
         \registers[36][28] , \registers[36][27] , \registers[36][26] ,
         \registers[36][25] , \registers[36][24] , \registers[36][23] ,
         \registers[36][22] , \registers[36][21] , \registers[36][20] ,
         \registers[36][19] , \registers[36][18] , \registers[36][17] ,
         \registers[36][16] , \registers[36][15] , \registers[36][14] ,
         \registers[36][13] , \registers[36][12] , \registers[36][11] ,
         \registers[36][10] , \registers[36][9] , \registers[36][8] ,
         \registers[36][7] , \registers[36][6] , \registers[36][5] ,
         \registers[36][4] , \registers[36][3] , \registers[36][2] ,
         \registers[36][1] , \registers[36][0] , \registers[37][31] ,
         \registers[37][30] , \registers[37][29] , \registers[37][28] ,
         \registers[37][27] , \registers[37][26] , \registers[37][25] ,
         \registers[37][24] , \registers[37][23] , \registers[37][22] ,
         \registers[37][21] , \registers[37][20] , \registers[37][19] ,
         \registers[37][18] , \registers[37][17] , \registers[37][16] ,
         \registers[37][15] , \registers[37][14] , \registers[37][13] ,
         \registers[37][12] , \registers[37][11] , \registers[37][10] ,
         \registers[37][9] , \registers[37][8] , \registers[37][7] ,
         \registers[37][6] , \registers[37][5] , \registers[37][4] ,
         \registers[37][3] , \registers[37][2] , \registers[37][1] ,
         \registers[37][0] , \registers[38][31] , \registers[38][30] ,
         \registers[38][29] , \registers[38][28] , \registers[38][27] ,
         \registers[38][26] , \registers[38][25] , \registers[38][24] ,
         \registers[38][23] , \registers[38][22] , \registers[38][21] ,
         \registers[38][20] , \registers[38][19] , \registers[38][18] ,
         \registers[38][17] , \registers[38][16] , \registers[38][15] ,
         \registers[38][14] , \registers[38][13] , \registers[38][12] ,
         \registers[38][11] , \registers[38][10] , \registers[38][9] ,
         \registers[38][8] , \registers[38][7] , \registers[38][6] ,
         \registers[38][5] , \registers[38][4] , \registers[38][3] ,
         \registers[38][2] , \registers[38][1] , \registers[38][0] ,
         \registers[40][31] , \registers[40][30] , \registers[40][29] ,
         \registers[40][28] , \registers[40][27] , \registers[40][26] ,
         \registers[40][25] , \registers[40][24] , \registers[40][23] ,
         \registers[40][22] , \registers[40][21] , \registers[40][20] ,
         \registers[40][19] , \registers[40][18] , \registers[40][17] ,
         \registers[40][16] , \registers[40][15] , \registers[40][14] ,
         \registers[40][13] , \registers[40][12] , \registers[40][11] ,
         \registers[40][10] , \registers[40][9] , \registers[40][8] ,
         \registers[40][7] , \registers[40][6] , \registers[40][5] ,
         \registers[40][4] , \registers[40][3] , \registers[40][2] ,
         \registers[40][1] , \registers[40][0] , \registers[41][31] ,
         \registers[41][30] , \registers[41][29] , \registers[41][28] ,
         \registers[41][27] , \registers[41][26] , \registers[41][25] ,
         \registers[41][24] , \registers[41][23] , \registers[41][22] ,
         \registers[41][21] , \registers[41][20] , \registers[41][19] ,
         \registers[41][18] , \registers[41][17] , \registers[41][16] ,
         \registers[41][15] , \registers[41][14] , \registers[41][13] ,
         \registers[41][12] , \registers[41][11] , \registers[41][10] ,
         \registers[41][9] , \registers[41][8] , \registers[41][7] ,
         \registers[41][6] , \registers[41][5] , \registers[41][4] ,
         \registers[41][3] , \registers[41][2] , \registers[41][1] ,
         \registers[41][0] , \registers[42][31] , \registers[42][30] ,
         \registers[42][29] , \registers[42][28] , \registers[42][27] ,
         \registers[42][26] , \registers[42][25] , \registers[42][24] ,
         \registers[42][23] , \registers[42][22] , \registers[42][21] ,
         \registers[42][20] , \registers[42][19] , \registers[42][18] ,
         \registers[42][17] , \registers[42][16] , \registers[42][15] ,
         \registers[42][14] , \registers[42][13] , \registers[42][12] ,
         \registers[42][11] , \registers[42][10] , \registers[42][9] ,
         \registers[42][8] , \registers[42][7] , \registers[42][6] ,
         \registers[42][5] , \registers[42][4] , \registers[42][3] ,
         \registers[42][2] , \registers[42][1] , \registers[42][0] ,
         \registers[43][31] , \registers[43][30] , \registers[43][29] ,
         \registers[43][28] , \registers[43][27] , \registers[43][26] ,
         \registers[43][25] , \registers[43][24] , \registers[43][23] ,
         \registers[43][22] , \registers[43][21] , \registers[43][20] ,
         \registers[43][19] , \registers[43][18] , \registers[43][17] ,
         \registers[43][16] , \registers[43][15] , \registers[43][14] ,
         \registers[43][13] , \registers[43][12] , \registers[43][11] ,
         \registers[43][10] , \registers[43][9] , \registers[43][8] ,
         \registers[43][7] , \registers[43][6] , \registers[43][5] ,
         \registers[43][4] , \registers[43][3] , \registers[43][2] ,
         \registers[43][1] , \registers[43][0] , \registers[44][31] ,
         \registers[44][30] , \registers[44][29] , \registers[44][28] ,
         \registers[44][27] , \registers[44][26] , \registers[44][25] ,
         \registers[44][24] , \registers[44][23] , \registers[44][22] ,
         \registers[44][21] , \registers[44][20] , \registers[44][19] ,
         \registers[44][18] , \registers[44][17] , \registers[44][16] ,
         \registers[44][15] , \registers[44][14] , \registers[44][13] ,
         \registers[44][12] , \registers[44][11] , \registers[44][10] ,
         \registers[44][9] , \registers[44][8] , \registers[44][7] ,
         \registers[44][6] , \registers[44][5] , \registers[44][4] ,
         \registers[44][3] , \registers[44][2] , \registers[44][1] ,
         \registers[44][0] , \registers[45][31] , \registers[45][30] ,
         \registers[45][29] , \registers[45][28] , \registers[45][27] ,
         \registers[45][26] , \registers[45][25] , \registers[45][24] ,
         \registers[45][23] , \registers[45][22] , \registers[45][21] ,
         \registers[45][20] , \registers[45][19] , \registers[45][18] ,
         \registers[45][17] , \registers[45][16] , \registers[45][15] ,
         \registers[45][14] , \registers[45][13] , \registers[45][12] ,
         \registers[45][11] , \registers[45][10] , \registers[45][9] ,
         \registers[45][8] , \registers[45][7] , \registers[45][6] ,
         \registers[45][5] , \registers[45][4] , \registers[45][3] ,
         \registers[45][2] , \registers[45][1] , \registers[45][0] ,
         \registers[47][31] , \registers[47][30] , \registers[47][29] ,
         \registers[47][28] , \registers[47][27] , \registers[47][26] ,
         \registers[47][25] , \registers[47][24] , \registers[47][23] ,
         \registers[47][22] , \registers[47][21] , \registers[47][20] ,
         \registers[47][19] , \registers[47][18] , \registers[47][17] ,
         \registers[47][16] , \registers[47][15] , \registers[47][14] ,
         \registers[47][13] , \registers[47][12] , \registers[47][11] ,
         \registers[47][10] , \registers[47][9] , \registers[47][8] ,
         \registers[47][7] , \registers[47][6] , \registers[47][5] ,
         \registers[47][4] , \registers[47][3] , \registers[47][2] ,
         \registers[47][1] , \registers[47][0] , \registers[48][31] ,
         \registers[48][30] , \registers[48][29] , \registers[48][28] ,
         \registers[48][27] , \registers[48][26] , \registers[48][25] ,
         \registers[48][24] , \registers[48][23] , \registers[48][22] ,
         \registers[48][21] , \registers[48][20] , \registers[48][19] ,
         \registers[48][18] , \registers[48][17] , \registers[48][16] ,
         \registers[48][15] , \registers[48][14] , \registers[48][13] ,
         \registers[48][12] , \registers[48][11] , \registers[48][10] ,
         \registers[48][9] , \registers[48][8] , \registers[48][7] ,
         \registers[48][6] , \registers[48][5] , \registers[48][4] ,
         \registers[48][3] , \registers[48][2] , \registers[48][1] ,
         \registers[48][0] , \registers[49][31] , \registers[49][30] ,
         \registers[49][29] , \registers[49][28] , \registers[49][27] ,
         \registers[49][26] , \registers[49][25] , \registers[49][24] ,
         \registers[49][23] , \registers[49][22] , \registers[49][21] ,
         \registers[49][20] , \registers[49][19] , \registers[49][18] ,
         \registers[49][17] , \registers[49][16] , \registers[49][15] ,
         \registers[49][14] , \registers[49][13] , \registers[49][12] ,
         \registers[49][11] , \registers[49][10] , \registers[49][9] ,
         \registers[49][8] , \registers[49][7] , \registers[49][6] ,
         \registers[49][5] , \registers[49][4] , \registers[49][3] ,
         \registers[49][2] , \registers[49][1] , \registers[49][0] ,
         \registers[50][31] , \registers[50][30] , \registers[50][29] ,
         \registers[50][28] , \registers[50][27] , \registers[50][26] ,
         \registers[50][25] , \registers[50][24] , \registers[50][23] ,
         \registers[50][22] , \registers[50][21] , \registers[50][20] ,
         \registers[50][19] , \registers[50][18] , \registers[50][17] ,
         \registers[50][16] , \registers[50][15] , \registers[50][14] ,
         \registers[50][13] , \registers[50][12] , \registers[50][11] ,
         \registers[50][10] , \registers[50][9] , \registers[50][8] ,
         \registers[50][7] , \registers[50][6] , \registers[50][5] ,
         \registers[50][4] , \registers[50][3] , \registers[50][2] ,
         \registers[50][1] , \registers[50][0] , \registers[51][31] ,
         \registers[51][30] , \registers[51][29] , \registers[51][28] ,
         \registers[51][27] , \registers[51][26] , \registers[51][25] ,
         \registers[51][24] , \registers[51][23] , \registers[51][22] ,
         \registers[51][21] , \registers[51][20] , \registers[51][19] ,
         \registers[51][18] , \registers[51][17] , \registers[51][16] ,
         \registers[51][15] , \registers[51][14] , \registers[51][13] ,
         \registers[51][12] , \registers[51][11] , \registers[51][10] ,
         \registers[51][9] , \registers[51][8] , \registers[51][7] ,
         \registers[51][6] , \registers[51][5] , \registers[51][4] ,
         \registers[51][3] , \registers[51][2] , \registers[51][1] ,
         \registers[51][0] , \registers[54][31] , \registers[54][30] ,
         \registers[54][29] , \registers[54][28] , \registers[54][27] ,
         \registers[54][26] , \registers[54][25] , \registers[54][24] ,
         \registers[54][23] , \registers[54][22] , \registers[54][21] ,
         \registers[54][20] , \registers[54][19] , \registers[54][18] ,
         \registers[54][17] , \registers[54][16] , \registers[54][15] ,
         \registers[54][14] , \registers[54][13] , \registers[54][12] ,
         \registers[54][11] , \registers[54][10] , \registers[54][9] ,
         \registers[54][8] , \registers[54][7] , \registers[54][6] ,
         \registers[54][5] , \registers[54][4] , \registers[54][3] ,
         \registers[54][2] , \registers[54][1] , \registers[54][0] ,
         \registers[55][31] , \registers[55][30] , \registers[55][29] ,
         \registers[55][28] , \registers[55][27] , \registers[55][26] ,
         \registers[55][25] , \registers[55][24] , \registers[55][23] ,
         \registers[55][22] , \registers[55][21] , \registers[55][20] ,
         \registers[55][19] , \registers[55][18] , \registers[55][17] ,
         \registers[55][16] , \registers[55][15] , \registers[55][14] ,
         \registers[55][13] , \registers[55][12] , \registers[55][11] ,
         \registers[55][10] , \registers[55][9] , \registers[55][8] ,
         \registers[55][7] , \registers[55][6] , \registers[55][5] ,
         \registers[55][4] , \registers[55][3] , \registers[55][2] ,
         \registers[55][1] , \registers[55][0] , \registers[56][31] ,
         \registers[56][30] , \registers[56][29] , \registers[56][28] ,
         \registers[56][27] , \registers[56][26] , \registers[56][25] ,
         \registers[56][24] , \registers[56][23] , \registers[56][22] ,
         \registers[56][21] , \registers[56][20] , \registers[56][19] ,
         \registers[56][18] , \registers[56][17] , \registers[56][16] ,
         \registers[56][15] , \registers[56][14] , \registers[56][13] ,
         \registers[56][12] , \registers[56][11] , \registers[56][10] ,
         \registers[56][9] , \registers[56][8] , \registers[56][7] ,
         \registers[56][6] , \registers[56][5] , \registers[56][4] ,
         \registers[56][3] , \registers[56][2] , \registers[56][1] ,
         \registers[56][0] , \registers[59][31] , \registers[59][30] ,
         \registers[59][29] , \registers[59][28] , \registers[59][27] ,
         \registers[59][26] , \registers[59][25] , \registers[59][24] ,
         \registers[59][23] , \registers[59][22] , \registers[59][21] ,
         \registers[59][20] , \registers[59][19] , \registers[59][18] ,
         \registers[59][17] , \registers[59][16] , \registers[59][15] ,
         \registers[59][14] , \registers[59][13] , \registers[59][12] ,
         \registers[59][11] , \registers[59][10] , \registers[59][9] ,
         \registers[59][8] , \registers[59][7] , \registers[59][6] ,
         \registers[59][5] , \registers[59][4] , \registers[59][3] ,
         \registers[59][2] , \registers[59][1] , \registers[59][0] ,
         \registers[60][31] , \registers[60][30] , \registers[60][29] ,
         \registers[60][28] , \registers[60][27] , \registers[60][26] ,
         \registers[60][25] , \registers[60][24] , \registers[60][23] ,
         \registers[60][22] , \registers[60][21] , \registers[60][20] ,
         \registers[60][19] , \registers[60][18] , \registers[60][17] ,
         \registers[60][16] , \registers[60][15] , \registers[60][14] ,
         \registers[60][13] , \registers[60][12] , \registers[60][11] ,
         \registers[60][10] , \registers[60][9] , \registers[60][8] ,
         \registers[60][7] , \registers[60][6] , \registers[60][5] ,
         \registers[60][4] , \registers[60][3] , \registers[60][2] ,
         \registers[60][1] , \registers[60][0] , \registers[62][31] ,
         \registers[62][30] , \registers[62][29] , \registers[62][28] ,
         \registers[62][27] , \registers[62][26] , \registers[62][25] ,
         \registers[62][24] , \registers[62][23] , \registers[62][22] ,
         \registers[62][21] , \registers[62][20] , \registers[62][19] ,
         \registers[62][18] , \registers[62][17] , \registers[62][16] ,
         \registers[62][15] , \registers[62][14] , \registers[62][13] ,
         \registers[62][12] , \registers[62][11] , \registers[62][10] ,
         \registers[62][9] , \registers[62][8] , \registers[62][7] ,
         \registers[62][6] , \registers[62][5] , \registers[62][4] ,
         \registers[62][3] , \registers[62][2] , \registers[62][1] ,
         \registers[62][0] , \registers[63][31] , \registers[63][30] ,
         \registers[63][29] , \registers[63][28] , \registers[63][27] ,
         \registers[63][26] , \registers[63][25] , \registers[63][24] ,
         \registers[63][23] , \registers[63][22] , \registers[63][21] ,
         \registers[63][20] , \registers[63][19] , \registers[63][18] ,
         \registers[63][17] , \registers[63][16] , \registers[63][15] ,
         \registers[63][14] , \registers[63][13] , \registers[63][12] ,
         \registers[63][11] , \registers[63][10] , \registers[63][9] ,
         \registers[63][8] , \registers[63][7] , \registers[63][6] ,
         \registers[63][5] , \registers[63][4] , \registers[63][3] ,
         \registers[63][2] , \registers[63][1] , \registers[63][0] ,
         \registers[68][31] , \registers[68][30] , \registers[68][29] ,
         \registers[68][28] , \registers[68][27] , \registers[68][26] ,
         \registers[68][25] , \registers[68][24] , \registers[68][23] ,
         \registers[68][22] , \registers[68][21] , \registers[68][20] ,
         \registers[68][19] , \registers[68][18] , \registers[68][17] ,
         \registers[68][16] , \registers[68][15] , \registers[68][14] ,
         \registers[68][13] , \registers[68][12] , \registers[68][11] ,
         \registers[68][10] , \registers[68][9] , \registers[68][8] ,
         \registers[68][7] , \registers[68][6] , \registers[68][5] ,
         \registers[68][4] , \registers[68][3] , \registers[68][2] ,
         \registers[68][1] , \registers[68][0] , N190, N191, N192,
         \lastcwp[4] , \lastcwp[3] , \lastcwp[2] , \lastcwp[1] , N273, N274,
         N275, N276, N9641, N9908, N9909, N9910, N9921, N9922, N9923, N9924,
         N9925, N9926, N45542, N45543, N45544, N45784, N45785, N45786, N45787,
         N45788, N45789, N46056, N46057, N46058, N46298, N46299, N46300,
         N46301, N46302, N46303, N51637, n7587, n7588, n7589, n7590, n7591,
         n7592, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10187,
         n10188, n10189, n10190, \sub_146/carry[4] , \sub_132/carry[4] ,
         \add_73/carry[1] , \add_73/carry[2] , \add_73/carry[3] ,
         \add_73/carry[4] , \add_73/carry[5] , \sub_71/carry[4] ,
         \r590/carry[5] , n3043, n5522, n6613, n6620, n6621, n6624, n6630,
         n6632, n6634, n6641, n6642, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6671,
         n6674, n6676, n6683, n6684, n6687, n6693, n6695, net226799, net226800,
         net226801, net226802, net226803, net226804, net226805, net226806,
         net226807, net226808, net226809, net226810, net226811, net226812,
         net226813, net226814, net226815, net226816, net226817, net226818,
         net226819, net226820, net226821, net226822, net226823, net226824,
         net226825, net226826, net226827, net226828, net226829, net226830,
         net226831, net226833, net226834, net226835, net226836, net226837,
         net226839, net226840, net226841, net226842, net226843, net226844,
         net226845, net226846, net226847, net226848, net226849, net226850,
         net226851, net226853, net226854, net226855, net226856, net226857,
         net226858, net226859, net226860, net226861, net226862, net226863,
         net226864, net226865, net226866, net226868, net226869, net226870,
         net226871, net226873, net226874, net226875, net226876, net226877,
         net226878, net226879, net226880, net226881, net226882, net226883,
         net226884, net226885, net226886, net226888, net226889, net226890,
         net226891, net226893, net226894, net226895, net226896, net226897,
         net226898, net226899, net226900, net226901, net226902, net226903,
         net226904, net226905, net226906, net226908, net226909, net226910,
         net226911, net226913, net226915, net226917, net226919, net226921,
         net226923, net226925, net226927, net226929, net226931, net226933,
         net226935, net226937, net226939, net226941, net226943, net226945,
         net226947, net226949, net226951, net226953, net226955, net226957,
         net226959, net226961, net226963, net226965, net226967, net226968,
         net226969, net226970, net226971, net226973, net226974, net226975,
         net226976, net226977, net226978, net226979, net226980, net226981,
         net226982, net226983, net226984, net226985, net226986, net226987,
         net226988, net226989, net226990, net226991, net226992, net226993,
         net226994, net226995, net226996, net226997, net226998, net226999,
         net227000, net227001, net227003, net227004, net227005, net227006,
         net227007, net227008, net227009, net227010, net227011, net227012,
         net227014, net227015, net227016, net227017, net227018, net227019,
         net227020, net227021, net227022, net227023, net227024, net227025,
         net227026, net227027, net227028, net227029, net227030, net227032,
         net227033, net227034, net227035, net227036, net227037, net227038,
         net227039, net227040, net227041, net227042, net227043, net227044,
         net227045, net227046, net227047, net227048, net227050, net227051,
         net227052, net227053, net227054, net227055, net227056, net227057,
         net227058, net227059, net227060, net227061, net227062, net227063,
         net227064, net227065, net227066, net227068, net227069, net227070,
         net227071, net227072, net227073, net227074, net227075, net227076,
         net227077, net227078, net227079, net227080, net227081, net227082,
         net227083, net227084, net227086, net227087, net227088, net227089,
         net227090, net227091, net227092, net227093, net227094, net227095,
         net227096, net227097, net227098, net227099, net227100, net227101,
         net227102, net227104, net227105, net227106, net227107, net227108,
         net227109, net227110, net227111, net227112, net227113, net227114,
         net227115, net227116, net227117, net227118, net227119, net227120,
         net227122, net227123, net227124, net227125, net227126, net227127,
         net227128, net227129, net227130, net227131, net227132, net227133,
         net227134, net227135, net227136, net227137, net227138, net227140,
         net227141, net227142, net227143, net227144, net227145, net227146,
         net227147, net227148, net227149, net227150, net227151, net227152,
         net227153, net227154, net227155, net227156, net227158, net227159,
         net227160, net227161, net227162, net227163, net227164, net227165,
         net227166, net227167, net227168, net227169, net227170, net227171,
         net227172, net227173, net227174, net227176, net227177, net227178,
         net227179, net227180, net227181, net227182, net227183, net227184,
         net227185, net227186, net227187, net227188, net227189, net227190,
         net227191, net227192, net227194, net227195, net227196, net227197,
         net227198, net227199, net227200, net227201, net227202, net227203,
         net227204, net227205, net227206, net227207, net227208, net227209,
         net227210, net227212, net227213, net227214, net227215, net227216,
         net227217, net227218, net227219, net227220, net227221, net227222,
         net227223, net227224, net227225, net227226, net227227, net227228,
         net227230, net227231, net227232, net227233, net227234, net227235,
         net227236, net227237, net227238, net227239, net227240, net227241,
         net227242, net227243, net227244, net227245, net227246, net227248,
         net227249, net227250, net227251, net227252, net227253, net227254,
         net227255, net227256, net227257, net227258, net227259, net227260,
         net227261, net227262, net227263, net227264, net227266, net227267,
         net227268, net227269, net227270, net227271, net227272, net227273,
         net227274, net227275, net227276, net227277, net227278, net227279,
         net227280, net227281, net227282, net227284, net227285, net227286,
         net227287, net227288, net227289, net227290, net227291, net227292,
         net227293, net227294, net227295, net227296, net227297, net227298,
         net227299, net227300, net227302, net227303, net227304, net227305,
         net227306, net227307, net227308, net227309, net227310, net227311,
         net227312, net227313, net227314, net227315, net227316, net227317,
         net227318, net227320, net227321, net227322, net227323, net227324,
         net227325, net227326, net227327, net227328, net227329, net227330,
         net227331, net227332, net227333, net227334, net227335, net227336,
         net227338, net227339, net227340, net227341, net227342, net227343,
         net227344, net227345, net227346, net227347, net227348, net227349,
         net227350, net227351, net227352, net227353, net227354, net227356,
         net227357, net227358, net227359, net227360, net227361, net227362,
         net227363, net227364, net227365, net227366, net227367, net227368,
         net227369, net227370, net227371, net227372, net227374, net227375,
         net227376, net227377, net227378, net227379, net227380, net227381,
         net227382, net227383, net227384, net227385, net227386, net227387,
         net227388, net227389, net227390, net227392, net227393, net227394,
         net227395, net227396, net227397, net227398, net227399, net227400,
         net227401, net227402, net227403, net227404, net227405, net227406,
         net227407, net227408, net227410, net227411, net227412, net227413,
         net227414, net227415, net227416, net227417, net227418, net227419,
         net227420, net227421, net227422, net227423, net227424, net227425,
         net227426, net227428, net227429, net227430, net227431, net227432,
         net227433, net227434, net227435, net227436, net227437, net227438,
         net227439, net227440, net227441, net227442, net227443, net227444,
         net227446, net227447, net227448, net227449, net227450, net227451,
         net227452, net227453, net227454, net227455, net227456, net227457,
         net227458, net227459, net227460, net227461, net227462, net227464,
         net227465, net227466, net227467, net227468, net227469, net227470,
         net227471, net227472, net227473, net227474, net227475, net227476,
         n4058, n4059, n4062, n4067, n4070, n4073, n4076, n4079, n4082, n4085,
         n4088, n4090, n4091, n4095, n4098, n4099, n4100, n4101, n4102, n4103,
         n4106, n4107, n4108, n4109, n4110, n4112, n4114, n4117, n4118, n4119,
         n4121, n4123, n4124, n4125, n4126, n4128, n4130, n4131, n4132, n4133,
         n4135, n4137, n4138, n4139, n4140, n4141, n4142, n4145, n4148, n4150,
         n4152, n4153, n4156, n4157, n4159, n4161, n4162, n4163, n4164, n4168,
         n4170, n4171, n4172, n4173, n4175, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4186, n4188, n4189, n4190, n4191, n4192, n4195,
         n4198, n4199, n4200, n4202, n4206, n4207, n4208, n4209, n4211, n4213,
         n4214, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4225, n4226,
         n4227, n4228, n4230, n4232, n4233, n4234, n4235, n4237, n4239, n4240,
         n4241, n4242, n4248, n4251, n4256, n4259, n4262, n4267, n4270, n4273,
         n4275, n4278, n4279, n4282, n4285, n4288, n4291, n4298, n4301, n4306,
         n4309, n4312, n4317, n4320, n4323, n4326, n4329, n4332, n4335, n4338,
         n4341, n4348, n4351, n4356, n4359, n4362, n4367, n4370, n4373, n4376,
         n4379, n4382, n4385, n4388, n4391, n4398, n4401, n4406, n4409, n4412,
         n4417, n4420, n4423, n4426, n4429, n4432, n4435, n4438, n4441, n4448,
         n4451, n4456, n4459, n4462, n4467, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4495, n4498,
         n4499, n4500, n4501, n4502, n4503, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4533, n4611, n4612, n4613, n4614, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4645, n4648, n4649, n4650, n4651, n4652, n4653,
         n4664, n4738, n4739, n4740, n4741, n4742, n4745, n4748, n4749, n4750,
         n4751, n4752, n4753, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4791, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4895, n4898, n4899, n4900, n4901, n4902, n4903, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4924, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5040, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5146, n5147, n5157, n5257, n5259, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5285, n5286, n5288, n5290, n5291,
         n5292, n5293, n5294, n5295, n5298, n5299, n5301, n5302, n5303, n5304,
         n5305, n5307, n5309, n5311, n5312, n5313, n5314, n5315, n5316, n5319,
         n5343, n5442, n5443, n5446, n5447, n5448, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5475, n5476, n5478, n5480,
         n5481, n5482, n5483, n5484, n5485, n5488, n5489, n5491, n5492, n5493,
         n5494, n5495, n5497, n5499, n5501, n5502, n5503, n5504, n5530, n5629,
         n5630, n5631, n5632, n5635, n5636, n5637, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5664, n5665, n5667, n5669,
         n5670, n5671, n5672, n5673, n5674, n5677, n5678, n5680, n5681, n5682,
         n5683, n5684, n5686, n5688, n5690, n5691, n5717, n5816, n5817, n5818,
         n5819, n5820, n5821, n5824, n5825, n5826, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5853, n5854, n5856, n5858,
         n5859, n5860, n5861, n5862, n5863, n5866, n5867, n5869, n5870, n5871,
         n5872, n5873, n5875, n5877, n5889, n6001, n6003, n6005, n6006, n6007,
         n6008, n6009, n6010, n6013, n6014, n6015, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6042, n6043, n6045, n6047,
         n6048, n6049, n6050, n6051, n6052, n6055, n6056, n6058, n6059, n6060,
         n6061, n6062, n6076, n6187, n6188, n6190, n6192, n6194, n6195, n6196,
         n6197, n6198, n6199, n6202, n6203, n6204, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6231, n6232, n6234, n6236,
         n6237, n6238, n6239, n6240, n6241, n6244, n6245, n6247, n6248, n6249,
         n6261, n6374, n6375, n6376, n6377, n6379, n6381, n6383, n6384, n6385,
         n6386, n6387, n6388, n6391, n6392, n6393, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6420, n6421, n6423, n6425,
         n6426, n6427, n6428, n6429, n6430, n6433, n6434, n6436, n6448, n6560,
         n6562, n6563, n6564, n6565, n6566, n6568, n6570, n6572, n6573, n6574,
         n6575, n6576, n6577, n6580, n6581, n6582, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6609, n6610, n6612, n6614,
         n6615, n6616, n6617, n6618, n6619, n6622, n6635, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6769, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6878, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6987, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7096, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7205, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7319, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7428, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7537, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7652, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10282, n10283, n10285,
         n10286, n10287, n10288, n10290, n10292, n10300, n10303, n10306,
         n10315, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10400, n10405,
         n10410, n10413, n10416, n10425, n10444, n10448, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10510, n10511, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10540, n10542,
         n10543, n10544, n10545, n10547, n10549, n10550, n10551, n10552,
         n10554, n10556, n10557, n10558, n10560, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10571, n10573, n10575,
         n10576, n10577, n10578, n10580, n10582, n10583, n10584, n10585,
         n10587, n10589, n10590, n10591, n10592, n10594, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10605, n10607,
         n10608, n10609, n10610, n10612, n10614, n10615, n10616, n10617,
         n10619, n10621, n10622, n10623, n10624, n10626, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10637, n10639,
         n10641, n10642, n10643, n10644, n10646, n10648, n10649, n10650,
         n10651, n10653, n10655, n10656, n10657, n10658, n10660, n10662,
         n10663, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10682, n10683, n10685, n10687, n10688, n10689, n10690, n10691,
         n10694, n10695, n10698, n10700, n10701, n10702, n10703, n10704,
         n10707, n10709, n10711, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11455, n11456, n11457,
         n11458, n11459, n11460, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11843,
         n11848, n11853, n11859, n11868, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11996, n12029, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12149, n12184, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12302, n12338, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12601,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13997,
         n13998, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14009, n14010, n14011, n14012, n14013, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14033, n14034,
         n14058, n14059, n14061, n14062, n14063, n14064, n14066, n14067,
         n14068, n14070, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14213, n14214,
         n14215, n14217, n14218, n14220, n14221, n14222, n14223, n14224,
         n14226, n14228, n14229, n14231, n14232, n14233, n14234, n14236,
         n14237, n14238, n14239, n14240, n14241, n14244, n14245, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14256,
         n14257, n14258, n14259, n14260, n14262, n14263, n14265, n14266,
         n14267, n11498, n11541, n11584, n11627, n11670, n11713, n11756,
         n11799, n11842, n11844, n11845, n11846, n11847, n11849, n11850,
         n11851, n11852, n11854, n11855, n11856, n11857, n11858, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11995, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12148, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12253, n12254, n12255, n12256, n12257, n12258, n12301, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12407, n12408, n12409, n12410, n12411, n12551, n12600,
         n12602, n12652, n12669, n13996, n13999, n14008, n14014, n14015,
         n14032, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14060, n14065, n14069, n14071, n14212, n14216, n14219, n14225,
         n14227, n14230, n14235, n14242, n14243, n14246, n14255, n14261,
         n14264, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055;
  wire   [5:0] swp;
  wire   [31:0] i;
  tri   [31:0] to_mem;
  assign N190 = add_wr[0];
  assign N191 = add_wr[1];
  assign N192 = add_wr[2];
  assign N45542 = add_rd1[0];
  assign N45543 = add_rd1[1];
  assign N45544 = add_rd1[2];
  assign N46056 = add_rd2[0];
  assign N46057 = add_rd2[1];
  assign N46058 = add_rd2[2];
  assign \sub_146/carry[4]  = add_rd2[3];
  assign \sub_132/carry[4]  = add_rd1[3];
  assign \sub_71/carry[4]  = add_wr[3];

  DFF_X1 imspilling_reg ( .D(n10185), .CK(clk), .Q(spill), .QN(n14821) );
  DFF_X1 \swp_reg[0]  ( .D(n10184), .CK(clk), .Q(swp[0]) );
  DFF_X1 imfilling_reg ( .D(n10183), .CK(clk), .Q(fill), .QN(n5522) );
  DFF_X1 \cwp_reg[5]  ( .D(n10181), .CK(clk), .Q(N51637), .QN(n3043) );
  DFF_X1 \swp_reg[1]  ( .D(n10178), .CK(clk), .Q(swp[1]) );
  DFF_X1 \swp_reg[2]  ( .D(n10176), .CK(clk), .Q(swp[2]) );
  DFF_X1 \swp_reg[3]  ( .D(n10174), .CK(clk), .Q(swp[3]) );
  DFF_X1 \swp_reg[5]  ( .D(n10173), .CK(clk), .Q(swp[5]) );
  DFF_X1 \swp_reg[4]  ( .D(n10172), .CK(clk), .Q(swp[4]) );
  DFF_X1 \to_mem_tri_enable_reg[31]  ( .D(n10171), .CK(clk), .Q(n6613), .QN(
        n7662) );
  DFF_X1 \to_mem_tri_enable_reg[30]  ( .D(n10170), .CK(clk), .Q(n6620), .QN(
        n7663) );
  DFF_X1 \to_mem_tri_enable_reg[29]  ( .D(n10169), .CK(clk), .Q(n6621), .QN(
        n7664) );
  DFF_X1 \to_mem_tri_enable_reg[28]  ( .D(n10168), .CK(clk), .Q(n6624), .QN(
        n7665) );
  DFF_X1 \to_mem_tri_enable_reg[27]  ( .D(n10167), .CK(clk), .Q(n6630), .QN(
        n7666) );
  DFF_X1 \to_mem_tri_enable_reg[26]  ( .D(n10166), .CK(clk), .Q(n6632), .QN(
        n7667) );
  DFF_X1 \to_mem_tri_enable_reg[25]  ( .D(n10165), .CK(clk), .Q(n6634), .QN(
        n7668) );
  DFF_X1 \to_mem_tri_enable_reg[24]  ( .D(n10164), .CK(clk), .Q(n6641), .QN(
        n7669) );
  DFF_X1 \to_mem_tri_enable_reg[23]  ( .D(n10163), .CK(clk), .Q(n6642), .QN(
        n7670) );
  DFF_X1 \to_mem_tri_enable_reg[22]  ( .D(n10162), .CK(clk), .Q(n6646), .QN(
        n7671) );
  DFF_X1 \to_mem_tri_enable_reg[21]  ( .D(n10161), .CK(clk), .Q(n6647), .QN(
        n7672) );
  DFF_X1 \to_mem_tri_enable_reg[20]  ( .D(n10160), .CK(clk), .Q(n6648), .QN(
        n7673) );
  DFF_X1 \to_mem_tri_enable_reg[19]  ( .D(n10159), .CK(clk), .Q(n6649), .QN(
        n7674) );
  DFF_X1 \to_mem_tri_enable_reg[18]  ( .D(n10158), .CK(clk), .Q(n6650), .QN(
        n7675) );
  DFF_X1 \to_mem_tri_enable_reg[17]  ( .D(n10157), .CK(clk), .Q(n6651), .QN(
        n7676) );
  DFF_X1 \to_mem_tri_enable_reg[16]  ( .D(n10156), .CK(clk), .Q(n6652), .QN(
        n7677) );
  DFF_X1 \to_mem_tri_enable_reg[15]  ( .D(n10155), .CK(clk), .Q(n6653), .QN(
        n7678) );
  DFF_X1 \to_mem_tri_enable_reg[14]  ( .D(n10154), .CK(clk), .Q(n6654), .QN(
        n7679) );
  DFF_X1 \to_mem_tri_enable_reg[13]  ( .D(n10153), .CK(clk), .Q(n6655), .QN(
        n7680) );
  DFF_X1 \to_mem_tri_enable_reg[12]  ( .D(n10152), .CK(clk), .Q(n6656), .QN(
        n7681) );
  DFF_X1 \to_mem_tri_enable_reg[11]  ( .D(n10151), .CK(clk), .Q(n6657), .QN(
        n7682) );
  DFF_X1 \to_mem_tri_enable_reg[10]  ( .D(n10150), .CK(clk), .Q(n6658), .QN(
        n7683) );
  DFF_X1 \to_mem_tri_enable_reg[9]  ( .D(n10149), .CK(clk), .Q(n6659), .QN(
        n7684) );
  DFF_X1 \to_mem_tri_enable_reg[8]  ( .D(n10148), .CK(clk), .Q(n6660), .QN(
        n7685) );
  DFF_X1 \to_mem_tri_enable_reg[7]  ( .D(n10147), .CK(clk), .Q(n6671), .QN(
        n7686) );
  DFF_X1 \to_mem_tri_enable_reg[6]  ( .D(n10146), .CK(clk), .Q(n6674), .QN(
        n7687) );
  DFF_X1 \to_mem_tri_enable_reg[5]  ( .D(n10145), .CK(clk), .Q(n6676), .QN(
        n7688) );
  DFF_X1 \to_mem_tri_enable_reg[4]  ( .D(n10144), .CK(clk), .Q(n6683), .QN(
        n7689) );
  DFF_X1 \to_mem_tri_enable_reg[3]  ( .D(n10143), .CK(clk), .Q(n6684), .QN(
        n7690) );
  DFF_X1 \to_mem_tri_enable_reg[2]  ( .D(n10142), .CK(clk), .Q(n6687), .QN(
        n7691) );
  DFF_X1 \to_mem_tri_enable_reg[1]  ( .D(n10141), .CK(clk), .Q(n6693), .QN(
        n7692) );
  DFF_X1 \to_mem_tri_enable_reg[0]  ( .D(n10140), .CK(clk), .Q(n6695), .QN(
        n7693) );
  DFF_X1 \i_reg[0]  ( .D(n10138), .CK(clk), .Q(i[0]), .QN(net227476) );
  DFF_X1 \i_reg[5]  ( .D(n10137), .CK(clk), .Q(i[5]), .QN(net227475) );
  DFF_X1 \i_reg[1]  ( .D(n10136), .CK(clk), .Q(i[1]), .QN(net227474) );
  DFF_X1 \i_reg[2]  ( .D(n10135), .CK(clk), .Q(i[2]), .QN(net227473) );
  DFF_X1 \i_reg[3]  ( .D(n10134), .CK(clk), .Q(i[3]), .QN(net227472) );
  DFF_X1 \i_reg[4]  ( .D(n10133), .CK(clk), .Q(i[4]), .QN(net227471) );
  DFF_X1 \lastcwp_reg[5]  ( .D(n10132), .CK(clk), .QN(n7592) );
  DFF_X1 \lastcwp_reg[4]  ( .D(n10131), .CK(clk), .Q(\lastcwp[4] ), .QN(n7591)
         );
  DFF_X1 \lastcwp_reg[3]  ( .D(n10130), .CK(clk), .Q(\lastcwp[3] ), .QN(n7590)
         );
  DFF_X1 \lastcwp_reg[2]  ( .D(n10129), .CK(clk), .Q(\lastcwp[2] ), .QN(n7589)
         );
  DFF_X1 \lastcwp_reg[1]  ( .D(n10128), .CK(clk), .Q(\lastcwp[1] ), .QN(n7588)
         );
  DFF_X1 \lastcwp_reg[0]  ( .D(n10127), .CK(clk), .QN(n7587) );
  DFF_X1 \registers_reg[0][31]  ( .D(n10125), .CK(clk), .Q(\registers[0][31] ), 
        .QN(n15801) );
  DFF_X1 \registers_reg[1][31]  ( .D(n10124), .CK(clk), .Q(\registers[1][31] ), 
        .QN(n15585) );
  DFF_X1 \registers_reg[2][31]  ( .D(n10123), .CK(clk), .Q(\registers[2][31] ), 
        .QN(n14815) );
  DFF_X1 \registers_reg[3][31]  ( .D(n10122), .CK(clk), .Q(net227470), .QN(
        n15781) );
  DFF_X1 \registers_reg[4][31]  ( .D(n10121), .CK(clk), .Q(\registers[4][31] ), 
        .QN(n15458) );
  DFF_X1 \registers_reg[5][31]  ( .D(n10120), .CK(clk), .Q(\registers[5][31] ), 
        .QN(n15318) );
  DFF_X1 \registers_reg[6][31]  ( .D(n10119), .CK(clk), .QN(n12348) );
  DFF_X1 \registers_reg[7][31]  ( .D(n10118), .CK(clk), .Q(\registers[7][31] ), 
        .QN(n15349) );
  DFF_X1 \registers_reg[8][31]  ( .D(n10117), .CK(clk), .Q(net227469), .QN(
        n15239) );
  DFF_X1 \registers_reg[9][31]  ( .D(n10116), .CK(clk), .Q(\registers[9][31] ), 
        .QN(n14358) );
  DFF_X1 \registers_reg[10][31]  ( .D(n10115), .CK(clk), .Q(
        \registers[10][31] ), .QN(n14756) );
  DFF_X1 \registers_reg[11][31]  ( .D(n10114), .CK(clk), .Q(
        \registers[11][31] ), .QN(n14425) );
  DFF_X1 \registers_reg[12][31]  ( .D(n10113), .CK(clk), .Q(
        \registers[12][31] ), .QN(n15691) );
  DFF_X1 \registers_reg[13][31]  ( .D(n10112), .CK(clk), .Q(net227468), .QN(
        n15071) );
  DFF_X1 \registers_reg[14][31]  ( .D(n10111), .CK(clk), .QN(n11903) );
  DFF_X1 \registers_reg[15][31]  ( .D(n10110), .CK(clk), .Q(
        \registers[15][31] ), .QN(n15314) );
  DFF_X1 \registers_reg[16][31]  ( .D(n10109), .CK(clk), .Q(
        \registers[16][31] ), .QN(n15721) );
  DFF_X1 \registers_reg[17][31]  ( .D(n10108), .CK(clk), .Q(
        \registers[17][31] ), .QN(n14627) );
  DFF_X1 \registers_reg[18][31]  ( .D(n10107), .CK(clk), .Q(
        \registers[18][31] ), .QN(n14371) );
  DFF_X1 \registers_reg[19][31]  ( .D(n10106), .CK(clk), .Q(
        \registers[19][31] ), .QN(n15814) );
  DFF_X1 \registers_reg[20][31]  ( .D(n10105), .CK(clk), .QN(n14853) );
  DFF_X1 \registers_reg[21][31]  ( .D(n10104), .CK(clk), .QN(n12307) );
  DFF_X1 \registers_reg[22][31]  ( .D(n10103), .CK(clk), .Q(
        \registers[22][31] ), .QN(n15377) );
  DFF_X1 \registers_reg[23][31]  ( .D(n10102), .CK(clk), .Q(
        \registers[23][31] ), .QN(n15889) );
  DFF_X1 \registers_reg[24][31]  ( .D(n10101), .CK(clk), .Q(net227467), .QN(
        n15209) );
  DFF_X1 \registers_reg[25][31]  ( .D(n10100), .CK(clk), .Q(
        \registers[25][31] ), .QN(n14328) );
  DFF_X1 \registers_reg[26][31]  ( .D(n10099), .CK(clk), .QN(n12355) );
  DFF_X1 \registers_reg[27][31]  ( .D(n10098), .CK(clk), .QN(n12047) );
  DFF_X1 \registers_reg[28][31]  ( .D(n10097), .CK(clk), .Q(net227466), .QN(
        n15032) );
  DFF_X1 \registers_reg[29][31]  ( .D(n10096), .CK(clk), .Q(
        \registers[29][31] ), .QN(n15813) );
  DFF_X1 \registers_reg[30][31]  ( .D(n10095), .CK(clk), .Q(
        \registers[30][31] ), .QN(n14699) );
  DFF_X1 \registers_reg[31][31]  ( .D(n10094), .CK(clk), .Q(net227465), .QN(
        n15757) );
  DFF_X1 \registers_reg[32][31]  ( .D(n10093), .CK(clk), .QN(n12314) );
  DFF_X1 \registers_reg[33][31]  ( .D(n10092), .CK(clk), .QN(n11845) );
  DFF_X1 \registers_reg[34][31]  ( .D(n10091), .CK(clk), .Q(
        \registers[34][31] ), .QN(n15517) );
  DFF_X1 \registers_reg[35][31]  ( .D(n10090), .CK(clk), .Q(net227464), .QN(
        n15590) );
  DFF_X1 \registers_reg[36][31]  ( .D(n10089), .CK(clk), .Q(
        \registers[36][31] ), .QN(n15156) );
  DFF_X1 \registers_reg[37][31]  ( .D(n10088), .CK(clk), .Q(
        \registers[37][31] ), .QN(n14370) );
  DFF_X1 \registers_reg[38][31]  ( .D(n10087), .CK(clk), .Q(
        \registers[38][31] ), .QN(n15041) );
  DFF_X1 \registers_reg[39][31]  ( .D(n10086), .CK(clk), .QN(n12194) );
  DFF_X1 \registers_reg[40][31]  ( .D(n10085), .CK(clk), .Q(
        \registers[40][31] ), .QN(n15150) );
  DFF_X1 \registers_reg[41][31]  ( .D(n10084), .CK(clk), .Q(
        \registers[41][31] ), .QN(n14533) );
  DFF_X1 \registers_reg[42][31]  ( .D(n10083), .CK(clk), .Q(
        \registers[42][31] ), .QN(n15926) );
  DFF_X1 \registers_reg[43][31]  ( .D(n10082), .CK(clk), .Q(
        \registers[43][31] ), .QN(n14887) );
  DFF_X1 \registers_reg[44][31]  ( .D(n10081), .CK(clk), .Q(
        \registers[44][31] ), .QN(n15487) );
  DFF_X1 \registers_reg[45][31]  ( .D(n10080), .CK(clk), .Q(
        \registers[45][31] ), .QN(n14816) );
  DFF_X1 \registers_reg[46][31]  ( .D(n10079), .CK(clk), .QN(n11950) );
  DFF_X1 \registers_reg[47][31]  ( .D(n10078), .CK(clk), .Q(
        \registers[47][31] ), .QN(n14546) );
  DFF_X1 \registers_reg[48][31]  ( .D(n10077), .CK(clk), .Q(
        \registers[48][31] ), .QN(n15551) );
  DFF_X1 \registers_reg[49][31]  ( .D(n10076), .CK(clk), .Q(
        \registers[49][31] ), .QN(n14477) );
  DFF_X1 \registers_reg[50][31]  ( .D(n10075), .CK(clk), .Q(
        \registers[50][31] ), .QN(n15975) );
  DFF_X1 \registers_reg[51][31]  ( .D(n10074), .CK(clk), .Q(
        \registers[51][31] ), .QN(n15427) );
  DFF_X1 \registers_reg[52][31]  ( .D(n10073), .CK(clk), .Q(net227462), .QN(
        n14937) );
  DFF_X1 \registers_reg[53][31]  ( .D(n10072), .CK(clk), .Q(net227461), .QN(
        n15920) );
  DFF_X1 \registers_reg[54][31]  ( .D(n10071), .CK(clk), .Q(
        \registers[54][31] ), .QN(n14535) );
  DFF_X1 \registers_reg[55][31]  ( .D(n10070), .CK(clk), .Q(
        \registers[55][31] ), .QN(n12049) );
  DFF_X1 \registers_reg[56][31]  ( .D(n10069), .CK(clk), .Q(
        \registers[56][31] ), .QN(n15790) );
  DFF_X1 \registers_reg[57][31]  ( .D(n10068), .CK(clk), .Q(net227460), .QN(
        n15034) );
  DFF_X1 \registers_reg[58][31]  ( .D(n10067), .CK(clk), .Q(net227459), .QN(
        n14859) );
  DFF_X1 \registers_reg[59][31]  ( .D(n10066), .CK(clk), .Q(
        \registers[59][31] ), .QN(n14670) );
  DFF_X1 \registers_reg[60][31]  ( .D(n10065), .CK(clk), .Q(
        \registers[60][31] ), .QN(n14634) );
  DFF_X1 \registers_reg[61][31]  ( .D(n10064), .CK(clk), .Q(net227458), .QN(
        n15317) );
  DFF_X1 \registers_reg[62][31]  ( .D(n10063), .CK(clk), .Q(
        \registers[62][31] ), .QN(n14992) );
  DFF_X1 \registers_reg[63][31]  ( .D(n10062), .CK(clk), .Q(
        \registers[63][31] ), .QN(n14281) );
  DFF_X1 \to_mem_reg[31]  ( .D(n10061), .CK(clk), .QN(n7694) );
  DFF_X1 \registers_reg[64][31]  ( .D(n10060), .CK(clk), .Q(net227457), .QN(
        n16034) );
  DFF_X1 \registers_reg[65][31]  ( .D(n10059), .CK(clk), .Q(net227456), .QN(
        n16028) );
  DFF_X1 \registers_reg[66][31]  ( .D(n10058), .CK(clk), .Q(net227455), .QN(
        n16029) );
  DFF_X1 \registers_reg[67][31]  ( .D(n10057), .CK(clk), .QN(n14856) );
  DFF_X1 \registers_reg[68][31]  ( .D(n10056), .CK(clk), .Q(
        \registers[68][31] ), .QN(n16035) );
  DFF_X1 \registers_reg[69][31]  ( .D(n10055), .CK(clk), .Q(net227454), .QN(
        n16033) );
  DFF_X1 \registers_reg[70][31]  ( .D(n10054), .CK(clk), .Q(net227453), .QN(
        n16123) );
  DFF_X1 \registers_reg[0][30]  ( .D(n10053), .CK(clk), .Q(\registers[0][30] ), 
        .QN(n15785) );
  DFF_X1 \registers_reg[1][30]  ( .D(n10052), .CK(clk), .Q(\registers[1][30] ), 
        .QN(n15279) );
  DFF_X1 \registers_reg[2][30]  ( .D(n10051), .CK(clk), .Q(\registers[2][30] ), 
        .QN(n14630) );
  DFF_X1 \registers_reg[3][30]  ( .D(n10050), .CK(clk), .Q(net227452), .QN(
        n15283) );
  DFF_X1 \registers_reg[4][30]  ( .D(n10049), .CK(clk), .Q(\registers[4][30] ), 
        .QN(n15274) );
  DFF_X1 \registers_reg[5][30]  ( .D(n10048), .CK(clk), .Q(\registers[5][30] ), 
        .QN(n14632) );
  DFF_X1 \registers_reg[6][30]  ( .D(n10047), .CK(clk), .QN(n12196) );
  DFF_X1 \registers_reg[7][30]  ( .D(n10046), .CK(clk), .Q(\registers[7][30] ), 
        .QN(n15271) );
  DFF_X1 \registers_reg[8][30]  ( .D(n10045), .CK(clk), .Q(net227451), .QN(
        n14874) );
  DFF_X1 \registers_reg[9][30]  ( .D(n10044), .CK(clk), .Q(\registers[9][30] ), 
        .QN(n14055) );
  DFF_X1 \registers_reg[10][30]  ( .D(n10043), .CK(clk), .Q(
        \registers[10][30] ), .QN(n14629) );
  DFF_X1 \registers_reg[11][30]  ( .D(n10042), .CK(clk), .Q(
        \registers[11][30] ), .QN(n14060) );
  DFF_X1 \registers_reg[12][30]  ( .D(n10041), .CK(clk), .Q(
        \registers[12][30] ), .QN(n15280) );
  DFF_X1 \registers_reg[13][30]  ( .D(n10040), .CK(clk), .Q(net227450), .QN(
        n14870) );
  DFF_X1 \registers_reg[14][30]  ( .D(n10039), .CK(clk), .QN(n11541) );
  DFF_X1 \registers_reg[15][30]  ( .D(n10038), .CK(clk), .Q(
        \registers[15][30] ), .QN(n15270) );
  DFF_X1 \registers_reg[16][30]  ( .D(n10037), .CK(clk), .Q(
        \registers[16][30] ), .QN(n15281) );
  DFF_X1 \registers_reg[17][30]  ( .D(n10036), .CK(clk), .Q(
        \registers[17][30] ), .QN(n14299) );
  DFF_X1 \registers_reg[18][30]  ( .D(n10035), .CK(clk), .Q(
        \registers[18][30] ), .QN(n14057) );
  DFF_X1 \registers_reg[19][30]  ( .D(n10034), .CK(clk), .Q(
        \registers[19][30] ), .QN(n15784) );
  DFF_X1 \registers_reg[20][30]  ( .D(n10033), .CK(clk), .QN(n14822) );
  DFF_X1 \registers_reg[21][30]  ( .D(n10032), .CK(clk), .QN(n12161) );
  DFF_X1 \registers_reg[22][30]  ( .D(n10031), .CK(clk), .Q(
        \registers[22][30] ), .QN(n15273) );
  DFF_X1 \registers_reg[23][30]  ( .D(n10030), .CK(clk), .Q(
        \registers[23][30] ), .QN(n15786) );
  DFF_X1 \registers_reg[24][30]  ( .D(n10029), .CK(clk), .Q(net227449), .QN(
        n14873) );
  DFF_X1 \registers_reg[25][30]  ( .D(n10028), .CK(clk), .Q(
        \registers[25][30] ), .QN(n14054) );
  DFF_X1 \registers_reg[26][30]  ( .D(n10027), .CK(clk), .QN(n12197) );
  DFF_X1 \registers_reg[27][30]  ( .D(n10026), .CK(clk), .QN(n11904) );
  DFF_X1 \registers_reg[28][30]  ( .D(n10025), .CK(clk), .Q(net227448), .QN(
        n14857) );
  DFF_X1 \registers_reg[29][30]  ( .D(n10024), .CK(clk), .Q(
        \registers[29][30] ), .QN(n15783) );
  DFF_X1 \registers_reg[30][30]  ( .D(n10023), .CK(clk), .Q(
        \registers[30][30] ), .QN(n14628) );
  DFF_X1 \registers_reg[31][30]  ( .D(n10022), .CK(clk), .Q(net227447), .QN(
        n15282) );
  DFF_X1 \registers_reg[32][30]  ( .D(n10021), .CK(clk), .QN(n12163) );
  DFF_X1 \registers_reg[33][30]  ( .D(n10020), .CK(clk), .QN(n11498) );
  DFF_X1 \registers_reg[34][30]  ( .D(n10019), .CK(clk), .Q(
        \registers[34][30] ), .QN(n15276) );
  DFF_X1 \registers_reg[35][30]  ( .D(n10018), .CK(clk), .Q(net227446), .QN(
        n15278) );
  DFF_X1 \registers_reg[36][30]  ( .D(n10017), .CK(clk), .Q(
        \registers[36][30] ), .QN(n14872) );
  DFF_X1 \registers_reg[37][30]  ( .D(n10016), .CK(clk), .Q(
        \registers[37][30] ), .QN(n14056) );
  DFF_X1 \registers_reg[38][30]  ( .D(n10015), .CK(clk), .Q(
        \registers[38][30] ), .QN(n14869) );
  DFF_X1 \registers_reg[39][30]  ( .D(n10014), .CK(clk), .QN(n12160) );
  DFF_X1 \registers_reg[40][30]  ( .D(n10013), .CK(clk), .Q(
        \registers[40][30] ), .QN(n14871) );
  DFF_X1 \registers_reg[41][30]  ( .D(n10012), .CK(clk), .Q(
        \registers[41][30] ), .QN(n14069) );
  DFF_X1 \registers_reg[42][30]  ( .D(n10011), .CK(clk), .Q(
        \registers[42][30] ), .QN(n15787) );
  DFF_X1 \registers_reg[43][30]  ( .D(n10010), .CK(clk), .Q(
        \registers[43][30] ), .QN(n14854) );
  DFF_X1 \registers_reg[44][30]  ( .D(n10009), .CK(clk), .Q(
        \registers[44][30] ), .QN(n15275) );
  DFF_X1 \registers_reg[45][30]  ( .D(n10008), .CK(clk), .Q(
        \registers[45][30] ), .QN(n14631) );
  DFF_X1 \registers_reg[46][30]  ( .D(n10007), .CK(clk), .QN(n11670) );
  DFF_X1 \registers_reg[47][30]  ( .D(n10006), .CK(clk), .Q(
        \registers[47][30] ), .QN(n14279) );
  DFF_X1 \registers_reg[48][30]  ( .D(n10005), .CK(clk), .Q(
        \registers[48][30] ), .QN(n15277) );
  DFF_X1 \registers_reg[49][30]  ( .D(n10004), .CK(clk), .Q(
        \registers[49][30] ), .QN(n14065) );
  DFF_X1 \registers_reg[50][30]  ( .D(n10003), .CK(clk), .Q(
        \registers[50][30] ), .QN(n15788) );
  DFF_X1 \registers_reg[51][30]  ( .D(n10002), .CK(clk), .Q(
        \registers[51][30] ), .QN(n15272) );
  DFF_X1 \registers_reg[52][30]  ( .D(n10001), .CK(clk), .Q(net227444), .QN(
        n14855) );
  DFF_X1 \registers_reg[53][30]  ( .D(n10000), .CK(clk), .Q(net227443), .QN(
        n15782) );
  DFF_X1 \registers_reg[54][30]  ( .D(n9999), .CK(clk), .Q(\registers[54][30] ), .QN(n14534) );
  DFF_X1 \registers_reg[55][30]  ( .D(n9998), .CK(clk), .Q(\registers[55][30] ), .QN(n12048) );
  DFF_X1 \registers_reg[56][30]  ( .D(n9997), .CK(clk), .Q(\registers[56][30] ), .QN(n15789) );
  DFF_X1 \registers_reg[57][30]  ( .D(n9996), .CK(clk), .Q(net227442), .QN(
        n15033) );
  DFF_X1 \registers_reg[58][30]  ( .D(n9995), .CK(clk), .Q(net227441), .QN(
        n14858) );
  DFF_X1 \registers_reg[59][30]  ( .D(n9994), .CK(clk), .Q(\registers[59][30] ), .QN(n15315) );
  DFF_X1 \registers_reg[60][30]  ( .D(n9993), .CK(clk), .Q(\registers[60][30] ), .QN(n14633) );
  DFF_X1 \registers_reg[61][30]  ( .D(n9992), .CK(clk), .Q(net227440), .QN(
        n15316) );
  DFF_X1 \registers_reg[62][30]  ( .D(n9991), .CK(clk), .Q(\registers[62][30] ), .QN(n14991) );
  DFF_X1 \registers_reg[63][30]  ( .D(n9990), .CK(clk), .Q(\registers[63][30] ), .QN(n14280) );
  DFF_X1 \to_mem_reg[30]  ( .D(n9989), .CK(clk), .QN(n7695) );
  DFF_X1 \registers_reg[64][30]  ( .D(n9988), .CK(clk), .Q(net227439), .QN(
        n16031) );
  DFF_X1 \registers_reg[65][30]  ( .D(n9987), .CK(clk), .Q(net227438), .QN(
        n16027) );
  DFF_X1 \registers_reg[66][30]  ( .D(n9986), .CK(clk), .Q(net227437), .QN(
        n16026) );
  DFF_X1 \registers_reg[67][30]  ( .D(n9985), .CK(clk), .QN(n14052) );
  DFF_X1 \registers_reg[68][30]  ( .D(n9984), .CK(clk), .Q(\registers[68][30] ), .QN(n16032) );
  DFF_X1 \registers_reg[69][30]  ( .D(n9983), .CK(clk), .Q(net227436), .QN(
        n16030) );
  DFF_X1 \registers_reg[70][30]  ( .D(n9982), .CK(clk), .Q(net227435), .QN(
        n16025) );
  DFF_X1 \registers_reg[0][29]  ( .D(n9981), .CK(clk), .Q(\registers[0][29] ), 
        .QN(n15880) );
  DFF_X1 \registers_reg[1][29]  ( .D(n9980), .CK(clk), .Q(\registers[1][29] ), 
        .QN(n15615) );
  DFF_X1 \registers_reg[2][29]  ( .D(n9979), .CK(clk), .Q(\registers[2][29] ), 
        .QN(n14769) );
  DFF_X1 \registers_reg[3][29]  ( .D(n9978), .CK(clk), .Q(net227434), .QN(
        n15735) );
  DFF_X1 \registers_reg[4][29]  ( .D(n9977), .CK(clk), .Q(\registers[4][29] ), 
        .QN(n15457) );
  DFF_X1 \registers_reg[5][29]  ( .D(n9976), .CK(clk), .Q(\registers[5][29] ), 
        .QN(n14709) );
  DFF_X1 \registers_reg[6][29]  ( .D(n9975), .CK(clk), .QN(n12347) );
  DFF_X1 \registers_reg[7][29]  ( .D(n9974), .CK(clk), .Q(\registers[7][29] ), 
        .QN(n15325) );
  DFF_X1 \registers_reg[8][29]  ( .D(n9973), .CK(clk), .Q(net227433), .QN(
        n15238) );
  DFF_X1 \registers_reg[9][29]  ( .D(n9972), .CK(clk), .Q(\registers[9][29] ), 
        .QN(n14357) );
  DFF_X1 \registers_reg[10][29]  ( .D(n9971), .CK(clk), .Q(\registers[10][29] ), .QN(n14710) );
  DFF_X1 \registers_reg[11][29]  ( .D(n9970), .CK(clk), .Q(\registers[11][29] ), .QN(n14424) );
  DFF_X1 \registers_reg[12][29]  ( .D(n9969), .CK(clk), .Q(\registers[12][29] ), .QN(n15668) );
  DFF_X1 \registers_reg[13][29]  ( .D(n9968), .CK(clk), .Q(net227432), .QN(
        n15070) );
  DFF_X1 \registers_reg[14][29]  ( .D(n9967), .CK(clk), .QN(n11880) );
  DFF_X1 \registers_reg[15][29]  ( .D(n9966), .CK(clk), .Q(\registers[15][29] ), .QN(n15291) );
  DFF_X1 \registers_reg[16][29]  ( .D(n9965), .CK(clk), .Q(\registers[16][29] ), .QN(n15698) );
  DFF_X1 \registers_reg[17][29]  ( .D(n9964), .CK(clk), .Q(\registers[17][29] ), .QN(n14604) );
  DFF_X1 \registers_reg[18][29]  ( .D(n9963), .CK(clk), .Q(\registers[18][29] ), .QN(n14397) );
  DFF_X1 \registers_reg[19][29]  ( .D(n9962), .CK(clk), .Q(\registers[19][29] ), .QN(n15840) );
  DFF_X1 \registers_reg[20][29]  ( .D(n9961), .CK(clk), .QN(n14830) );
  DFF_X1 \registers_reg[21][29]  ( .D(n9960), .CK(clk), .QN(n12204) );
  DFF_X1 \registers_reg[22][29]  ( .D(n9959), .CK(clk), .Q(\registers[22][29] ), .QN(n15390) );
  DFF_X1 \registers_reg[23][29]  ( .D(n9958), .CK(clk), .Q(\registers[23][29] ), .QN(n15902) );
  DFF_X1 \registers_reg[24][29]  ( .D(n9957), .CK(clk), .Q(net227431), .QN(
        n15208) );
  DFF_X1 \registers_reg[25][29]  ( .D(n9956), .CK(clk), .Q(\registers[25][29] ), .QN(n14327) );
  DFF_X1 \registers_reg[26][29]  ( .D(n9955), .CK(clk), .QN(n12354) );
  DFF_X1 \registers_reg[27][29]  ( .D(n9954), .CK(clk), .QN(n12046) );
  DFF_X1 \registers_reg[28][29]  ( .D(n9953), .CK(clk), .Q(net227430), .QN(
        n15031) );
  DFF_X1 \registers_reg[29][29]  ( .D(n9952), .CK(clk), .Q(\registers[29][29] ), .QN(n15839) );
  DFF_X1 \registers_reg[30][29]  ( .D(n9951), .CK(clk), .Q(\registers[30][29] ), .QN(n14677) );
  DFF_X1 \registers_reg[31][29]  ( .D(n9950), .CK(clk), .Q(net227429), .QN(
        n15734) );
  DFF_X1 \registers_reg[32][29]  ( .D(n9949), .CK(clk), .QN(n12339) );
  DFF_X1 \registers_reg[33][29]  ( .D(n9948), .CK(clk), .QN(n11861) );
  DFF_X1 \registers_reg[34][29]  ( .D(n9947), .CK(clk), .Q(\registers[34][29] ), .QN(n15494) );
  DFF_X1 \registers_reg[35][29]  ( .D(n9946), .CK(clk), .Q(net227428), .QN(
        n15614) );
  DFF_X1 \registers_reg[36][29]  ( .D(n9945), .CK(clk), .Q(\registers[36][29] ), .QN(n15169) );
  DFF_X1 \registers_reg[37][29]  ( .D(n9944), .CK(clk), .Q(\registers[37][29] ), .QN(n14396) );
  DFF_X1 \registers_reg[38][29]  ( .D(n9943), .CK(clk), .Q(\registers[38][29] ), .QN(n15054) );
  DFF_X1 \registers_reg[39][29]  ( .D(n9942), .CK(clk), .QN(n12170) );
  DFF_X1 \registers_reg[40][29]  ( .D(n9941), .CK(clk), .Q(\registers[40][29] ), .QN(n15149) );
  DFF_X1 \registers_reg[41][29]  ( .D(n9940), .CK(clk), .Q(\registers[41][29] ), .QN(n14532) );
  DFF_X1 \registers_reg[42][29]  ( .D(n9939), .CK(clk), .Q(\registers[42][29] ), .QN(n15939) );
  DFF_X1 \registers_reg[43][29]  ( .D(n9938), .CK(clk), .Q(\registers[43][29] ), .QN(n14885) );
  DFF_X1 \registers_reg[44][29]  ( .D(n9937), .CK(clk), .Q(\registers[44][29] ), .QN(n15465) );
  DFF_X1 \registers_reg[45][29]  ( .D(n9936), .CK(clk), .Q(\registers[45][29] ), .QN(n14770) );
  DFF_X1 \registers_reg[46][29]  ( .D(n9935), .CK(clk), .QN(n11949) );
  DFF_X1 \registers_reg[47][29]  ( .D(n9934), .CK(clk), .Q(\registers[47][29] ), .QN(n14545) );
  DFF_X1 \registers_reg[48][29]  ( .D(n9933), .CK(clk), .Q(\registers[48][29] ), .QN(n15550) );
  DFF_X1 \registers_reg[49][29]  ( .D(n9932), .CK(clk), .Q(\registers[49][29] ), .QN(n14476) );
  DFF_X1 \registers_reg[50][29]  ( .D(n9931), .CK(clk), .Q(\registers[50][29] ), .QN(n15988) );
  DFF_X1 \registers_reg[51][29]  ( .D(n9930), .CK(clk), .Q(\registers[51][29] ), .QN(n15426) );
  DFF_X1 \registers_reg[52][29]  ( .D(n9929), .CK(clk), .Q(net227426), .QN(
        n14936) );
  DFF_X1 \registers_reg[53][29]  ( .D(n9928), .CK(clk), .Q(net227425), .QN(
        n15968) );
  DFF_X1 \registers_reg[54][29]  ( .D(n9927), .CK(clk), .Q(\registers[54][29] ), .QN(n14597) );
  DFF_X1 \registers_reg[55][29]  ( .D(n9926), .CK(clk), .Q(\registers[55][29] ), .QN(n12159) );
  DFF_X1 \registers_reg[56][29]  ( .D(n9925), .CK(clk), .Q(\registers[56][29] ), .QN(n16012) );
  DFF_X1 \registers_reg[57][29]  ( .D(n9924), .CK(clk), .Q(net227424), .QN(
        n15269) );
  DFF_X1 \registers_reg[58][29]  ( .D(n9923), .CK(clk), .Q(net227423), .QN(
        n14886) );
  DFF_X1 \registers_reg[59][29]  ( .D(n9922), .CK(clk), .Q(\registers[59][29] ), .QN(n15431) );
  DFF_X1 \registers_reg[60][29]  ( .D(n9921), .CK(clk), .Q(\registers[60][29] ), .QN(n14644) );
  DFF_X1 \registers_reg[61][29]  ( .D(n9920), .CK(clk), .Q(net227422), .QN(
        n15660) );
  DFF_X1 \registers_reg[62][29]  ( .D(n9919), .CK(clk), .Q(\registers[62][29] ), .QN(n15122) );
  DFF_X1 \registers_reg[63][29]  ( .D(n9918), .CK(clk), .Q(\registers[63][29] ), .QN(n14483) );
  DFF_X1 \to_mem_reg[29]  ( .D(n9917), .CK(clk), .QN(n7696) );
  DFF_X1 \registers_reg[64][29]  ( .D(n9916), .CK(clk), .Q(net227421), .QN(
        n16148) );
  DFF_X1 \registers_reg[65][29]  ( .D(n9915), .CK(clk), .Q(net227420), .QN(
        n16097) );
  DFF_X1 \registers_reg[66][29]  ( .D(n9914), .CK(clk), .Q(net227419), .QN(
        n16059) );
  DFF_X1 \registers_reg[67][29]  ( .D(n9913), .CK(clk), .QN(n14278) );
  DFF_X1 \registers_reg[68][29]  ( .D(n9912), .CK(clk), .Q(\registers[68][29] ), .QN(n16185) );
  DFF_X1 \registers_reg[69][29]  ( .D(n9911), .CK(clk), .Q(net227418), .QN(
        n16137) );
  DFF_X1 \registers_reg[70][29]  ( .D(n9910), .CK(clk), .Q(net227417), .QN(
        n16049) );
  DFF_X1 \registers_reg[0][28]  ( .D(n9909), .CK(clk), .Q(\registers[0][28] ), 
        .QN(n15879) );
  DFF_X1 \registers_reg[1][28]  ( .D(n9908), .CK(clk), .Q(\registers[1][28] ), 
        .QN(n15636) );
  DFF_X1 \registers_reg[2][28]  ( .D(n9907), .CK(clk), .Q(\registers[2][28] ), 
        .QN(n14767) );
  DFF_X1 \registers_reg[3][28]  ( .D(n9906), .CK(clk), .Q(net227416), .QN(
        n15733) );
  DFF_X1 \registers_reg[4][28]  ( .D(n9905), .CK(clk), .Q(\registers[4][28] ), 
        .QN(n15456) );
  DFF_X1 \registers_reg[5][28]  ( .D(n9904), .CK(clk), .Q(\registers[5][28] ), 
        .QN(n14707) );
  DFF_X1 \registers_reg[6][28]  ( .D(n9903), .CK(clk), .QN(n12346) );
  DFF_X1 \registers_reg[7][28]  ( .D(n9902), .CK(clk), .Q(\registers[7][28] ), 
        .QN(n15324) );
  DFF_X1 \registers_reg[8][28]  ( .D(n9901), .CK(clk), .Q(net227415), .QN(
        n15237) );
  DFF_X1 \registers_reg[9][28]  ( .D(n9900), .CK(clk), .Q(\registers[9][28] ), 
        .QN(n14356) );
  DFF_X1 \registers_reg[10][28]  ( .D(n9899), .CK(clk), .Q(\registers[10][28] ), .QN(n14708) );
  DFF_X1 \registers_reg[11][28]  ( .D(n9898), .CK(clk), .Q(\registers[11][28] ), .QN(n14423) );
  DFF_X1 \registers_reg[12][28]  ( .D(n9897), .CK(clk), .Q(\registers[12][28] ), .QN(n15667) );
  DFF_X1 \registers_reg[13][28]  ( .D(n9896), .CK(clk), .Q(net227414), .QN(
        n15069) );
  DFF_X1 \registers_reg[14][28]  ( .D(n9895), .CK(clk), .QN(n11879) );
  DFF_X1 \registers_reg[15][28]  ( .D(n9894), .CK(clk), .Q(\registers[15][28] ), .QN(n15290) );
  DFF_X1 \registers_reg[16][28]  ( .D(n9893), .CK(clk), .Q(\registers[16][28] ), .QN(n15697) );
  DFF_X1 \registers_reg[17][28]  ( .D(n9892), .CK(clk), .Q(\registers[17][28] ), .QN(n14603) );
  DFF_X1 \registers_reg[18][28]  ( .D(n9891), .CK(clk), .Q(\registers[18][28] ), .QN(n14418) );
  DFF_X1 \registers_reg[19][28]  ( .D(n9890), .CK(clk), .Q(\registers[19][28] ), .QN(n15857) );
  DFF_X1 \registers_reg[20][28]  ( .D(n9889), .CK(clk), .QN(n14829) );
  DFF_X1 \registers_reg[21][28]  ( .D(n9888), .CK(clk), .QN(n12203) );
  DFF_X1 \registers_reg[22][28]  ( .D(n9887), .CK(clk), .Q(\registers[22][28] ), .QN(n15400) );
  DFF_X1 \registers_reg[23][28]  ( .D(n9886), .CK(clk), .Q(\registers[23][28] ), .QN(n15910) );
  DFF_X1 \registers_reg[24][28]  ( .D(n9885), .CK(clk), .Q(net227413), .QN(
        n15207) );
  DFF_X1 \registers_reg[25][28]  ( .D(n9884), .CK(clk), .Q(\registers[25][28] ), .QN(n14326) );
  DFF_X1 \registers_reg[26][28]  ( .D(n9883), .CK(clk), .QN(n12353) );
  DFF_X1 \registers_reg[27][28]  ( .D(n9882), .CK(clk), .QN(n12045) );
  DFF_X1 \registers_reg[28][28]  ( .D(n9881), .CK(clk), .Q(net227412), .QN(
        n15030) );
  DFF_X1 \registers_reg[29][28]  ( .D(n9880), .CK(clk), .Q(\registers[29][28] ), .QN(n15848) );
  DFF_X1 \registers_reg[30][28]  ( .D(n9879), .CK(clk), .Q(\registers[30][28] ), .QN(n14676) );
  DFF_X1 \registers_reg[31][28]  ( .D(n9878), .CK(clk), .Q(net227411), .QN(
        n15732) );
  DFF_X1 \registers_reg[32][28]  ( .D(n9877), .CK(clk), .QN(n12337) );
  DFF_X1 \registers_reg[33][28]  ( .D(n9876), .CK(clk), .QN(n11873) );
  DFF_X1 \registers_reg[34][28]  ( .D(n9875), .CK(clk), .Q(\registers[34][28] ), .QN(n15493) );
  DFF_X1 \registers_reg[35][28]  ( .D(n9874), .CK(clk), .Q(net227410), .QN(
        n15625) );
  DFF_X1 \registers_reg[36][28]  ( .D(n9873), .CK(clk), .Q(\registers[36][28] ), .QN(n15180) );
  DFF_X1 \registers_reg[37][28]  ( .D(n9872), .CK(clk), .Q(\registers[37][28] ), .QN(n14407) );
  DFF_X1 \registers_reg[38][28]  ( .D(n9871), .CK(clk), .Q(\registers[38][28] ), .QN(n15064) );
  DFF_X1 \registers_reg[39][28]  ( .D(n9870), .CK(clk), .QN(n12169) );
  DFF_X1 \registers_reg[40][28]  ( .D(n9869), .CK(clk), .Q(\registers[40][28] ), .QN(n15148) );
  DFF_X1 \registers_reg[41][28]  ( .D(n9868), .CK(clk), .Q(\registers[41][28] ), .QN(n14531) );
  DFF_X1 \registers_reg[42][28]  ( .D(n9867), .CK(clk), .Q(\registers[42][28] ), .QN(n15955) );
  DFF_X1 \registers_reg[43][28]  ( .D(n9866), .CK(clk), .Q(\registers[43][28] ), .QN(n14883) );
  DFF_X1 \registers_reg[44][28]  ( .D(n9865), .CK(clk), .Q(\registers[44][28] ), .QN(n15464) );
  DFF_X1 \registers_reg[45][28]  ( .D(n9864), .CK(clk), .Q(\registers[45][28] ), .QN(n14768) );
  DFF_X1 \registers_reg[46][28]  ( .D(n9863), .CK(clk), .QN(n11948) );
  DFF_X1 \registers_reg[47][28]  ( .D(n9862), .CK(clk), .Q(\registers[47][28] ), .QN(n14544) );
  DFF_X1 \registers_reg[48][28]  ( .D(n9861), .CK(clk), .Q(\registers[48][28] ), .QN(n15549) );
  DFF_X1 \registers_reg[49][28]  ( .D(n9860), .CK(clk), .Q(\registers[49][28] ), .QN(n14475) );
  DFF_X1 \registers_reg[50][28]  ( .D(n9859), .CK(clk), .Q(\registers[50][28] ), .QN(n15997) );
  DFF_X1 \registers_reg[51][28]  ( .D(n9858), .CK(clk), .Q(\registers[51][28] ), .QN(n15425) );
  DFF_X1 \registers_reg[52][28]  ( .D(n9857), .CK(clk), .Q(net227408), .QN(
        n14935) );
  DFF_X1 \registers_reg[53][28]  ( .D(n9856), .CK(clk), .Q(net227407), .QN(
        n15946) );
  DFF_X1 \registers_reg[54][28]  ( .D(n9855), .CK(clk), .Q(\registers[54][28] ), .QN(n14596) );
  DFF_X1 \registers_reg[55][28]  ( .D(n9854), .CK(clk), .Q(\registers[55][28] ), .QN(n12158) );
  DFF_X1 \registers_reg[56][28]  ( .D(n9853), .CK(clk), .Q(\registers[56][28] ), .QN(n16011) );
  DFF_X1 \registers_reg[57][28]  ( .D(n9852), .CK(clk), .Q(net227406), .QN(
        n15268) );
  DFF_X1 \registers_reg[58][28]  ( .D(n9851), .CK(clk), .Q(net227405), .QN(
        n14884) );
  DFF_X1 \registers_reg[59][28]  ( .D(n9850), .CK(clk), .Q(\registers[59][28] ), .QN(n15430) );
  DFF_X1 \registers_reg[60][28]  ( .D(n9849), .CK(clk), .Q(\registers[60][28] ), .QN(n14668) );
  DFF_X1 \registers_reg[61][28]  ( .D(n9848), .CK(clk), .Q(net227404), .QN(
        n15659) );
  DFF_X1 \registers_reg[62][28]  ( .D(n9847), .CK(clk), .Q(\registers[62][28] ), .QN(n15121) );
  DFF_X1 \registers_reg[63][28]  ( .D(n9846), .CK(clk), .Q(\registers[63][28] ), .QN(n14482) );
  DFF_X1 \to_mem_reg[28]  ( .D(n9845), .CK(clk), .QN(n7697) );
  DFF_X1 \registers_reg[64][28]  ( .D(n9844), .CK(clk), .Q(net227403), .QN(
        n16147) );
  DFF_X1 \registers_reg[65][28]  ( .D(n9843), .CK(clk), .Q(net227402), .QN(
        n16096) );
  DFF_X1 \registers_reg[66][28]  ( .D(n9842), .CK(clk), .Q(net227401), .QN(
        n16058) );
  DFF_X1 \registers_reg[67][28]  ( .D(n9841), .CK(clk), .QN(n14277) );
  DFF_X1 \registers_reg[68][28]  ( .D(n9840), .CK(clk), .Q(\registers[68][28] ), .QN(n16184) );
  DFF_X1 \registers_reg[69][28]  ( .D(n9839), .CK(clk), .Q(net227400), .QN(
        n16136) );
  DFF_X1 \registers_reg[70][28]  ( .D(n9838), .CK(clk), .Q(net227399), .QN(
        n16048) );
  DFF_X1 \registers_reg[0][27]  ( .D(n9837), .CK(clk), .Q(\registers[0][27] ), 
        .QN(n15878) );
  DFF_X1 \registers_reg[1][27]  ( .D(n9836), .CK(clk), .Q(\registers[1][27] ), 
        .QN(n15635) );
  DFF_X1 \registers_reg[2][27]  ( .D(n9835), .CK(clk), .Q(\registers[2][27] ), 
        .QN(n14765) );
  DFF_X1 \registers_reg[3][27]  ( .D(n9834), .CK(clk), .Q(net227398), .QN(
        n15731) );
  DFF_X1 \registers_reg[4][27]  ( .D(n9833), .CK(clk), .Q(\registers[4][27] ), 
        .QN(n15455) );
  DFF_X1 \registers_reg[5][27]  ( .D(n9832), .CK(clk), .Q(\registers[5][27] ), 
        .QN(n14705) );
  DFF_X1 \registers_reg[6][27]  ( .D(n9831), .CK(clk), .QN(n12345) );
  DFF_X1 \registers_reg[7][27]  ( .D(n9830), .CK(clk), .Q(\registers[7][27] ), 
        .QN(n15323) );
  DFF_X1 \registers_reg[8][27]  ( .D(n9829), .CK(clk), .Q(net227397), .QN(
        n15236) );
  DFF_X1 \registers_reg[9][27]  ( .D(n9828), .CK(clk), .Q(\registers[9][27] ), 
        .QN(n14355) );
  DFF_X1 \registers_reg[10][27]  ( .D(n9827), .CK(clk), .Q(\registers[10][27] ), .QN(n14706) );
  DFF_X1 \registers_reg[11][27]  ( .D(n9826), .CK(clk), .Q(\registers[11][27] ), .QN(n14422) );
  DFF_X1 \registers_reg[12][27]  ( .D(n9825), .CK(clk), .Q(\registers[12][27] ), .QN(n15666) );
  DFF_X1 \registers_reg[13][27]  ( .D(n9824), .CK(clk), .Q(net227396), .QN(
        n15068) );
  DFF_X1 \registers_reg[14][27]  ( .D(n9823), .CK(clk), .QN(n11878) );
  DFF_X1 \registers_reg[15][27]  ( .D(n9822), .CK(clk), .Q(\registers[15][27] ), .QN(n15289) );
  DFF_X1 \registers_reg[16][27]  ( .D(n9821), .CK(clk), .Q(\registers[16][27] ), .QN(n15696) );
  DFF_X1 \registers_reg[17][27]  ( .D(n9820), .CK(clk), .Q(\registers[17][27] ), .QN(n14602) );
  DFF_X1 \registers_reg[18][27]  ( .D(n9819), .CK(clk), .Q(\registers[18][27] ), .QN(n14417) );
  DFF_X1 \registers_reg[19][27]  ( .D(n9818), .CK(clk), .Q(\registers[19][27] ), .QN(n15856) );
  DFF_X1 \registers_reg[20][27]  ( .D(n9817), .CK(clk), .QN(n14828) );
  DFF_X1 \registers_reg[21][27]  ( .D(n9816), .CK(clk), .QN(n12202) );
  DFF_X1 \registers_reg[22][27]  ( .D(n9815), .CK(clk), .Q(\registers[22][27] ), .QN(n15399) );
  DFF_X1 \registers_reg[23][27]  ( .D(n9814), .CK(clk), .Q(\registers[23][27] ), .QN(n15909) );
  DFF_X1 \registers_reg[24][27]  ( .D(n9813), .CK(clk), .Q(net227395), .QN(
        n15206) );
  DFF_X1 \registers_reg[25][27]  ( .D(n9812), .CK(clk), .Q(\registers[25][27] ), .QN(n14325) );
  DFF_X1 \registers_reg[26][27]  ( .D(n9811), .CK(clk), .QN(n12352) );
  DFF_X1 \registers_reg[27][27]  ( .D(n9810), .CK(clk), .QN(n12044) );
  DFF_X1 \registers_reg[28][27]  ( .D(n9809), .CK(clk), .Q(net227394), .QN(
        n15029) );
  DFF_X1 \registers_reg[29][27]  ( .D(n9808), .CK(clk), .Q(\registers[29][27] ), .QN(n15847) );
  DFF_X1 \registers_reg[30][27]  ( .D(n9807), .CK(clk), .Q(\registers[30][27] ), .QN(n14675) );
  DFF_X1 \registers_reg[31][27]  ( .D(n9806), .CK(clk), .Q(net227393), .QN(
        n15730) );
  DFF_X1 \registers_reg[32][27]  ( .D(n9805), .CK(clk), .QN(n12336) );
  DFF_X1 \registers_reg[33][27]  ( .D(n9804), .CK(clk), .QN(n11872) );
  DFF_X1 \registers_reg[34][27]  ( .D(n9803), .CK(clk), .Q(\registers[34][27] ), .QN(n15492) );
  DFF_X1 \registers_reg[35][27]  ( .D(n9802), .CK(clk), .Q(net227392), .QN(
        n15624) );
  DFF_X1 \registers_reg[36][27]  ( .D(n9801), .CK(clk), .Q(\registers[36][27] ), .QN(n15179) );
  DFF_X1 \registers_reg[37][27]  ( .D(n9800), .CK(clk), .Q(\registers[37][27] ), .QN(n14406) );
  DFF_X1 \registers_reg[38][27]  ( .D(n9799), .CK(clk), .Q(\registers[38][27] ), .QN(n15063) );
  DFF_X1 \registers_reg[39][27]  ( .D(n9798), .CK(clk), .QN(n12168) );
  DFF_X1 \registers_reg[40][27]  ( .D(n9797), .CK(clk), .Q(\registers[40][27] ), .QN(n15147) );
  DFF_X1 \registers_reg[41][27]  ( .D(n9796), .CK(clk), .Q(\registers[41][27] ), .QN(n14530) );
  DFF_X1 \registers_reg[42][27]  ( .D(n9795), .CK(clk), .Q(\registers[42][27] ), .QN(n15954) );
  DFF_X1 \registers_reg[43][27]  ( .D(n9794), .CK(clk), .Q(\registers[43][27] ), .QN(n14881) );
  DFF_X1 \registers_reg[44][27]  ( .D(n9793), .CK(clk), .Q(\registers[44][27] ), .QN(n15463) );
  DFF_X1 \registers_reg[45][27]  ( .D(n9792), .CK(clk), .Q(\registers[45][27] ), .QN(n14766) );
  DFF_X1 \registers_reg[46][27]  ( .D(n9791), .CK(clk), .QN(n11947) );
  DFF_X1 \registers_reg[47][27]  ( .D(n9790), .CK(clk), .Q(\registers[47][27] ), .QN(n14543) );
  DFF_X1 \registers_reg[48][27]  ( .D(n9789), .CK(clk), .Q(\registers[48][27] ), .QN(n15548) );
  DFF_X1 \registers_reg[49][27]  ( .D(n9788), .CK(clk), .Q(\registers[49][27] ), .QN(n14474) );
  DFF_X1 \registers_reg[50][27]  ( .D(n9787), .CK(clk), .Q(\registers[50][27] ), .QN(n15996) );
  DFF_X1 \registers_reg[51][27]  ( .D(n9786), .CK(clk), .Q(\registers[51][27] ), .QN(n15424) );
  DFF_X1 \registers_reg[52][27]  ( .D(n9785), .CK(clk), .Q(net227390), .QN(
        n14934) );
  DFF_X1 \registers_reg[53][27]  ( .D(n9784), .CK(clk), .Q(net227389), .QN(
        n15945) );
  DFF_X1 \registers_reg[54][27]  ( .D(n9783), .CK(clk), .Q(\registers[54][27] ), .QN(n14595) );
  DFF_X1 \registers_reg[55][27]  ( .D(n9782), .CK(clk), .Q(\registers[55][27] ), .QN(n12157) );
  DFF_X1 \registers_reg[56][27]  ( .D(n9781), .CK(clk), .Q(\registers[56][27] ), .QN(n16010) );
  DFF_X1 \registers_reg[57][27]  ( .D(n9780), .CK(clk), .Q(net227388), .QN(
        n15267) );
  DFF_X1 \registers_reg[58][27]  ( .D(n9779), .CK(clk), .Q(net227387), .QN(
        n14882) );
  DFF_X1 \registers_reg[59][27]  ( .D(n9778), .CK(clk), .Q(\registers[59][27] ), .QN(n15429) );
  DFF_X1 \registers_reg[60][27]  ( .D(n9777), .CK(clk), .Q(\registers[60][27] ), .QN(n14667) );
  DFF_X1 \registers_reg[61][27]  ( .D(n9776), .CK(clk), .Q(net227386), .QN(
        n15658) );
  DFF_X1 \registers_reg[62][27]  ( .D(n9775), .CK(clk), .Q(\registers[62][27] ), .QN(n15120) );
  DFF_X1 \registers_reg[63][27]  ( .D(n9774), .CK(clk), .Q(\registers[63][27] ), .QN(n14481) );
  DFF_X1 \to_mem_reg[27]  ( .D(n9773), .CK(clk), .QN(n7698) );
  DFF_X1 \registers_reg[64][27]  ( .D(n9772), .CK(clk), .Q(net227385), .QN(
        n16146) );
  DFF_X1 \registers_reg[65][27]  ( .D(n9771), .CK(clk), .Q(net227384), .QN(
        n16095) );
  DFF_X1 \registers_reg[66][27]  ( .D(n9770), .CK(clk), .Q(net227383), .QN(
        n16057) );
  DFF_X1 \registers_reg[67][27]  ( .D(n9769), .CK(clk), .QN(n14276) );
  DFF_X1 \registers_reg[68][27]  ( .D(n9768), .CK(clk), .Q(\registers[68][27] ), .QN(n16183) );
  DFF_X1 \registers_reg[69][27]  ( .D(n9767), .CK(clk), .Q(net227382), .QN(
        n16135) );
  DFF_X1 \registers_reg[70][27]  ( .D(n9766), .CK(clk), .Q(net227381), .QN(
        n16047) );
  DFF_X1 \registers_reg[0][26]  ( .D(n9765), .CK(clk), .Q(\registers[0][26] ), 
        .QN(n15877) );
  DFF_X1 \registers_reg[1][26]  ( .D(n9764), .CK(clk), .Q(\registers[1][26] ), 
        .QN(n15634) );
  DFF_X1 \registers_reg[2][26]  ( .D(n9763), .CK(clk), .Q(\registers[2][26] ), 
        .QN(n14763) );
  DFF_X1 \registers_reg[3][26]  ( .D(n9762), .CK(clk), .Q(net227380), .QN(
        n15729) );
  DFF_X1 \registers_reg[4][26]  ( .D(n9761), .CK(clk), .Q(\registers[4][26] ), 
        .QN(n15454) );
  DFF_X1 \registers_reg[5][26]  ( .D(n9760), .CK(clk), .Q(\registers[5][26] ), 
        .QN(n14703) );
  DFF_X1 \registers_reg[6][26]  ( .D(n9759), .CK(clk), .QN(n12344) );
  DFF_X1 \registers_reg[7][26]  ( .D(n9758), .CK(clk), .Q(\registers[7][26] ), 
        .QN(n15322) );
  DFF_X1 \registers_reg[8][26]  ( .D(n9757), .CK(clk), .Q(net227379), .QN(
        n15235) );
  DFF_X1 \registers_reg[9][26]  ( .D(n9756), .CK(clk), .Q(\registers[9][26] ), 
        .QN(n14354) );
  DFF_X1 \registers_reg[10][26]  ( .D(n9755), .CK(clk), .Q(\registers[10][26] ), .QN(n14704) );
  DFF_X1 \registers_reg[11][26]  ( .D(n9754), .CK(clk), .Q(\registers[11][26] ), .QN(n14421) );
  DFF_X1 \registers_reg[12][26]  ( .D(n9753), .CK(clk), .Q(\registers[12][26] ), .QN(n15665) );
  DFF_X1 \registers_reg[13][26]  ( .D(n9752), .CK(clk), .Q(net227378), .QN(
        n15067) );
  DFF_X1 \registers_reg[14][26]  ( .D(n9751), .CK(clk), .QN(n11877) );
  DFF_X1 \registers_reg[15][26]  ( .D(n9750), .CK(clk), .Q(\registers[15][26] ), .QN(n15288) );
  DFF_X1 \registers_reg[16][26]  ( .D(n9749), .CK(clk), .Q(\registers[16][26] ), .QN(n15695) );
  DFF_X1 \registers_reg[17][26]  ( .D(n9748), .CK(clk), .Q(\registers[17][26] ), .QN(n14601) );
  DFF_X1 \registers_reg[18][26]  ( .D(n9747), .CK(clk), .Q(\registers[18][26] ), .QN(n14416) );
  DFF_X1 \registers_reg[19][26]  ( .D(n9746), .CK(clk), .Q(\registers[19][26] ), .QN(n15855) );
  DFF_X1 \registers_reg[20][26]  ( .D(n9745), .CK(clk), .QN(n14827) );
  DFF_X1 \registers_reg[21][26]  ( .D(n9744), .CK(clk), .QN(n12201) );
  DFF_X1 \registers_reg[22][26]  ( .D(n9743), .CK(clk), .Q(\registers[22][26] ), .QN(n15398) );
  DFF_X1 \registers_reg[23][26]  ( .D(n9742), .CK(clk), .Q(\registers[23][26] ), .QN(n15908) );
  DFF_X1 \registers_reg[24][26]  ( .D(n9741), .CK(clk), .Q(net227377), .QN(
        n15205) );
  DFF_X1 \registers_reg[25][26]  ( .D(n9740), .CK(clk), .Q(\registers[25][26] ), .QN(n14324) );
  DFF_X1 \registers_reg[26][26]  ( .D(n9739), .CK(clk), .QN(n12351) );
  DFF_X1 \registers_reg[27][26]  ( .D(n9738), .CK(clk), .QN(n12043) );
  DFF_X1 \registers_reg[28][26]  ( .D(n9737), .CK(clk), .Q(net227376), .QN(
        n15028) );
  DFF_X1 \registers_reg[29][26]  ( .D(n9736), .CK(clk), .Q(\registers[29][26] ), .QN(n15846) );
  DFF_X1 \registers_reg[30][26]  ( .D(n9735), .CK(clk), .Q(\registers[30][26] ), .QN(n14674) );
  DFF_X1 \registers_reg[31][26]  ( .D(n9734), .CK(clk), .Q(net227375), .QN(
        n15728) );
  DFF_X1 \registers_reg[32][26]  ( .D(n9733), .CK(clk), .QN(n12335) );
  DFF_X1 \registers_reg[33][26]  ( .D(n9732), .CK(clk), .QN(n11871) );
  DFF_X1 \registers_reg[34][26]  ( .D(n9731), .CK(clk), .Q(\registers[34][26] ), .QN(n15491) );
  DFF_X1 \registers_reg[35][26]  ( .D(n9730), .CK(clk), .Q(net227374), .QN(
        n15623) );
  DFF_X1 \registers_reg[36][26]  ( .D(n9729), .CK(clk), .Q(\registers[36][26] ), .QN(n15178) );
  DFF_X1 \registers_reg[37][26]  ( .D(n9728), .CK(clk), .Q(\registers[37][26] ), .QN(n14405) );
  DFF_X1 \registers_reg[38][26]  ( .D(n9727), .CK(clk), .Q(\registers[38][26] ), .QN(n15062) );
  DFF_X1 \registers_reg[39][26]  ( .D(n9726), .CK(clk), .QN(n12167) );
  DFF_X1 \registers_reg[40][26]  ( .D(n9725), .CK(clk), .Q(\registers[40][26] ), .QN(n15146) );
  DFF_X1 \registers_reg[41][26]  ( .D(n9724), .CK(clk), .Q(\registers[41][26] ), .QN(n14529) );
  DFF_X1 \registers_reg[42][26]  ( .D(n9723), .CK(clk), .Q(\registers[42][26] ), .QN(n15953) );
  DFF_X1 \registers_reg[43][26]  ( .D(n9722), .CK(clk), .Q(\registers[43][26] ), .QN(n14879) );
  DFF_X1 \registers_reg[44][26]  ( .D(n9721), .CK(clk), .Q(\registers[44][26] ), .QN(n15462) );
  DFF_X1 \registers_reg[45][26]  ( .D(n9720), .CK(clk), .Q(\registers[45][26] ), .QN(n14764) );
  DFF_X1 \registers_reg[46][26]  ( .D(n9719), .CK(clk), .QN(n11946) );
  DFF_X1 \registers_reg[47][26]  ( .D(n9718), .CK(clk), .Q(\registers[47][26] ), .QN(n14542) );
  DFF_X1 \registers_reg[48][26]  ( .D(n9717), .CK(clk), .Q(\registers[48][26] ), .QN(n15547) );
  DFF_X1 \registers_reg[49][26]  ( .D(n9716), .CK(clk), .Q(\registers[49][26] ), .QN(n14473) );
  DFF_X1 \registers_reg[50][26]  ( .D(n9715), .CK(clk), .Q(\registers[50][26] ), .QN(n15995) );
  DFF_X1 \registers_reg[51][26]  ( .D(n9714), .CK(clk), .Q(\registers[51][26] ), .QN(n15423) );
  DFF_X1 \registers_reg[52][26]  ( .D(n9713), .CK(clk), .Q(net227372), .QN(
        n14933) );
  DFF_X1 \registers_reg[53][26]  ( .D(n9712), .CK(clk), .Q(net227371), .QN(
        n15944) );
  DFF_X1 \registers_reg[54][26]  ( .D(n9711), .CK(clk), .Q(\registers[54][26] ), .QN(n14594) );
  DFF_X1 \registers_reg[55][26]  ( .D(n9710), .CK(clk), .Q(\registers[55][26] ), .QN(n12156) );
  DFF_X1 \registers_reg[56][26]  ( .D(n9709), .CK(clk), .Q(\registers[56][26] ), .QN(n16009) );
  DFF_X1 \registers_reg[57][26]  ( .D(n9708), .CK(clk), .Q(net227370), .QN(
        n15266) );
  DFF_X1 \registers_reg[58][26]  ( .D(n9707), .CK(clk), .Q(net227369), .QN(
        n14880) );
  DFF_X1 \registers_reg[59][26]  ( .D(n9706), .CK(clk), .Q(\registers[59][26] ), .QN(n15428) );
  DFF_X1 \registers_reg[60][26]  ( .D(n9705), .CK(clk), .Q(\registers[60][26] ), .QN(n14666) );
  DFF_X1 \registers_reg[61][26]  ( .D(n9704), .CK(clk), .Q(net227368), .QN(
        n15657) );
  DFF_X1 \registers_reg[62][26]  ( .D(n9703), .CK(clk), .Q(\registers[62][26] ), .QN(n15119) );
  DFF_X1 \registers_reg[63][26]  ( .D(n9702), .CK(clk), .Q(\registers[63][26] ), .QN(n14480) );
  DFF_X1 \to_mem_reg[26]  ( .D(n9701), .CK(clk), .QN(n7699) );
  DFF_X1 \registers_reg[64][26]  ( .D(n9700), .CK(clk), .Q(net227367), .QN(
        n16145) );
  DFF_X1 \registers_reg[65][26]  ( .D(n9699), .CK(clk), .Q(net227366), .QN(
        n16094) );
  DFF_X1 \registers_reg[66][26]  ( .D(n9698), .CK(clk), .Q(net227365), .QN(
        n16056) );
  DFF_X1 \registers_reg[67][26]  ( .D(n9697), .CK(clk), .QN(n14275) );
  DFF_X1 \registers_reg[68][26]  ( .D(n9696), .CK(clk), .Q(\registers[68][26] ), .QN(n16182) );
  DFF_X1 \registers_reg[69][26]  ( .D(n9695), .CK(clk), .Q(net227364), .QN(
        n16134) );
  DFF_X1 \registers_reg[70][26]  ( .D(n9694), .CK(clk), .Q(net227363), .QN(
        n16046) );
  DFF_X1 \registers_reg[0][25]  ( .D(n9693), .CK(clk), .Q(\registers[0][25] ), 
        .QN(n15876) );
  DFF_X1 \registers_reg[1][25]  ( .D(n9692), .CK(clk), .Q(\registers[1][25] ), 
        .QN(n15633) );
  DFF_X1 \registers_reg[2][25]  ( .D(n9691), .CK(clk), .Q(\registers[2][25] ), 
        .QN(n14761) );
  DFF_X1 \registers_reg[3][25]  ( .D(n9690), .CK(clk), .Q(net227362), .QN(
        n15727) );
  DFF_X1 \registers_reg[4][25]  ( .D(n9689), .CK(clk), .Q(\registers[4][25] ), 
        .QN(n15453) );
  DFF_X1 \registers_reg[5][25]  ( .D(n9688), .CK(clk), .Q(\registers[5][25] ), 
        .QN(n14819) );
  DFF_X1 \registers_reg[6][25]  ( .D(n9687), .CK(clk), .QN(n12343) );
  DFF_X1 \registers_reg[7][25]  ( .D(n9686), .CK(clk), .Q(\registers[7][25] ), 
        .QN(n15321) );
  DFF_X1 \registers_reg[8][25]  ( .D(n9685), .CK(clk), .Q(net227361), .QN(
        n15234) );
  DFF_X1 \registers_reg[9][25]  ( .D(n9684), .CK(clk), .Q(\registers[9][25] ), 
        .QN(n14353) );
  DFF_X1 \registers_reg[10][25]  ( .D(n9683), .CK(clk), .Q(\registers[10][25] ), .QN(n14702) );
  DFF_X1 \registers_reg[11][25]  ( .D(n9682), .CK(clk), .Q(\registers[11][25] ), .QN(n14420) );
  DFF_X1 \registers_reg[12][25]  ( .D(n9681), .CK(clk), .Q(\registers[12][25] ), .QN(n15664) );
  DFF_X1 \registers_reg[13][25]  ( .D(n9680), .CK(clk), .Q(net227360), .QN(
        n15066) );
  DFF_X1 \registers_reg[14][25]  ( .D(n9679), .CK(clk), .QN(n11876) );
  DFF_X1 \registers_reg[15][25]  ( .D(n9678), .CK(clk), .Q(\registers[15][25] ), .QN(n15287) );
  DFF_X1 \registers_reg[16][25]  ( .D(n9677), .CK(clk), .Q(\registers[16][25] ), .QN(n15694) );
  DFF_X1 \registers_reg[17][25]  ( .D(n9676), .CK(clk), .Q(\registers[17][25] ), .QN(n14600) );
  DFF_X1 \registers_reg[18][25]  ( .D(n9675), .CK(clk), .Q(\registers[18][25] ), .QN(n14415) );
  DFF_X1 \registers_reg[19][25]  ( .D(n9674), .CK(clk), .Q(\registers[19][25] ), .QN(n15854) );
  DFF_X1 \registers_reg[20][25]  ( .D(n9673), .CK(clk), .QN(n14826) );
  DFF_X1 \registers_reg[21][25]  ( .D(n9672), .CK(clk), .QN(n12200) );
  DFF_X1 \registers_reg[22][25]  ( .D(n9671), .CK(clk), .Q(\registers[22][25] ), .QN(n15397) );
  DFF_X1 \registers_reg[23][25]  ( .D(n9670), .CK(clk), .Q(\registers[23][25] ), .QN(n15907) );
  DFF_X1 \registers_reg[24][25]  ( .D(n9669), .CK(clk), .Q(net227359), .QN(
        n15204) );
  DFF_X1 \registers_reg[25][25]  ( .D(n9668), .CK(clk), .Q(\registers[25][25] ), .QN(n14323) );
  DFF_X1 \registers_reg[26][25]  ( .D(n9667), .CK(clk), .QN(n12350) );
  DFF_X1 \registers_reg[27][25]  ( .D(n9666), .CK(clk), .QN(n12042) );
  DFF_X1 \registers_reg[28][25]  ( .D(n9665), .CK(clk), .Q(net227358), .QN(
        n15027) );
  DFF_X1 \registers_reg[29][25]  ( .D(n9664), .CK(clk), .Q(\registers[29][25] ), .QN(n15845) );
  DFF_X1 \registers_reg[30][25]  ( .D(n9663), .CK(clk), .Q(\registers[30][25] ), .QN(n14673) );
  DFF_X1 \registers_reg[31][25]  ( .D(n9662), .CK(clk), .Q(net227357), .QN(
        n15726) );
  DFF_X1 \registers_reg[32][25]  ( .D(n9661), .CK(clk), .QN(n12334) );
  DFF_X1 \registers_reg[33][25]  ( .D(n9660), .CK(clk), .QN(n11870) );
  DFF_X1 \registers_reg[34][25]  ( .D(n9659), .CK(clk), .Q(\registers[34][25] ), .QN(n15490) );
  DFF_X1 \registers_reg[35][25]  ( .D(n9658), .CK(clk), .Q(net227356), .QN(
        n15622) );
  DFF_X1 \registers_reg[36][25]  ( .D(n9657), .CK(clk), .Q(\registers[36][25] ), .QN(n15177) );
  DFF_X1 \registers_reg[37][25]  ( .D(n9656), .CK(clk), .Q(\registers[37][25] ), .QN(n14404) );
  DFF_X1 \registers_reg[38][25]  ( .D(n9655), .CK(clk), .Q(\registers[38][25] ), .QN(n15061) );
  DFF_X1 \registers_reg[39][25]  ( .D(n9654), .CK(clk), .QN(n12166) );
  DFF_X1 \registers_reg[40][25]  ( .D(n9653), .CK(clk), .Q(\registers[40][25] ), .QN(n15145) );
  DFF_X1 \registers_reg[41][25]  ( .D(n9652), .CK(clk), .Q(\registers[41][25] ), .QN(n14528) );
  DFF_X1 \registers_reg[42][25]  ( .D(n9651), .CK(clk), .Q(\registers[42][25] ), .QN(n15952) );
  DFF_X1 \registers_reg[43][25]  ( .D(n9650), .CK(clk), .Q(\registers[43][25] ), .QN(n14877) );
  DFF_X1 \registers_reg[44][25]  ( .D(n9649), .CK(clk), .Q(\registers[44][25] ), .QN(n15461) );
  DFF_X1 \registers_reg[45][25]  ( .D(n9648), .CK(clk), .Q(\registers[45][25] ), .QN(n14762) );
  DFF_X1 \registers_reg[46][25]  ( .D(n9647), .CK(clk), .QN(n11945) );
  DFF_X1 \registers_reg[47][25]  ( .D(n9646), .CK(clk), .Q(\registers[47][25] ), .QN(n14541) );
  DFF_X1 \registers_reg[48][25]  ( .D(n9645), .CK(clk), .Q(\registers[48][25] ), .QN(n15546) );
  DFF_X1 \registers_reg[49][25]  ( .D(n9644), .CK(clk), .Q(\registers[49][25] ), .QN(n14472) );
  DFF_X1 \registers_reg[50][25]  ( .D(n9643), .CK(clk), .Q(\registers[50][25] ), .QN(n15994) );
  DFF_X1 \registers_reg[51][25]  ( .D(n9642), .CK(clk), .Q(\registers[51][25] ), .QN(n15422) );
  DFF_X1 \registers_reg[52][25]  ( .D(n9641), .CK(clk), .Q(net227354), .QN(
        n14932) );
  DFF_X1 \registers_reg[53][25]  ( .D(n9640), .CK(clk), .Q(net227353), .QN(
        n15943) );
  DFF_X1 \registers_reg[54][25]  ( .D(n9639), .CK(clk), .Q(\registers[54][25] ), .QN(n14593) );
  DFF_X1 \registers_reg[55][25]  ( .D(n9638), .CK(clk), .Q(\registers[55][25] ), .QN(n12155) );
  DFF_X1 \registers_reg[56][25]  ( .D(n9637), .CK(clk), .Q(\registers[56][25] ), .QN(n16008) );
  DFF_X1 \registers_reg[57][25]  ( .D(n9636), .CK(clk), .Q(net227352), .QN(
        n15265) );
  DFF_X1 \registers_reg[58][25]  ( .D(n9635), .CK(clk), .Q(net227351), .QN(
        n14878) );
  DFF_X1 \registers_reg[59][25]  ( .D(n9634), .CK(clk), .Q(\registers[59][25] ), .QN(n15520) );
  DFF_X1 \registers_reg[60][25]  ( .D(n9633), .CK(clk), .Q(\registers[60][25] ), .QN(n14665) );
  DFF_X1 \registers_reg[61][25]  ( .D(n9632), .CK(clk), .Q(net227350), .QN(
        n15656) );
  DFF_X1 \registers_reg[62][25]  ( .D(n9631), .CK(clk), .Q(\registers[62][25] ), .QN(n15118) );
  DFF_X1 \registers_reg[63][25]  ( .D(n9630), .CK(clk), .Q(\registers[63][25] ), .QN(n14479) );
  DFF_X1 \to_mem_reg[25]  ( .D(n9629), .CK(clk), .QN(n7700) );
  DFF_X1 \registers_reg[64][25]  ( .D(n9628), .CK(clk), .Q(net227349), .QN(
        n16144) );
  DFF_X1 \registers_reg[65][25]  ( .D(n9627), .CK(clk), .Q(net227348), .QN(
        n16093) );
  DFF_X1 \registers_reg[66][25]  ( .D(n9626), .CK(clk), .Q(net227347), .QN(
        n16055) );
  DFF_X1 \registers_reg[67][25]  ( .D(n9625), .CK(clk), .QN(n14274) );
  DFF_X1 \registers_reg[68][25]  ( .D(n9624), .CK(clk), .Q(\registers[68][25] ), .QN(n16181) );
  DFF_X1 \registers_reg[69][25]  ( .D(n9623), .CK(clk), .Q(net227346), .QN(
        n16133) );
  DFF_X1 \registers_reg[70][25]  ( .D(n9622), .CK(clk), .Q(net227345), .QN(
        n16045) );
  DFF_X1 \registers_reg[0][24]  ( .D(n9621), .CK(clk), .Q(\registers[0][24] ), 
        .QN(n15875) );
  DFF_X1 \registers_reg[1][24]  ( .D(n9620), .CK(clk), .Q(\registers[1][24] ), 
        .QN(n15632) );
  DFF_X1 \registers_reg[2][24]  ( .D(n9619), .CK(clk), .Q(\registers[2][24] ), 
        .QN(n14759) );
  DFF_X1 \registers_reg[3][24]  ( .D(n9618), .CK(clk), .Q(net227344), .QN(
        n15725) );
  DFF_X1 \registers_reg[4][24]  ( .D(n9617), .CK(clk), .Q(\registers[4][24] ), 
        .QN(n15452) );
  DFF_X1 \registers_reg[5][24]  ( .D(n9616), .CK(clk), .Q(\registers[5][24] ), 
        .QN(n14818) );
  DFF_X1 \registers_reg[6][24]  ( .D(n9615), .CK(clk), .QN(n12342) );
  DFF_X1 \registers_reg[7][24]  ( .D(n9614), .CK(clk), .Q(\registers[7][24] ), 
        .QN(n15320) );
  DFF_X1 \registers_reg[8][24]  ( .D(n9613), .CK(clk), .Q(net227343), .QN(
        n15233) );
  DFF_X1 \registers_reg[9][24]  ( .D(n9612), .CK(clk), .Q(\registers[9][24] ), 
        .QN(n14352) );
  DFF_X1 \registers_reg[10][24]  ( .D(n9611), .CK(clk), .Q(\registers[10][24] ), .QN(n14701) );
  DFF_X1 \registers_reg[11][24]  ( .D(n9610), .CK(clk), .Q(\registers[11][24] ), .QN(n14419) );
  DFF_X1 \registers_reg[12][24]  ( .D(n9609), .CK(clk), .Q(\registers[12][24] ), .QN(n15663) );
  DFF_X1 \registers_reg[13][24]  ( .D(n9608), .CK(clk), .Q(net227342), .QN(
        n15065) );
  DFF_X1 \registers_reg[14][24]  ( .D(n9607), .CK(clk), .QN(n11875) );
  DFF_X1 \registers_reg[15][24]  ( .D(n9606), .CK(clk), .Q(\registers[15][24] ), .QN(n15286) );
  DFF_X1 \registers_reg[16][24]  ( .D(n9605), .CK(clk), .Q(\registers[16][24] ), .QN(n15693) );
  DFF_X1 \registers_reg[17][24]  ( .D(n9604), .CK(clk), .Q(\registers[17][24] ), .QN(n14599) );
  DFF_X1 \registers_reg[18][24]  ( .D(n9603), .CK(clk), .Q(\registers[18][24] ), .QN(n14414) );
  DFF_X1 \registers_reg[19][24]  ( .D(n9602), .CK(clk), .Q(\registers[19][24] ), .QN(n15853) );
  DFF_X1 \registers_reg[20][24]  ( .D(n9601), .CK(clk), .QN(n14825) );
  DFF_X1 \registers_reg[21][24]  ( .D(n9600), .CK(clk), .QN(n12199) );
  DFF_X1 \registers_reg[22][24]  ( .D(n9599), .CK(clk), .Q(\registers[22][24] ), .QN(n15396) );
  DFF_X1 \registers_reg[23][24]  ( .D(n9598), .CK(clk), .Q(\registers[23][24] ), .QN(n15906) );
  DFF_X1 \registers_reg[24][24]  ( .D(n9597), .CK(clk), .Q(net227341), .QN(
        n15203) );
  DFF_X1 \registers_reg[25][24]  ( .D(n9596), .CK(clk), .Q(\registers[25][24] ), .QN(n14322) );
  DFF_X1 \registers_reg[26][24]  ( .D(n9595), .CK(clk), .QN(n12349) );
  DFF_X1 \registers_reg[27][24]  ( .D(n9594), .CK(clk), .QN(n12041) );
  DFF_X1 \registers_reg[28][24]  ( .D(n9593), .CK(clk), .Q(net227340), .QN(
        n15026) );
  DFF_X1 \registers_reg[29][24]  ( .D(n9592), .CK(clk), .Q(\registers[29][24] ), .QN(n15844) );
  DFF_X1 \registers_reg[30][24]  ( .D(n9591), .CK(clk), .Q(\registers[30][24] ), .QN(n14672) );
  DFF_X1 \registers_reg[31][24]  ( .D(n9590), .CK(clk), .Q(net227339), .QN(
        n15724) );
  DFF_X1 \registers_reg[32][24]  ( .D(n9589), .CK(clk), .QN(n12333) );
  DFF_X1 \registers_reg[33][24]  ( .D(n9588), .CK(clk), .QN(n11869) );
  DFF_X1 \registers_reg[34][24]  ( .D(n9587), .CK(clk), .Q(\registers[34][24] ), .QN(n15489) );
  DFF_X1 \registers_reg[35][24]  ( .D(n9586), .CK(clk), .Q(net227338), .QN(
        n15621) );
  DFF_X1 \registers_reg[36][24]  ( .D(n9585), .CK(clk), .Q(\registers[36][24] ), .QN(n15176) );
  DFF_X1 \registers_reg[37][24]  ( .D(n9584), .CK(clk), .Q(\registers[37][24] ), .QN(n14403) );
  DFF_X1 \registers_reg[38][24]  ( .D(n9583), .CK(clk), .Q(\registers[38][24] ), .QN(n15060) );
  DFF_X1 \registers_reg[39][24]  ( .D(n9582), .CK(clk), .QN(n12165) );
  DFF_X1 \registers_reg[40][24]  ( .D(n9581), .CK(clk), .Q(\registers[40][24] ), .QN(n15144) );
  DFF_X1 \registers_reg[41][24]  ( .D(n9580), .CK(clk), .Q(\registers[41][24] ), .QN(n14527) );
  DFF_X1 \registers_reg[42][24]  ( .D(n9579), .CK(clk), .Q(\registers[42][24] ), .QN(n15951) );
  DFF_X1 \registers_reg[43][24]  ( .D(n9578), .CK(clk), .Q(\registers[43][24] ), .QN(n14875) );
  DFF_X1 \registers_reg[44][24]  ( .D(n9577), .CK(clk), .Q(\registers[44][24] ), .QN(n15460) );
  DFF_X1 \registers_reg[45][24]  ( .D(n9576), .CK(clk), .Q(\registers[45][24] ), .QN(n14760) );
  DFF_X1 \registers_reg[46][24]  ( .D(n9575), .CK(clk), .QN(n11907) );
  DFF_X1 \registers_reg[47][24]  ( .D(n9574), .CK(clk), .Q(\registers[47][24] ), .QN(n14540) );
  DFF_X1 \registers_reg[48][24]  ( .D(n9573), .CK(clk), .Q(\registers[48][24] ), .QN(n15545) );
  DFF_X1 \registers_reg[49][24]  ( .D(n9572), .CK(clk), .Q(\registers[49][24] ), .QN(n14471) );
  DFF_X1 \registers_reg[50][24]  ( .D(n9571), .CK(clk), .Q(\registers[50][24] ), .QN(n15993) );
  DFF_X1 \registers_reg[51][24]  ( .D(n9570), .CK(clk), .Q(\registers[51][24] ), .QN(n15421) );
  DFF_X1 \registers_reg[52][24]  ( .D(n9569), .CK(clk), .Q(net227336), .QN(
        n14931) );
  DFF_X1 \registers_reg[53][24]  ( .D(n9568), .CK(clk), .Q(net227335), .QN(
        n15942) );
  DFF_X1 \registers_reg[54][24]  ( .D(n9567), .CK(clk), .Q(\registers[54][24] ), .QN(n14592) );
  DFF_X1 \registers_reg[55][24]  ( .D(n9566), .CK(clk), .Q(\registers[55][24] ), .QN(n12154) );
  DFF_X1 \registers_reg[56][24]  ( .D(n9565), .CK(clk), .Q(\registers[56][24] ), .QN(n16007) );
  DFF_X1 \registers_reg[57][24]  ( .D(n9564), .CK(clk), .Q(net227334), .QN(
        n15264) );
  DFF_X1 \registers_reg[58][24]  ( .D(n9563), .CK(clk), .Q(net227333), .QN(
        n14876) );
  DFF_X1 \registers_reg[59][24]  ( .D(n9562), .CK(clk), .Q(\registers[59][24] ), .QN(n15519) );
  DFF_X1 \registers_reg[60][24]  ( .D(n9561), .CK(clk), .Q(\registers[60][24] ), .QN(n14664) );
  DFF_X1 \registers_reg[61][24]  ( .D(n9560), .CK(clk), .Q(net227332), .QN(
        n15655) );
  DFF_X1 \registers_reg[62][24]  ( .D(n9559), .CK(clk), .Q(\registers[62][24] ), .QN(n15117) );
  DFF_X1 \registers_reg[63][24]  ( .D(n9558), .CK(clk), .Q(\registers[63][24] ), .QN(n14478) );
  DFF_X1 \to_mem_reg[24]  ( .D(n9557), .CK(clk), .QN(n7701) );
  DFF_X1 \registers_reg[64][24]  ( .D(n9556), .CK(clk), .Q(net227331), .QN(
        n16143) );
  DFF_X1 \registers_reg[65][24]  ( .D(n9555), .CK(clk), .Q(net227330), .QN(
        n16092) );
  DFF_X1 \registers_reg[66][24]  ( .D(n9554), .CK(clk), .Q(net227329), .QN(
        n16054) );
  DFF_X1 \registers_reg[67][24]  ( .D(n9553), .CK(clk), .QN(n14273) );
  DFF_X1 \registers_reg[68][24]  ( .D(n9552), .CK(clk), .Q(\registers[68][24] ), .QN(n16180) );
  DFF_X1 \registers_reg[69][24]  ( .D(n9551), .CK(clk), .Q(net227328), .QN(
        n16132) );
  DFF_X1 \registers_reg[70][24]  ( .D(n9550), .CK(clk), .Q(net227327), .QN(
        n16044) );
  DFF_X1 \registers_reg[0][23]  ( .D(n9549), .CK(clk), .Q(\registers[0][23] ), 
        .QN(n15874) );
  DFF_X1 \registers_reg[1][23]  ( .D(n9548), .CK(clk), .Q(\registers[1][23] ), 
        .QN(n15631) );
  DFF_X1 \registers_reg[2][23]  ( .D(n9547), .CK(clk), .Q(\registers[2][23] ), 
        .QN(n14757) );
  DFF_X1 \registers_reg[3][23]  ( .D(n9546), .CK(clk), .Q(net227326), .QN(
        n15723) );
  DFF_X1 \registers_reg[4][23]  ( .D(n9545), .CK(clk), .Q(\registers[4][23] ), 
        .QN(n15544) );
  DFF_X1 \registers_reg[5][23]  ( .D(n9544), .CK(clk), .Q(\registers[5][23] ), 
        .QN(n14817) );
  DFF_X1 \registers_reg[6][23]  ( .D(n9543), .CK(clk), .QN(n14050) );
  DFF_X1 \registers_reg[7][23]  ( .D(n9542), .CK(clk), .Q(\registers[7][23] ), 
        .QN(n15319) );
  DFF_X1 \registers_reg[8][23]  ( .D(n9541), .CK(clk), .Q(net227325), .QN(
        n15232) );
  DFF_X1 \registers_reg[9][23]  ( .D(n9540), .CK(clk), .Q(\registers[9][23] ), 
        .QN(n14351) );
  DFF_X1 \registers_reg[10][23]  ( .D(n9539), .CK(clk), .Q(\registers[10][23] ), .QN(n14700) );
  DFF_X1 \registers_reg[11][23]  ( .D(n9538), .CK(clk), .Q(\registers[11][23] ), .QN(n14469) );
  DFF_X1 \registers_reg[12][23]  ( .D(n9537), .CK(clk), .Q(\registers[12][23] ), .QN(n15662) );
  DFF_X1 \registers_reg[13][23]  ( .D(n9536), .CK(clk), .Q(net227324), .QN(
        n15115) );
  DFF_X1 \registers_reg[14][23]  ( .D(n9535), .CK(clk), .QN(n11874) );
  DFF_X1 \registers_reg[15][23]  ( .D(n9534), .CK(clk), .Q(\registers[15][23] ), .QN(n15285) );
  DFF_X1 \registers_reg[16][23]  ( .D(n9533), .CK(clk), .Q(\registers[16][23] ), .QN(n15692) );
  DFF_X1 \registers_reg[17][23]  ( .D(n9532), .CK(clk), .Q(\registers[17][23] ), .QN(n14598) );
  DFF_X1 \registers_reg[18][23]  ( .D(n9531), .CK(clk), .Q(\registers[18][23] ), .QN(n14413) );
  DFF_X1 \registers_reg[19][23]  ( .D(n9530), .CK(clk), .Q(\registers[19][23] ), .QN(n15852) );
  DFF_X1 \registers_reg[20][23]  ( .D(n9529), .CK(clk), .QN(n14824) );
  DFF_X1 \registers_reg[21][23]  ( .D(n9528), .CK(clk), .QN(n12198) );
  DFF_X1 \registers_reg[22][23]  ( .D(n9527), .CK(clk), .Q(\registers[22][23] ), .QN(n15395) );
  DFF_X1 \registers_reg[23][23]  ( .D(n9526), .CK(clk), .Q(\registers[23][23] ), .QN(n15905) );
  DFF_X1 \registers_reg[24][23]  ( .D(n9525), .CK(clk), .Q(net227323), .QN(
        n15202) );
  DFF_X1 \registers_reg[25][23]  ( .D(n9524), .CK(clk), .Q(\registers[25][23] ), .QN(n14321) );
  DFF_X1 \registers_reg[26][23]  ( .D(n9523), .CK(clk), .QN(n14049) );
  DFF_X1 \registers_reg[27][23]  ( .D(n9522), .CK(clk), .QN(n12040) );
  DFF_X1 \registers_reg[28][23]  ( .D(n9521), .CK(clk), .Q(net227322), .QN(
        n15025) );
  DFF_X1 \registers_reg[29][23]  ( .D(n9520), .CK(clk), .Q(\registers[29][23] ), .QN(n15843) );
  DFF_X1 \registers_reg[30][23]  ( .D(n9519), .CK(clk), .Q(\registers[30][23] ), .QN(n14671) );
  DFF_X1 \registers_reg[31][23]  ( .D(n9518), .CK(clk), .Q(net227321), .QN(
        n15722) );
  DFF_X1 \registers_reg[32][23]  ( .D(n9517), .CK(clk), .QN(n12332) );
  DFF_X1 \registers_reg[33][23]  ( .D(n9516), .CK(clk), .QN(n11867) );
  DFF_X1 \registers_reg[34][23]  ( .D(n9515), .CK(clk), .Q(\registers[34][23] ), .QN(n15488) );
  DFF_X1 \registers_reg[35][23]  ( .D(n9514), .CK(clk), .Q(net227320), .QN(
        n15620) );
  DFF_X1 \registers_reg[36][23]  ( .D(n9513), .CK(clk), .Q(\registers[36][23] ), .QN(n15175) );
  DFF_X1 \registers_reg[37][23]  ( .D(n9512), .CK(clk), .Q(\registers[37][23] ), .QN(n14402) );
  DFF_X1 \registers_reg[38][23]  ( .D(n9511), .CK(clk), .Q(\registers[38][23] ), .QN(n15059) );
  DFF_X1 \registers_reg[39][23]  ( .D(n9510), .CK(clk), .QN(n12164) );
  DFF_X1 \registers_reg[40][23]  ( .D(n9509), .CK(clk), .Q(\registers[40][23] ), .QN(n15116) );
  DFF_X1 \registers_reg[41][23]  ( .D(n9508), .CK(clk), .Q(\registers[41][23] ), .QN(n14470) );
  DFF_X1 \registers_reg[42][23]  ( .D(n9507), .CK(clk), .Q(\registers[42][23] ), .QN(n15950) );
  DFF_X1 \registers_reg[43][23]  ( .D(n9506), .CK(clk), .Q(\registers[43][23] ), .QN(n14909) );
  DFF_X1 \registers_reg[44][23]  ( .D(n9505), .CK(clk), .Q(\registers[44][23] ), .QN(n15459) );
  DFF_X1 \registers_reg[45][23]  ( .D(n9504), .CK(clk), .Q(\registers[45][23] ), .QN(n14758) );
  DFF_X1 \registers_reg[46][23]  ( .D(n9503), .CK(clk), .QN(n12015) );
  DFF_X1 \registers_reg[47][23]  ( .D(n9502), .CK(clk), .Q(\registers[47][23] ), .QN(n14568) );
  DFF_X1 \registers_reg[48][23]  ( .D(n9501), .CK(clk), .Q(\registers[48][23] ), .QN(n15573) );
  DFF_X1 \registers_reg[49][23]  ( .D(n9500), .CK(clk), .Q(\registers[49][23] ), .QN(n14505) );
  DFF_X1 \registers_reg[50][23]  ( .D(n9499), .CK(clk), .Q(\registers[50][23] ), .QN(n15992) );
  DFF_X1 \registers_reg[51][23]  ( .D(n9498), .CK(clk), .Q(\registers[51][23] ), .QN(n15420) );
  DFF_X1 \registers_reg[52][23]  ( .D(n9497), .CK(clk), .Q(net227318), .QN(
        n14959) );
  DFF_X1 \registers_reg[53][23]  ( .D(n9496), .CK(clk), .Q(net227317), .QN(
        n15941) );
  DFF_X1 \registers_reg[54][23]  ( .D(n9495), .CK(clk), .Q(\registers[54][23] ), .QN(n14591) );
  DFF_X1 \registers_reg[55][23]  ( .D(n9494), .CK(clk), .Q(\registers[55][23] ), .QN(n12153) );
  DFF_X1 \registers_reg[56][23]  ( .D(n9493), .CK(clk), .Q(\registers[56][23] ), .QN(n16006) );
  DFF_X1 \registers_reg[57][23]  ( .D(n9492), .CK(clk), .Q(net227316), .QN(
        n15263) );
  DFF_X1 \registers_reg[58][23]  ( .D(n9491), .CK(clk), .Q(net227315), .QN(
        n14930) );
  DFF_X1 \registers_reg[59][23]  ( .D(n9490), .CK(clk), .Q(\registers[59][23] ), .QN(n15518) );
  DFF_X1 \registers_reg[60][23]  ( .D(n9489), .CK(clk), .Q(\registers[60][23] ), .QN(n14663) );
  DFF_X1 \registers_reg[61][23]  ( .D(n9488), .CK(clk), .Q(net227314), .QN(
        n15654) );
  DFF_X1 \registers_reg[62][23]  ( .D(n9487), .CK(clk), .Q(\registers[62][23] ), .QN(n15143) );
  DFF_X1 \registers_reg[63][23]  ( .D(n9486), .CK(clk), .Q(\registers[63][23] ), .QN(n14526) );
  DFF_X1 \to_mem_reg[23]  ( .D(n9485), .CK(clk), .QN(n7702) );
  DFF_X1 \registers_reg[64][23]  ( .D(n9484), .CK(clk), .Q(net227313), .QN(
        n16142) );
  DFF_X1 \registers_reg[65][23]  ( .D(n9483), .CK(clk), .Q(net227312), .QN(
        n16091) );
  DFF_X1 \registers_reg[66][23]  ( .D(n9482), .CK(clk), .Q(net227311), .QN(
        n16053) );
  DFF_X1 \registers_reg[67][23]  ( .D(n9481), .CK(clk), .QN(n14272) );
  DFF_X1 \registers_reg[68][23]  ( .D(n9480), .CK(clk), .Q(\registers[68][23] ), .QN(n16179) );
  DFF_X1 \registers_reg[69][23]  ( .D(n9479), .CK(clk), .Q(net227310), .QN(
        n16131) );
  DFF_X1 \registers_reg[70][23]  ( .D(n9478), .CK(clk), .Q(net227309), .QN(
        n16043) );
  DFF_X1 \registers_reg[0][22]  ( .D(n9477), .CK(clk), .Q(\registers[0][22] ), 
        .QN(n15873) );
  DFF_X1 \registers_reg[1][22]  ( .D(n9476), .CK(clk), .Q(\registers[1][22] ), 
        .QN(n15630) );
  DFF_X1 \registers_reg[2][22]  ( .D(n9475), .CK(clk), .Q(\registers[2][22] ), 
        .QN(n14813) );
  DFF_X1 \registers_reg[3][22]  ( .D(n9474), .CK(clk), .Q(net227308), .QN(
        n15780) );
  DFF_X1 \registers_reg[4][22]  ( .D(n9473), .CK(clk), .Q(\registers[4][22] ), 
        .QN(n15543) );
  DFF_X1 \registers_reg[5][22]  ( .D(n9472), .CK(clk), .Q(\registers[5][22] ), 
        .QN(n14754) );
  DFF_X1 \registers_reg[6][22]  ( .D(n9471), .CK(clk), .QN(n14048) );
  DFF_X1 \registers_reg[7][22]  ( .D(n9470), .CK(clk), .Q(\registers[7][22] ), 
        .QN(n15348) );
  DFF_X1 \registers_reg[8][22]  ( .D(n9469), .CK(clk), .Q(net227307), .QN(
        n15231) );
  DFF_X1 \registers_reg[9][22]  ( .D(n9468), .CK(clk), .Q(\registers[9][22] ), 
        .QN(n14350) );
  DFF_X1 \registers_reg[10][22]  ( .D(n9467), .CK(clk), .Q(\registers[10][22] ), .QN(n14755) );
  DFF_X1 \registers_reg[11][22]  ( .D(n9466), .CK(clk), .Q(\registers[11][22] ), .QN(n14467) );
  DFF_X1 \registers_reg[12][22]  ( .D(n9465), .CK(clk), .Q(\registers[12][22] ), .QN(n15690) );
  DFF_X1 \registers_reg[13][22]  ( .D(n9464), .CK(clk), .Q(net227306), .QN(
        n15113) );
  DFF_X1 \registers_reg[14][22]  ( .D(n9463), .CK(clk), .QN(n11902) );
  DFF_X1 \registers_reg[15][22]  ( .D(n9462), .CK(clk), .Q(\registers[15][22] ), .QN(n15313) );
  DFF_X1 \registers_reg[16][22]  ( .D(n9461), .CK(clk), .Q(\registers[16][22] ), .QN(n15720) );
  DFF_X1 \registers_reg[17][22]  ( .D(n9460), .CK(clk), .Q(\registers[17][22] ), .QN(n14626) );
  DFF_X1 \registers_reg[18][22]  ( .D(n9459), .CK(clk), .Q(\registers[18][22] ), .QN(n14412) );
  DFF_X1 \registers_reg[19][22]  ( .D(n9458), .CK(clk), .Q(\registers[19][22] ), .QN(n15851) );
  DFF_X1 \registers_reg[20][22]  ( .D(n9457), .CK(clk), .QN(n14852) );
  DFF_X1 \registers_reg[21][22]  ( .D(n9456), .CK(clk), .QN(n12306) );
  DFF_X1 \registers_reg[22][22]  ( .D(n9455), .CK(clk), .Q(\registers[22][22] ), .QN(n15394) );
  DFF_X1 \registers_reg[23][22]  ( .D(n9454), .CK(clk), .Q(\registers[23][22] ), .QN(n15904) );
  DFF_X1 \registers_reg[24][22]  ( .D(n9453), .CK(clk), .Q(net227305), .QN(
        n15201) );
  DFF_X1 \registers_reg[25][22]  ( .D(n9452), .CK(clk), .Q(\registers[25][22] ), .QN(n14320) );
  DFF_X1 \registers_reg[26][22]  ( .D(n9451), .CK(clk), .QN(n14047) );
  DFF_X1 \registers_reg[27][22]  ( .D(n9450), .CK(clk), .QN(n12039) );
  DFF_X1 \registers_reg[28][22]  ( .D(n9449), .CK(clk), .Q(net227304), .QN(
        n15024) );
  DFF_X1 \registers_reg[29][22]  ( .D(n9448), .CK(clk), .Q(\registers[29][22] ), .QN(n15842) );
  DFF_X1 \registers_reg[30][22]  ( .D(n9447), .CK(clk), .Q(\registers[30][22] ), .QN(n14698) );
  DFF_X1 \registers_reg[31][22]  ( .D(n9446), .CK(clk), .Q(net227303), .QN(
        n15756) );
  DFF_X1 \registers_reg[32][22]  ( .D(n9445), .CK(clk), .QN(n12331) );
  DFF_X1 \registers_reg[33][22]  ( .D(n9444), .CK(clk), .QN(n11866) );
  DFF_X1 \registers_reg[34][22]  ( .D(n9443), .CK(clk), .Q(\registers[34][22] ), .QN(n15516) );
  DFF_X1 \registers_reg[35][22]  ( .D(n9442), .CK(clk), .Q(net227302), .QN(
        n15619) );
  DFF_X1 \registers_reg[36][22]  ( .D(n9441), .CK(clk), .Q(\registers[36][22] ), .QN(n15174) );
  DFF_X1 \registers_reg[37][22]  ( .D(n9440), .CK(clk), .Q(\registers[37][22] ), .QN(n14401) );
  DFF_X1 \registers_reg[38][22]  ( .D(n9439), .CK(clk), .Q(\registers[38][22] ), .QN(n15058) );
  DFF_X1 \registers_reg[39][22]  ( .D(n9438), .CK(clk), .QN(n12193) );
  DFF_X1 \registers_reg[40][22]  ( .D(n9437), .CK(clk), .Q(\registers[40][22] ), .QN(n15114) );
  DFF_X1 \registers_reg[41][22]  ( .D(n9436), .CK(clk), .Q(\registers[41][22] ), .QN(n14468) );
  DFF_X1 \registers_reg[42][22]  ( .D(n9435), .CK(clk), .Q(\registers[42][22] ), .QN(n15949) );
  DFF_X1 \registers_reg[43][22]  ( .D(n9434), .CK(clk), .Q(\registers[43][22] ), .QN(n14908) );
  DFF_X1 \registers_reg[44][22]  ( .D(n9433), .CK(clk), .Q(\registers[44][22] ), .QN(n15486) );
  DFF_X1 \registers_reg[45][22]  ( .D(n9432), .CK(clk), .Q(\registers[45][22] ), .QN(n14814) );
  DFF_X1 \registers_reg[46][22]  ( .D(n9431), .CK(clk), .QN(n12014) );
  DFF_X1 \registers_reg[47][22]  ( .D(n9430), .CK(clk), .Q(\registers[47][22] ), .QN(n14567) );
  DFF_X1 \registers_reg[48][22]  ( .D(n9429), .CK(clk), .Q(\registers[48][22] ), .QN(n15572) );
  DFF_X1 \registers_reg[49][22]  ( .D(n9428), .CK(clk), .Q(\registers[49][22] ), .QN(n14504) );
  DFF_X1 \registers_reg[50][22]  ( .D(n9427), .CK(clk), .Q(\registers[50][22] ), .QN(n15991) );
  DFF_X1 \registers_reg[51][22]  ( .D(n9426), .CK(clk), .Q(\registers[51][22] ), .QN(n15419) );
  DFF_X1 \registers_reg[52][22]  ( .D(n9425), .CK(clk), .Q(net227300), .QN(
        n14958) );
  DFF_X1 \registers_reg[53][22]  ( .D(n9424), .CK(clk), .Q(net227299), .QN(
        n15940) );
  DFF_X1 \registers_reg[54][22]  ( .D(n9423), .CK(clk), .Q(\registers[54][22] ), .QN(n14590) );
  DFF_X1 \registers_reg[55][22]  ( .D(n9422), .CK(clk), .Q(\registers[55][22] ), .QN(n12152) );
  DFF_X1 \registers_reg[56][22]  ( .D(n9421), .CK(clk), .Q(\registers[56][22] ), .QN(n16024) );
  DFF_X1 \registers_reg[57][22]  ( .D(n9420), .CK(clk), .Q(net227298), .QN(
        n15262) );
  DFF_X1 \registers_reg[58][22]  ( .D(n9419), .CK(clk), .Q(net227297), .QN(
        n14929) );
  DFF_X1 \registers_reg[59][22]  ( .D(n9418), .CK(clk), .Q(\registers[59][22] ), .QN(n15451) );
  DFF_X1 \registers_reg[60][22]  ( .D(n9417), .CK(clk), .Q(\registers[60][22] ), .QN(n14662) );
  DFF_X1 \registers_reg[61][22]  ( .D(n9416), .CK(clk), .Q(net227296), .QN(
        n15653) );
  DFF_X1 \registers_reg[62][22]  ( .D(n9415), .CK(clk), .Q(\registers[62][22] ), .QN(n15142) );
  DFF_X1 \registers_reg[63][22]  ( .D(n9414), .CK(clk), .Q(\registers[63][22] ), .QN(n14525) );
  DFF_X1 \to_mem_reg[22]  ( .D(n9413), .CK(clk), .QN(n7703) );
  DFF_X1 \registers_reg[64][22]  ( .D(n9412), .CK(clk), .Q(net227295), .QN(
        n16160) );
  DFF_X1 \registers_reg[65][22]  ( .D(n9411), .CK(clk), .Q(net227294), .QN(
        n16110) );
  DFF_X1 \registers_reg[66][22]  ( .D(n9410), .CK(clk), .Q(net227293), .QN(
        n16084) );
  DFF_X1 \registers_reg[67][22]  ( .D(n9409), .CK(clk), .QN(n14268) );
  DFF_X1 \registers_reg[68][22]  ( .D(n9408), .CK(clk), .Q(\registers[68][22] ), .QN(n16198) );
  DFF_X1 \registers_reg[69][22]  ( .D(n9407), .CK(clk), .Q(net227292), .QN(
        n16173) );
  DFF_X1 \registers_reg[70][22]  ( .D(n9406), .CK(clk), .Q(net227291), .QN(
        n16083) );
  DFF_X1 \registers_reg[0][21]  ( .D(n9405), .CK(clk), .Q(\registers[0][21] ), 
        .QN(n15872) );
  DFF_X1 \registers_reg[1][21]  ( .D(n9404), .CK(clk), .Q(\registers[1][21] ), 
        .QN(n15629) );
  DFF_X1 \registers_reg[2][21]  ( .D(n9403), .CK(clk), .Q(\registers[2][21] ), 
        .QN(n14811) );
  DFF_X1 \registers_reg[3][21]  ( .D(n9402), .CK(clk), .Q(net227290), .QN(
        n15779) );
  DFF_X1 \registers_reg[4][21]  ( .D(n9401), .CK(clk), .Q(\registers[4][21] ), 
        .QN(n15542) );
  DFF_X1 \registers_reg[5][21]  ( .D(n9400), .CK(clk), .Q(\registers[5][21] ), 
        .QN(n14752) );
  DFF_X1 \registers_reg[6][21]  ( .D(n9399), .CK(clk), .QN(n14046) );
  DFF_X1 \registers_reg[7][21]  ( .D(n9398), .CK(clk), .Q(\registers[7][21] ), 
        .QN(n15347) );
  DFF_X1 \registers_reg[8][21]  ( .D(n9397), .CK(clk), .Q(net227289), .QN(
        n15230) );
  DFF_X1 \registers_reg[9][21]  ( .D(n9396), .CK(clk), .Q(\registers[9][21] ), 
        .QN(n14349) );
  DFF_X1 \registers_reg[10][21]  ( .D(n9395), .CK(clk), .Q(\registers[10][21] ), .QN(n14753) );
  DFF_X1 \registers_reg[11][21]  ( .D(n9394), .CK(clk), .Q(\registers[11][21] ), .QN(n14465) );
  DFF_X1 \registers_reg[12][21]  ( .D(n9393), .CK(clk), .Q(\registers[12][21] ), .QN(n15689) );
  DFF_X1 \registers_reg[13][21]  ( .D(n9392), .CK(clk), .Q(net227288), .QN(
        n15111) );
  DFF_X1 \registers_reg[14][21]  ( .D(n9391), .CK(clk), .QN(n11901) );
  DFF_X1 \registers_reg[15][21]  ( .D(n9390), .CK(clk), .Q(\registers[15][21] ), .QN(n15312) );
  DFF_X1 \registers_reg[16][21]  ( .D(n9389), .CK(clk), .Q(\registers[16][21] ), .QN(n15719) );
  DFF_X1 \registers_reg[17][21]  ( .D(n9388), .CK(clk), .Q(\registers[17][21] ), .QN(n14625) );
  DFF_X1 \registers_reg[18][21]  ( .D(n9387), .CK(clk), .Q(\registers[18][21] ), .QN(n14411) );
  DFF_X1 \registers_reg[19][21]  ( .D(n9386), .CK(clk), .Q(\registers[19][21] ), .QN(n15850) );
  DFF_X1 \registers_reg[20][21]  ( .D(n9385), .CK(clk), .QN(n14851) );
  DFF_X1 \registers_reg[21][21]  ( .D(n9384), .CK(clk), .QN(n12305) );
  DFF_X1 \registers_reg[22][21]  ( .D(n9383), .CK(clk), .Q(\registers[22][21] ), .QN(n15393) );
  DFF_X1 \registers_reg[23][21]  ( .D(n9382), .CK(clk), .Q(\registers[23][21] ), .QN(n15903) );
  DFF_X1 \registers_reg[24][21]  ( .D(n9381), .CK(clk), .Q(net227287), .QN(
        n15200) );
  DFF_X1 \registers_reg[25][21]  ( .D(n9380), .CK(clk), .Q(\registers[25][21] ), .QN(n14319) );
  DFF_X1 \registers_reg[26][21]  ( .D(n9379), .CK(clk), .QN(n14045) );
  DFF_X1 \registers_reg[27][21]  ( .D(n9378), .CK(clk), .QN(n12038) );
  DFF_X1 \registers_reg[28][21]  ( .D(n9377), .CK(clk), .Q(net227286), .QN(
        n15023) );
  DFF_X1 \registers_reg[29][21]  ( .D(n9376), .CK(clk), .Q(\registers[29][21] ), .QN(n15841) );
  DFF_X1 \registers_reg[30][21]  ( .D(n9375), .CK(clk), .Q(\registers[30][21] ), .QN(n14697) );
  DFF_X1 \registers_reg[31][21]  ( .D(n9374), .CK(clk), .Q(net227285), .QN(
        n15755) );
  DFF_X1 \registers_reg[32][21]  ( .D(n9373), .CK(clk), .QN(n12330) );
  DFF_X1 \registers_reg[33][21]  ( .D(n9372), .CK(clk), .QN(n11865) );
  DFF_X1 \registers_reg[34][21]  ( .D(n9371), .CK(clk), .Q(\registers[34][21] ), .QN(n15515) );
  DFF_X1 \registers_reg[35][21]  ( .D(n9370), .CK(clk), .Q(net227284), .QN(
        n15618) );
  DFF_X1 \registers_reg[36][21]  ( .D(n9369), .CK(clk), .Q(\registers[36][21] ), .QN(n15173) );
  DFF_X1 \registers_reg[37][21]  ( .D(n9368), .CK(clk), .Q(\registers[37][21] ), .QN(n14400) );
  DFF_X1 \registers_reg[38][21]  ( .D(n9367), .CK(clk), .Q(\registers[38][21] ), .QN(n15057) );
  DFF_X1 \registers_reg[39][21]  ( .D(n9366), .CK(clk), .QN(n12192) );
  DFF_X1 \registers_reg[40][21]  ( .D(n9365), .CK(clk), .Q(\registers[40][21] ), .QN(n15112) );
  DFF_X1 \registers_reg[41][21]  ( .D(n9364), .CK(clk), .Q(\registers[41][21] ), .QN(n14466) );
  DFF_X1 \registers_reg[42][21]  ( .D(n9363), .CK(clk), .Q(\registers[42][21] ), .QN(n15948) );
  DFF_X1 \registers_reg[43][21]  ( .D(n9362), .CK(clk), .Q(\registers[43][21] ), .QN(n14907) );
  DFF_X1 \registers_reg[44][21]  ( .D(n9361), .CK(clk), .Q(\registers[44][21] ), .QN(n15485) );
  DFF_X1 \registers_reg[45][21]  ( .D(n9360), .CK(clk), .Q(\registers[45][21] ), .QN(n14812) );
  DFF_X1 \registers_reg[46][21]  ( .D(n9359), .CK(clk), .QN(n12013) );
  DFF_X1 \registers_reg[47][21]  ( .D(n9358), .CK(clk), .Q(\registers[47][21] ), .QN(n14566) );
  DFF_X1 \registers_reg[48][21]  ( .D(n9357), .CK(clk), .Q(\registers[48][21] ), .QN(n15571) );
  DFF_X1 \registers_reg[49][21]  ( .D(n9356), .CK(clk), .Q(\registers[49][21] ), .QN(n14503) );
  DFF_X1 \registers_reg[50][21]  ( .D(n9355), .CK(clk), .Q(\registers[50][21] ), .QN(n15990) );
  DFF_X1 \registers_reg[51][21]  ( .D(n9354), .CK(clk), .Q(\registers[51][21] ), .QN(n15418) );
  DFF_X1 \registers_reg[52][21]  ( .D(n9353), .CK(clk), .Q(net227282), .QN(
        n14957) );
  DFF_X1 \registers_reg[53][21]  ( .D(n9352), .CK(clk), .Q(net227281), .QN(
        n15967) );
  DFF_X1 \registers_reg[54][21]  ( .D(n9351), .CK(clk), .Q(\registers[54][21] ), .QN(n14589) );
  DFF_X1 \registers_reg[55][21]  ( .D(n9350), .CK(clk), .Q(\registers[55][21] ), .QN(n12151) );
  DFF_X1 \registers_reg[56][21]  ( .D(n9349), .CK(clk), .Q(\registers[56][21] ), .QN(n16005) );
  DFF_X1 \registers_reg[57][21]  ( .D(n9348), .CK(clk), .Q(net227280), .QN(
        n15261) );
  DFF_X1 \registers_reg[58][21]  ( .D(n9347), .CK(clk), .Q(net227279), .QN(
        n14928) );
  DFF_X1 \registers_reg[59][21]  ( .D(n9346), .CK(clk), .Q(\registers[59][21] ), .QN(n15450) );
  DFF_X1 \registers_reg[60][21]  ( .D(n9345), .CK(clk), .Q(\registers[60][21] ), .QN(n14661) );
  DFF_X1 \registers_reg[61][21]  ( .D(n9344), .CK(clk), .Q(net227278), .QN(
        n15652) );
  DFF_X1 \registers_reg[62][21]  ( .D(n9343), .CK(clk), .Q(\registers[62][21] ), .QN(n15141) );
  DFF_X1 \registers_reg[63][21]  ( .D(n9342), .CK(clk), .Q(\registers[63][21] ), .QN(n14524) );
  DFF_X1 \to_mem_reg[21]  ( .D(n9341), .CK(clk), .QN(n7704) );
  DFF_X1 \registers_reg[64][21]  ( .D(n9340), .CK(clk), .Q(net227277), .QN(
        n16141) );
  DFF_X1 \registers_reg[65][21]  ( .D(n9339), .CK(clk), .Q(net227276), .QN(
        n16090) );
  DFF_X1 \registers_reg[66][21]  ( .D(n9338), .CK(clk), .Q(net227275), .QN(
        n16052) );
  DFF_X1 \registers_reg[67][21]  ( .D(n9337), .CK(clk), .QN(n14271) );
  DFF_X1 \registers_reg[68][21]  ( .D(n9336), .CK(clk), .Q(\registers[68][21] ), .QN(n16178) );
  DFF_X1 \registers_reg[69][21]  ( .D(n9335), .CK(clk), .Q(net227274), .QN(
        n16130) );
  DFF_X1 \registers_reg[70][21]  ( .D(n9334), .CK(clk), .Q(net227273), .QN(
        n16042) );
  DFF_X1 \registers_reg[0][20]  ( .D(n9333), .CK(clk), .Q(\registers[0][20] ), 
        .QN(n15871) );
  DFF_X1 \registers_reg[1][20]  ( .D(n9332), .CK(clk), .Q(\registers[1][20] ), 
        .QN(n15628) );
  DFF_X1 \registers_reg[2][20]  ( .D(n9331), .CK(clk), .Q(\registers[2][20] ), 
        .QN(n14809) );
  DFF_X1 \registers_reg[3][20]  ( .D(n9330), .CK(clk), .Q(net227272), .QN(
        n15778) );
  DFF_X1 \registers_reg[4][20]  ( .D(n9329), .CK(clk), .Q(\registers[4][20] ), 
        .QN(n15541) );
  DFF_X1 \registers_reg[5][20]  ( .D(n9328), .CK(clk), .Q(\registers[5][20] ), 
        .QN(n14750) );
  DFF_X1 \registers_reg[6][20]  ( .D(n9327), .CK(clk), .QN(n14044) );
  DFF_X1 \registers_reg[7][20]  ( .D(n9326), .CK(clk), .Q(\registers[7][20] ), 
        .QN(n15346) );
  DFF_X1 \registers_reg[8][20]  ( .D(n9325), .CK(clk), .Q(net227271), .QN(
        n15229) );
  DFF_X1 \registers_reg[9][20]  ( .D(n9324), .CK(clk), .Q(\registers[9][20] ), 
        .QN(n14348) );
  DFF_X1 \registers_reg[10][20]  ( .D(n9323), .CK(clk), .Q(\registers[10][20] ), .QN(n14751) );
  DFF_X1 \registers_reg[11][20]  ( .D(n9322), .CK(clk), .Q(\registers[11][20] ), .QN(n14463) );
  DFF_X1 \registers_reg[12][20]  ( .D(n9321), .CK(clk), .Q(\registers[12][20] ), .QN(n15688) );
  DFF_X1 \registers_reg[13][20]  ( .D(n9320), .CK(clk), .Q(net227270), .QN(
        n15109) );
  DFF_X1 \registers_reg[14][20]  ( .D(n9319), .CK(clk), .QN(n11900) );
  DFF_X1 \registers_reg[15][20]  ( .D(n9318), .CK(clk), .Q(\registers[15][20] ), .QN(n15311) );
  DFF_X1 \registers_reg[16][20]  ( .D(n9317), .CK(clk), .Q(\registers[16][20] ), .QN(n15718) );
  DFF_X1 \registers_reg[17][20]  ( .D(n9316), .CK(clk), .Q(\registers[17][20] ), .QN(n14624) );
  DFF_X1 \registers_reg[18][20]  ( .D(n9315), .CK(clk), .Q(\registers[18][20] ), .QN(n14410) );
  DFF_X1 \registers_reg[19][20]  ( .D(n9314), .CK(clk), .Q(\registers[19][20] ), .QN(n15849) );
  DFF_X1 \registers_reg[20][20]  ( .D(n9313), .CK(clk), .QN(n14850) );
  DFF_X1 \registers_reg[21][20]  ( .D(n9312), .CK(clk), .QN(n12304) );
  DFF_X1 \registers_reg[22][20]  ( .D(n9311), .CK(clk), .Q(\registers[22][20] ), .QN(n15392) );
  DFF_X1 \registers_reg[23][20]  ( .D(n9310), .CK(clk), .Q(\registers[23][20] ), .QN(n15901) );
  DFF_X1 \registers_reg[24][20]  ( .D(n9309), .CK(clk), .Q(net227269), .QN(
        n15199) );
  DFF_X1 \registers_reg[25][20]  ( .D(n9308), .CK(clk), .Q(\registers[25][20] ), .QN(n14318) );
  DFF_X1 \registers_reg[26][20]  ( .D(n9307), .CK(clk), .QN(n14043) );
  DFF_X1 \registers_reg[27][20]  ( .D(n9306), .CK(clk), .QN(n12037) );
  DFF_X1 \registers_reg[28][20]  ( .D(n9305), .CK(clk), .Q(net227268), .QN(
        n15022) );
  DFF_X1 \registers_reg[29][20]  ( .D(n9304), .CK(clk), .Q(\registers[29][20] ), .QN(n15838) );
  DFF_X1 \registers_reg[30][20]  ( .D(n9303), .CK(clk), .Q(\registers[30][20] ), .QN(n14696) );
  DFF_X1 \registers_reg[31][20]  ( .D(n9302), .CK(clk), .Q(net227267), .QN(
        n15754) );
  DFF_X1 \registers_reg[32][20]  ( .D(n9301), .CK(clk), .QN(n12329) );
  DFF_X1 \registers_reg[33][20]  ( .D(n9300), .CK(clk), .QN(n11864) );
  DFF_X1 \registers_reg[34][20]  ( .D(n9299), .CK(clk), .Q(\registers[34][20] ), .QN(n15514) );
  DFF_X1 \registers_reg[35][20]  ( .D(n9298), .CK(clk), .Q(net227266), .QN(
        n15617) );
  DFF_X1 \registers_reg[36][20]  ( .D(n9297), .CK(clk), .Q(\registers[36][20] ), .QN(n15172) );
  DFF_X1 \registers_reg[37][20]  ( .D(n9296), .CK(clk), .Q(\registers[37][20] ), .QN(n14399) );
  DFF_X1 \registers_reg[38][20]  ( .D(n9295), .CK(clk), .Q(\registers[38][20] ), .QN(n15056) );
  DFF_X1 \registers_reg[39][20]  ( .D(n9294), .CK(clk), .QN(n12191) );
  DFF_X1 \registers_reg[40][20]  ( .D(n9293), .CK(clk), .Q(\registers[40][20] ), .QN(n15110) );
  DFF_X1 \registers_reg[41][20]  ( .D(n9292), .CK(clk), .Q(\registers[41][20] ), .QN(n14464) );
  DFF_X1 \registers_reg[42][20]  ( .D(n9291), .CK(clk), .Q(\registers[42][20] ), .QN(n15947) );
  DFF_X1 \registers_reg[43][20]  ( .D(n9290), .CK(clk), .Q(\registers[43][20] ), .QN(n14906) );
  DFF_X1 \registers_reg[44][20]  ( .D(n9289), .CK(clk), .Q(\registers[44][20] ), .QN(n15484) );
  DFF_X1 \registers_reg[45][20]  ( .D(n9288), .CK(clk), .Q(\registers[45][20] ), .QN(n14810) );
  DFF_X1 \registers_reg[46][20]  ( .D(n9287), .CK(clk), .QN(n12012) );
  DFF_X1 \registers_reg[47][20]  ( .D(n9286), .CK(clk), .Q(\registers[47][20] ), .QN(n14565) );
  DFF_X1 \registers_reg[48][20]  ( .D(n9285), .CK(clk), .Q(\registers[48][20] ), .QN(n15570) );
  DFF_X1 \registers_reg[49][20]  ( .D(n9284), .CK(clk), .Q(\registers[49][20] ), .QN(n14502) );
  DFF_X1 \registers_reg[50][20]  ( .D(n9283), .CK(clk), .Q(\registers[50][20] ), .QN(n15989) );
  DFF_X1 \registers_reg[51][20]  ( .D(n9282), .CK(clk), .Q(\registers[51][20] ), .QN(n15417) );
  DFF_X1 \registers_reg[52][20]  ( .D(n9281), .CK(clk), .Q(net227264), .QN(
        n14956) );
  DFF_X1 \registers_reg[53][20]  ( .D(n9280), .CK(clk), .Q(net227263), .QN(
        n15966) );
  DFF_X1 \registers_reg[54][20]  ( .D(n9279), .CK(clk), .Q(\registers[54][20] ), .QN(n14588) );
  DFF_X1 \registers_reg[55][20]  ( .D(n9278), .CK(clk), .Q(\registers[55][20] ), .QN(n12150) );
  DFF_X1 \registers_reg[56][20]  ( .D(n9277), .CK(clk), .Q(\registers[56][20] ), .QN(n16004) );
  DFF_X1 \registers_reg[57][20]  ( .D(n9276), .CK(clk), .Q(net227262), .QN(
        n15260) );
  DFF_X1 \registers_reg[58][20]  ( .D(n9275), .CK(clk), .Q(net227261), .QN(
        n14927) );
  DFF_X1 \registers_reg[59][20]  ( .D(n9274), .CK(clk), .Q(\registers[59][20] ), .QN(n15449) );
  DFF_X1 \registers_reg[60][20]  ( .D(n9273), .CK(clk), .Q(\registers[60][20] ), .QN(n14660) );
  DFF_X1 \registers_reg[61][20]  ( .D(n9272), .CK(clk), .Q(net227260), .QN(
        n15651) );
  DFF_X1 \registers_reg[62][20]  ( .D(n9271), .CK(clk), .Q(\registers[62][20] ), .QN(n15140) );
  DFF_X1 \registers_reg[63][20]  ( .D(n9270), .CK(clk), .Q(\registers[63][20] ), .QN(n14523) );
  DFF_X1 \to_mem_reg[20]  ( .D(n9269), .CK(clk), .QN(n7705) );
  DFF_X1 \registers_reg[64][20]  ( .D(n9268), .CK(clk), .Q(net227259), .QN(
        n16140) );
  DFF_X1 \registers_reg[65][20]  ( .D(n9267), .CK(clk), .Q(net227258), .QN(
        n16089) );
  DFF_X1 \registers_reg[66][20]  ( .D(n9266), .CK(clk), .Q(net227257), .QN(
        n16051) );
  DFF_X1 \registers_reg[67][20]  ( .D(n9265), .CK(clk), .QN(n14270) );
  DFF_X1 \registers_reg[68][20]  ( .D(n9264), .CK(clk), .Q(\registers[68][20] ), .QN(n16177) );
  DFF_X1 \registers_reg[69][20]  ( .D(n9263), .CK(clk), .Q(net227256), .QN(
        n16129) );
  DFF_X1 \registers_reg[70][20]  ( .D(n9262), .CK(clk), .Q(net227255), .QN(
        n16082) );
  DFF_X1 \registers_reg[0][19]  ( .D(n9261), .CK(clk), .Q(\registers[0][19] ), 
        .QN(n15870) );
  DFF_X1 \registers_reg[1][19]  ( .D(n9260), .CK(clk), .Q(\registers[1][19] ), 
        .QN(n15627) );
  DFF_X1 \registers_reg[2][19]  ( .D(n9259), .CK(clk), .Q(\registers[2][19] ), 
        .QN(n14807) );
  DFF_X1 \registers_reg[3][19]  ( .D(n9258), .CK(clk), .Q(net227254), .QN(
        n15777) );
  DFF_X1 \registers_reg[4][19]  ( .D(n9257), .CK(clk), .Q(\registers[4][19] ), 
        .QN(n15540) );
  DFF_X1 \registers_reg[5][19]  ( .D(n9256), .CK(clk), .Q(\registers[5][19] ), 
        .QN(n14748) );
  DFF_X1 \registers_reg[6][19]  ( .D(n9255), .CK(clk), .QN(n14042) );
  DFF_X1 \registers_reg[7][19]  ( .D(n9254), .CK(clk), .Q(\registers[7][19] ), 
        .QN(n15345) );
  DFF_X1 \registers_reg[8][19]  ( .D(n9253), .CK(clk), .Q(net227253), .QN(
        n15228) );
  DFF_X1 \registers_reg[9][19]  ( .D(n9252), .CK(clk), .Q(\registers[9][19] ), 
        .QN(n14347) );
  DFF_X1 \registers_reg[10][19]  ( .D(n9251), .CK(clk), .Q(\registers[10][19] ), .QN(n14749) );
  DFF_X1 \registers_reg[11][19]  ( .D(n9250), .CK(clk), .Q(\registers[11][19] ), .QN(n14461) );
  DFF_X1 \registers_reg[12][19]  ( .D(n9249), .CK(clk), .Q(\registers[12][19] ), .QN(n15687) );
  DFF_X1 \registers_reg[13][19]  ( .D(n9248), .CK(clk), .Q(net227252), .QN(
        n15107) );
  DFF_X1 \registers_reg[14][19]  ( .D(n9247), .CK(clk), .QN(n11899) );
  DFF_X1 \registers_reg[15][19]  ( .D(n9246), .CK(clk), .Q(\registers[15][19] ), .QN(n15310) );
  DFF_X1 \registers_reg[16][19]  ( .D(n9245), .CK(clk), .Q(\registers[16][19] ), .QN(n15717) );
  DFF_X1 \registers_reg[17][19]  ( .D(n9244), .CK(clk), .Q(\registers[17][19] ), .QN(n14623) );
  DFF_X1 \registers_reg[18][19]  ( .D(n9243), .CK(clk), .Q(\registers[18][19] ), .QN(n14409) );
  DFF_X1 \registers_reg[19][19]  ( .D(n9242), .CK(clk), .Q(\registers[19][19] ), .QN(n15837) );
  DFF_X1 \registers_reg[20][19]  ( .D(n9241), .CK(clk), .QN(n14849) );
  DFF_X1 \registers_reg[21][19]  ( .D(n9240), .CK(clk), .QN(n12303) );
  DFF_X1 \registers_reg[22][19]  ( .D(n9239), .CK(clk), .Q(\registers[22][19] ), .QN(n15391) );
  DFF_X1 \registers_reg[23][19]  ( .D(n9238), .CK(clk), .Q(\registers[23][19] ), .QN(n15900) );
  DFF_X1 \registers_reg[24][19]  ( .D(n9237), .CK(clk), .Q(net227251), .QN(
        n15198) );
  DFF_X1 \registers_reg[25][19]  ( .D(n9236), .CK(clk), .Q(\registers[25][19] ), .QN(n14317) );
  DFF_X1 \registers_reg[26][19]  ( .D(n9235), .CK(clk), .QN(n14041) );
  DFF_X1 \registers_reg[27][19]  ( .D(n9234), .CK(clk), .QN(n12036) );
  DFF_X1 \registers_reg[28][19]  ( .D(n9233), .CK(clk), .Q(net227250), .QN(
        n15021) );
  DFF_X1 \registers_reg[29][19]  ( .D(n9232), .CK(clk), .Q(\registers[29][19] ), .QN(n15836) );
  DFF_X1 \registers_reg[30][19]  ( .D(n9231), .CK(clk), .Q(\registers[30][19] ), .QN(n14695) );
  DFF_X1 \registers_reg[31][19]  ( .D(n9230), .CK(clk), .Q(net227249), .QN(
        n15753) );
  DFF_X1 \registers_reg[32][19]  ( .D(n9229), .CK(clk), .QN(n12328) );
  DFF_X1 \registers_reg[33][19]  ( .D(n9228), .CK(clk), .QN(n11863) );
  DFF_X1 \registers_reg[34][19]  ( .D(n9227), .CK(clk), .Q(\registers[34][19] ), .QN(n15513) );
  DFF_X1 \registers_reg[35][19]  ( .D(n9226), .CK(clk), .Q(net227248), .QN(
        n15616) );
  DFF_X1 \registers_reg[36][19]  ( .D(n9225), .CK(clk), .Q(\registers[36][19] ), .QN(n15171) );
  DFF_X1 \registers_reg[37][19]  ( .D(n9224), .CK(clk), .Q(\registers[37][19] ), .QN(n14398) );
  DFF_X1 \registers_reg[38][19]  ( .D(n9223), .CK(clk), .Q(\registers[38][19] ), .QN(n15055) );
  DFF_X1 \registers_reg[39][19]  ( .D(n9222), .CK(clk), .QN(n12190) );
  DFF_X1 \registers_reg[40][19]  ( .D(n9221), .CK(clk), .Q(\registers[40][19] ), .QN(n15108) );
  DFF_X1 \registers_reg[41][19]  ( .D(n9220), .CK(clk), .Q(\registers[41][19] ), .QN(n14462) );
  DFF_X1 \registers_reg[42][19]  ( .D(n9219), .CK(clk), .Q(\registers[42][19] ), .QN(n15938) );
  DFF_X1 \registers_reg[43][19]  ( .D(n9218), .CK(clk), .Q(\registers[43][19] ), .QN(n14905) );
  DFF_X1 \registers_reg[44][19]  ( .D(n9217), .CK(clk), .Q(\registers[44][19] ), .QN(n15483) );
  DFF_X1 \registers_reg[45][19]  ( .D(n9216), .CK(clk), .Q(\registers[45][19] ), .QN(n14808) );
  DFF_X1 \registers_reg[46][19]  ( .D(n9215), .CK(clk), .QN(n12011) );
  DFF_X1 \registers_reg[47][19]  ( .D(n9214), .CK(clk), .Q(\registers[47][19] ), .QN(n14564) );
  DFF_X1 \registers_reg[48][19]  ( .D(n9213), .CK(clk), .Q(\registers[48][19] ), .QN(n15569) );
  DFF_X1 \registers_reg[49][19]  ( .D(n9212), .CK(clk), .Q(\registers[49][19] ), .QN(n14501) );
  DFF_X1 \registers_reg[50][19]  ( .D(n9211), .CK(clk), .Q(\registers[50][19] ), .QN(n15987) );
  DFF_X1 \registers_reg[51][19]  ( .D(n9210), .CK(clk), .Q(\registers[51][19] ), .QN(n15416) );
  DFF_X1 \registers_reg[52][19]  ( .D(n9209), .CK(clk), .Q(net227246), .QN(
        n14955) );
  DFF_X1 \registers_reg[53][19]  ( .D(n9208), .CK(clk), .Q(net227245), .QN(
        n15965) );
  DFF_X1 \registers_reg[54][19]  ( .D(n9207), .CK(clk), .Q(\registers[54][19] ), .QN(n14587) );
  DFF_X1 \registers_reg[55][19]  ( .D(n9206), .CK(clk), .Q(\registers[55][19] ), .QN(n12148) );
  DFF_X1 \registers_reg[56][19]  ( .D(n9205), .CK(clk), .Q(\registers[56][19] ), .QN(n16023) );
  DFF_X1 \registers_reg[57][19]  ( .D(n9204), .CK(clk), .Q(net227244), .QN(
        n15259) );
  DFF_X1 \registers_reg[58][19]  ( .D(n9203), .CK(clk), .Q(net227243), .QN(
        n14926) );
  DFF_X1 \registers_reg[59][19]  ( .D(n9202), .CK(clk), .Q(\registers[59][19] ), .QN(n15448) );
  DFF_X1 \registers_reg[60][19]  ( .D(n9201), .CK(clk), .Q(\registers[60][19] ), .QN(n14659) );
  DFF_X1 \registers_reg[61][19]  ( .D(n9200), .CK(clk), .Q(net227242), .QN(
        n15650) );
  DFF_X1 \registers_reg[62][19]  ( .D(n9199), .CK(clk), .Q(\registers[62][19] ), .QN(n15139) );
  DFF_X1 \registers_reg[63][19]  ( .D(n9198), .CK(clk), .Q(\registers[63][19] ), .QN(n14522) );
  DFF_X1 \to_mem_reg[19]  ( .D(n9197), .CK(clk), .QN(n7706) );
  DFF_X1 \registers_reg[64][19]  ( .D(n9196), .CK(clk), .Q(net227241), .QN(
        n16139) );
  DFF_X1 \registers_reg[65][19]  ( .D(n9195), .CK(clk), .Q(net227240), .QN(
        n16088) );
  DFF_X1 \registers_reg[66][19]  ( .D(n9194), .CK(clk), .Q(net227239), .QN(
        n16050) );
  DFF_X1 \registers_reg[67][19]  ( .D(n9193), .CK(clk), .QN(n14269) );
  DFF_X1 \registers_reg[68][19]  ( .D(n9192), .CK(clk), .Q(\registers[68][19] ), .QN(n16176) );
  DFF_X1 \registers_reg[69][19]  ( .D(n9191), .CK(clk), .Q(net227238), .QN(
        n16172) );
  DFF_X1 \registers_reg[70][19]  ( .D(n9190), .CK(clk), .Q(net227237), .QN(
        n16085) );
  DFF_X1 \registers_reg[0][18]  ( .D(n9189), .CK(clk), .Q(\registers[0][18] ), 
        .QN(n15869) );
  DFF_X1 \registers_reg[1][18]  ( .D(n9188), .CK(clk), .Q(\registers[1][18] ), 
        .QN(n15626) );
  DFF_X1 \registers_reg[2][18]  ( .D(n9187), .CK(clk), .Q(\registers[2][18] ), 
        .QN(n14805) );
  DFF_X1 \registers_reg[3][18]  ( .D(n9186), .CK(clk), .Q(net227236), .QN(
        n15776) );
  DFF_X1 \registers_reg[4][18]  ( .D(n9185), .CK(clk), .Q(\registers[4][18] ), 
        .QN(n15539) );
  DFF_X1 \registers_reg[5][18]  ( .D(n9184), .CK(clk), .Q(\registers[5][18] ), 
        .QN(n14746) );
  DFF_X1 \registers_reg[6][18]  ( .D(n9183), .CK(clk), .QN(n14040) );
  DFF_X1 \registers_reg[7][18]  ( .D(n9182), .CK(clk), .Q(\registers[7][18] ), 
        .QN(n15344) );
  DFF_X1 \registers_reg[8][18]  ( .D(n9181), .CK(clk), .Q(net227235), .QN(
        n15227) );
  DFF_X1 \registers_reg[9][18]  ( .D(n9180), .CK(clk), .Q(\registers[9][18] ), 
        .QN(n14346) );
  DFF_X1 \registers_reg[10][18]  ( .D(n9179), .CK(clk), .Q(\registers[10][18] ), .QN(n14747) );
  DFF_X1 \registers_reg[11][18]  ( .D(n9178), .CK(clk), .Q(\registers[11][18] ), .QN(n14459) );
  DFF_X1 \registers_reg[12][18]  ( .D(n9177), .CK(clk), .Q(\registers[12][18] ), .QN(n15686) );
  DFF_X1 \registers_reg[13][18]  ( .D(n9176), .CK(clk), .Q(net227234), .QN(
        n15105) );
  DFF_X1 \registers_reg[14][18]  ( .D(n9175), .CK(clk), .QN(n11898) );
  DFF_X1 \registers_reg[15][18]  ( .D(n9174), .CK(clk), .Q(\registers[15][18] ), .QN(n15309) );
  DFF_X1 \registers_reg[16][18]  ( .D(n9173), .CK(clk), .Q(\registers[16][18] ), .QN(n15716) );
  DFF_X1 \registers_reg[17][18]  ( .D(n9172), .CK(clk), .Q(\registers[17][18] ), .QN(n14622) );
  DFF_X1 \registers_reg[18][18]  ( .D(n9171), .CK(clk), .Q(\registers[18][18] ), .QN(n14408) );
  DFF_X1 \registers_reg[19][18]  ( .D(n9170), .CK(clk), .Q(\registers[19][18] ), .QN(n15835) );
  DFF_X1 \registers_reg[20][18]  ( .D(n9169), .CK(clk), .QN(n14848) );
  DFF_X1 \registers_reg[21][18]  ( .D(n9168), .CK(clk), .QN(n12301) );
  DFF_X1 \registers_reg[22][18]  ( .D(n9167), .CK(clk), .Q(\registers[22][18] ), .QN(n15389) );
  DFF_X1 \registers_reg[23][18]  ( .D(n9166), .CK(clk), .Q(\registers[23][18] ), .QN(n15899) );
  DFF_X1 \registers_reg[24][18]  ( .D(n9165), .CK(clk), .Q(net227233), .QN(
        n15197) );
  DFF_X1 \registers_reg[25][18]  ( .D(n9164), .CK(clk), .Q(\registers[25][18] ), .QN(n14316) );
  DFF_X1 \registers_reg[26][18]  ( .D(n9163), .CK(clk), .QN(n14039) );
  DFF_X1 \registers_reg[27][18]  ( .D(n9162), .CK(clk), .QN(n12035) );
  DFF_X1 \registers_reg[28][18]  ( .D(n9161), .CK(clk), .Q(net227232), .QN(
        n15020) );
  DFF_X1 \registers_reg[29][18]  ( .D(n9160), .CK(clk), .Q(\registers[29][18] ), .QN(n15834) );
  DFF_X1 \registers_reg[30][18]  ( .D(n9159), .CK(clk), .Q(\registers[30][18] ), .QN(n14694) );
  DFF_X1 \registers_reg[31][18]  ( .D(n9158), .CK(clk), .Q(net227231), .QN(
        n15752) );
  DFF_X1 \registers_reg[32][18]  ( .D(n9157), .CK(clk), .QN(n12327) );
  DFF_X1 \registers_reg[33][18]  ( .D(n9156), .CK(clk), .QN(n11862) );
  DFF_X1 \registers_reg[34][18]  ( .D(n9155), .CK(clk), .Q(\registers[34][18] ), .QN(n15512) );
  DFF_X1 \registers_reg[35][18]  ( .D(n9154), .CK(clk), .Q(net227230), .QN(
        n15613) );
  DFF_X1 \registers_reg[36][18]  ( .D(n9153), .CK(clk), .Q(\registers[36][18] ), .QN(n15170) );
  DFF_X1 \registers_reg[37][18]  ( .D(n9152), .CK(clk), .Q(\registers[37][18] ), .QN(n14395) );
  DFF_X1 \registers_reg[38][18]  ( .D(n9151), .CK(clk), .Q(\registers[38][18] ), .QN(n15053) );
  DFF_X1 \registers_reg[39][18]  ( .D(n9150), .CK(clk), .QN(n12189) );
  DFF_X1 \registers_reg[40][18]  ( .D(n9149), .CK(clk), .Q(\registers[40][18] ), .QN(n15106) );
  DFF_X1 \registers_reg[41][18]  ( .D(n9148), .CK(clk), .Q(\registers[41][18] ), .QN(n14460) );
  DFF_X1 \registers_reg[42][18]  ( .D(n9147), .CK(clk), .Q(\registers[42][18] ), .QN(n15937) );
  DFF_X1 \registers_reg[43][18]  ( .D(n9146), .CK(clk), .Q(\registers[43][18] ), .QN(n14904) );
  DFF_X1 \registers_reg[44][18]  ( .D(n9145), .CK(clk), .Q(\registers[44][18] ), .QN(n15482) );
  DFF_X1 \registers_reg[45][18]  ( .D(n9144), .CK(clk), .Q(\registers[45][18] ), .QN(n14806) );
  DFF_X1 \registers_reg[46][18]  ( .D(n9143), .CK(clk), .QN(n12010) );
  DFF_X1 \registers_reg[47][18]  ( .D(n9142), .CK(clk), .Q(\registers[47][18] ), .QN(n14563) );
  DFF_X1 \registers_reg[48][18]  ( .D(n9141), .CK(clk), .Q(\registers[48][18] ), .QN(n15568) );
  DFF_X1 \registers_reg[49][18]  ( .D(n9140), .CK(clk), .Q(\registers[49][18] ), .QN(n14500) );
  DFF_X1 \registers_reg[50][18]  ( .D(n9139), .CK(clk), .Q(\registers[50][18] ), .QN(n15986) );
  DFF_X1 \registers_reg[51][18]  ( .D(n9138), .CK(clk), .Q(\registers[51][18] ), .QN(n15415) );
  DFF_X1 \registers_reg[52][18]  ( .D(n9137), .CK(clk), .Q(net227228), .QN(
        n14954) );
  DFF_X1 \registers_reg[53][18]  ( .D(n9136), .CK(clk), .Q(net227227), .QN(
        n15964) );
  DFF_X1 \registers_reg[54][18]  ( .D(n9135), .CK(clk), .Q(\registers[54][18] ), .QN(n14586) );
  DFF_X1 \registers_reg[55][18]  ( .D(n9134), .CK(clk), .Q(\registers[55][18] ), .QN(n12105) );
  DFF_X1 \registers_reg[56][18]  ( .D(n9133), .CK(clk), .Q(\registers[56][18] ), .QN(n16022) );
  DFF_X1 \registers_reg[57][18]  ( .D(n9132), .CK(clk), .Q(net227226), .QN(
        n15258) );
  DFF_X1 \registers_reg[58][18]  ( .D(n9131), .CK(clk), .Q(net227225), .QN(
        n14925) );
  DFF_X1 \registers_reg[59][18]  ( .D(n9130), .CK(clk), .Q(\registers[59][18] ), .QN(n15447) );
  DFF_X1 \registers_reg[60][18]  ( .D(n9129), .CK(clk), .Q(\registers[60][18] ), .QN(n14658) );
  DFF_X1 \registers_reg[61][18]  ( .D(n9128), .CK(clk), .Q(net227224), .QN(
        n15649) );
  DFF_X1 \registers_reg[62][18]  ( .D(n9127), .CK(clk), .Q(\registers[62][18] ), .QN(n15138) );
  DFF_X1 \registers_reg[63][18]  ( .D(n9126), .CK(clk), .Q(\registers[63][18] ), .QN(n14521) );
  DFF_X1 \to_mem_reg[18]  ( .D(n9125), .CK(clk), .QN(n7707) );
  DFF_X1 \registers_reg[64][18]  ( .D(n9124), .CK(clk), .Q(net227223), .QN(
        n16138) );
  DFF_X1 \registers_reg[65][18]  ( .D(n9123), .CK(clk), .Q(net227222), .QN(
        n16109) );
  DFF_X1 \registers_reg[66][18]  ( .D(n9122), .CK(clk), .Q(net227221), .QN(
        n16081) );
  DFF_X1 \registers_reg[67][18]  ( .D(n9121), .CK(clk), .QN(n14264) );
  DFF_X1 \registers_reg[68][18]  ( .D(n9120), .CK(clk), .Q(\registers[68][18] ), .QN(n16197) );
  DFF_X1 \registers_reg[69][18]  ( .D(n9119), .CK(clk), .Q(net227220), .QN(
        n16171) );
  DFF_X1 \registers_reg[70][18]  ( .D(n9118), .CK(clk), .Q(net227219), .QN(
        n16080) );
  DFF_X1 \registers_reg[0][17]  ( .D(n9117), .CK(clk), .Q(\registers[0][17] ), 
        .QN(n15868) );
  DFF_X1 \registers_reg[1][17]  ( .D(n9116), .CK(clk), .Q(\registers[1][17] ), 
        .QN(n15612) );
  DFF_X1 \registers_reg[2][17]  ( .D(n9115), .CK(clk), .Q(\registers[2][17] ), 
        .QN(n14803) );
  DFF_X1 \registers_reg[3][17]  ( .D(n9114), .CK(clk), .Q(net227218), .QN(
        n15775) );
  DFF_X1 \registers_reg[4][17]  ( .D(n9113), .CK(clk), .Q(\registers[4][17] ), 
        .QN(n15538) );
  DFF_X1 \registers_reg[5][17]  ( .D(n9112), .CK(clk), .Q(\registers[5][17] ), 
        .QN(n14744) );
  DFF_X1 \registers_reg[6][17]  ( .D(n9111), .CK(clk), .QN(n14038) );
  DFF_X1 \registers_reg[7][17]  ( .D(n9110), .CK(clk), .Q(\registers[7][17] ), 
        .QN(n15343) );
  DFF_X1 \registers_reg[8][17]  ( .D(n9109), .CK(clk), .Q(net227217), .QN(
        n15226) );
  DFF_X1 \registers_reg[9][17]  ( .D(n9108), .CK(clk), .Q(\registers[9][17] ), 
        .QN(n14345) );
  DFF_X1 \registers_reg[10][17]  ( .D(n9107), .CK(clk), .Q(\registers[10][17] ), .QN(n14745) );
  DFF_X1 \registers_reg[11][17]  ( .D(n9106), .CK(clk), .Q(\registers[11][17] ), .QN(n14457) );
  DFF_X1 \registers_reg[12][17]  ( .D(n9105), .CK(clk), .Q(\registers[12][17] ), .QN(n15685) );
  DFF_X1 \registers_reg[13][17]  ( .D(n9104), .CK(clk), .Q(net227216), .QN(
        n15103) );
  DFF_X1 \registers_reg[14][17]  ( .D(n9103), .CK(clk), .QN(n11897) );
  DFF_X1 \registers_reg[15][17]  ( .D(n9102), .CK(clk), .Q(\registers[15][17] ), .QN(n15308) );
  DFF_X1 \registers_reg[16][17]  ( .D(n9101), .CK(clk), .Q(\registers[16][17] ), .QN(n15715) );
  DFF_X1 \registers_reg[17][17]  ( .D(n9100), .CK(clk), .Q(\registers[17][17] ), .QN(n14621) );
  DFF_X1 \registers_reg[18][17]  ( .D(n9099), .CK(clk), .Q(\registers[18][17] ), .QN(n14394) );
  DFF_X1 \registers_reg[19][17]  ( .D(n9098), .CK(clk), .Q(\registers[19][17] ), .QN(n15833) );
  DFF_X1 \registers_reg[20][17]  ( .D(n9097), .CK(clk), .QN(n14847) );
  DFF_X1 \registers_reg[21][17]  ( .D(n9096), .CK(clk), .QN(n12258) );
  DFF_X1 \registers_reg[22][17]  ( .D(n9095), .CK(clk), .Q(\registers[22][17] ), .QN(n15388) );
  DFF_X1 \registers_reg[23][17]  ( .D(n9094), .CK(clk), .Q(\registers[23][17] ), .QN(n15898) );
  DFF_X1 \registers_reg[24][17]  ( .D(n9093), .CK(clk), .Q(net227215), .QN(
        n15196) );
  DFF_X1 \registers_reg[25][17]  ( .D(n9092), .CK(clk), .Q(\registers[25][17] ), .QN(n14315) );
  DFF_X1 \registers_reg[26][17]  ( .D(n9091), .CK(clk), .QN(n14037) );
  DFF_X1 \registers_reg[27][17]  ( .D(n9090), .CK(clk), .QN(n12034) );
  DFF_X1 \registers_reg[28][17]  ( .D(n9089), .CK(clk), .Q(net227214), .QN(
        n15019) );
  DFF_X1 \registers_reg[29][17]  ( .D(n9088), .CK(clk), .Q(\registers[29][17] ), .QN(n15832) );
  DFF_X1 \registers_reg[30][17]  ( .D(n9087), .CK(clk), .Q(\registers[30][17] ), .QN(n14693) );
  DFF_X1 \registers_reg[31][17]  ( .D(n9086), .CK(clk), .Q(net227213), .QN(
        n15751) );
  DFF_X1 \registers_reg[32][17]  ( .D(n9085), .CK(clk), .QN(n12326) );
  DFF_X1 \registers_reg[33][17]  ( .D(n9084), .CK(clk), .QN(n11860) );
  DFF_X1 \registers_reg[34][17]  ( .D(n9083), .CK(clk), .Q(\registers[34][17] ), .QN(n15511) );
  DFF_X1 \registers_reg[35][17]  ( .D(n9082), .CK(clk), .Q(net227212), .QN(
        n15611) );
  DFF_X1 \registers_reg[36][17]  ( .D(n9081), .CK(clk), .Q(\registers[36][17] ), .QN(n15168) );
  DFF_X1 \registers_reg[37][17]  ( .D(n9080), .CK(clk), .Q(\registers[37][17] ), .QN(n14393) );
  DFF_X1 \registers_reg[38][17]  ( .D(n9079), .CK(clk), .Q(\registers[38][17] ), .QN(n15052) );
  DFF_X1 \registers_reg[39][17]  ( .D(n9078), .CK(clk), .QN(n12188) );
  DFF_X1 \registers_reg[40][17]  ( .D(n9077), .CK(clk), .Q(\registers[40][17] ), .QN(n15104) );
  DFF_X1 \registers_reg[41][17]  ( .D(n9076), .CK(clk), .Q(\registers[41][17] ), .QN(n14458) );
  DFF_X1 \registers_reg[42][17]  ( .D(n9075), .CK(clk), .Q(\registers[42][17] ), .QN(n15936) );
  DFF_X1 \registers_reg[43][17]  ( .D(n9074), .CK(clk), .Q(\registers[43][17] ), .QN(n14903) );
  DFF_X1 \registers_reg[44][17]  ( .D(n9073), .CK(clk), .Q(\registers[44][17] ), .QN(n15481) );
  DFF_X1 \registers_reg[45][17]  ( .D(n9072), .CK(clk), .Q(\registers[45][17] ), .QN(n14804) );
  DFF_X1 \registers_reg[46][17]  ( .D(n9071), .CK(clk), .QN(n12009) );
  DFF_X1 \registers_reg[47][17]  ( .D(n9070), .CK(clk), .Q(\registers[47][17] ), .QN(n14562) );
  DFF_X1 \registers_reg[48][17]  ( .D(n9069), .CK(clk), .Q(\registers[48][17] ), .QN(n15567) );
  DFF_X1 \registers_reg[49][17]  ( .D(n9068), .CK(clk), .Q(\registers[49][17] ), .QN(n14499) );
  DFF_X1 \registers_reg[50][17]  ( .D(n9067), .CK(clk), .Q(\registers[50][17] ), .QN(n15985) );
  DFF_X1 \registers_reg[51][17]  ( .D(n9066), .CK(clk), .Q(\registers[51][17] ), .QN(n15414) );
  DFF_X1 \registers_reg[52][17]  ( .D(n9065), .CK(clk), .Q(net227210), .QN(
        n14953) );
  DFF_X1 \registers_reg[53][17]  ( .D(n9064), .CK(clk), .Q(net227209), .QN(
        n15963) );
  DFF_X1 \registers_reg[54][17]  ( .D(n9063), .CK(clk), .Q(\registers[54][17] ), .QN(n14585) );
  DFF_X1 \registers_reg[55][17]  ( .D(n9062), .CK(clk), .Q(\registers[55][17] ), .QN(n12104) );
  DFF_X1 \registers_reg[56][17]  ( .D(n9061), .CK(clk), .Q(\registers[56][17] ), .QN(n16021) );
  DFF_X1 \registers_reg[57][17]  ( .D(n9060), .CK(clk), .Q(net227208), .QN(
        n15257) );
  DFF_X1 \registers_reg[58][17]  ( .D(n9059), .CK(clk), .Q(net227207), .QN(
        n14924) );
  DFF_X1 \registers_reg[59][17]  ( .D(n9058), .CK(clk), .Q(\registers[59][17] ), .QN(n15446) );
  DFF_X1 \registers_reg[60][17]  ( .D(n9057), .CK(clk), .Q(\registers[60][17] ), .QN(n14657) );
  DFF_X1 \registers_reg[61][17]  ( .D(n9056), .CK(clk), .Q(net227206), .QN(
        n15648) );
  DFF_X1 \registers_reg[62][17]  ( .D(n9055), .CK(clk), .Q(\registers[62][17] ), .QN(n15137) );
  DFF_X1 \registers_reg[63][17]  ( .D(n9054), .CK(clk), .Q(\registers[63][17] ), .QN(n14520) );
  DFF_X1 \to_mem_reg[17]  ( .D(n9053), .CK(clk), .QN(n7708) );
  DFF_X1 \registers_reg[64][17]  ( .D(n9052), .CK(clk), .Q(net227205), .QN(
        n16159) );
  DFF_X1 \registers_reg[65][17]  ( .D(n9051), .CK(clk), .Q(net227204), .QN(
        n16108) );
  DFF_X1 \registers_reg[66][17]  ( .D(n9050), .CK(clk), .Q(net227203), .QN(
        n16079) );
  DFF_X1 \registers_reg[67][17]  ( .D(n9049), .CK(clk), .QN(n14261) );
  DFF_X1 \registers_reg[68][17]  ( .D(n9048), .CK(clk), .Q(\registers[68][17] ), .QN(n16196) );
  DFF_X1 \registers_reg[69][17]  ( .D(n9047), .CK(clk), .Q(net227202), .QN(
        n16170) );
  DFF_X1 \registers_reg[70][17]  ( .D(n9046), .CK(clk), .Q(net227201), .QN(
        n16078) );
  DFF_X1 \registers_reg[0][16]  ( .D(n9045), .CK(clk), .Q(\registers[0][16] ), 
        .QN(n15867) );
  DFF_X1 \registers_reg[1][16]  ( .D(n9044), .CK(clk), .Q(\registers[1][16] ), 
        .QN(n15610) );
  DFF_X1 \registers_reg[2][16]  ( .D(n9043), .CK(clk), .Q(\registers[2][16] ), 
        .QN(n14801) );
  DFF_X1 \registers_reg[3][16]  ( .D(n9042), .CK(clk), .Q(net227200), .QN(
        n15774) );
  DFF_X1 \registers_reg[4][16]  ( .D(n9041), .CK(clk), .Q(\registers[4][16] ), 
        .QN(n15537) );
  DFF_X1 \registers_reg[5][16]  ( .D(n9040), .CK(clk), .Q(\registers[5][16] ), 
        .QN(n14742) );
  DFF_X1 \registers_reg[6][16]  ( .D(n9039), .CK(clk), .QN(n14036) );
  DFF_X1 \registers_reg[7][16]  ( .D(n9038), .CK(clk), .Q(\registers[7][16] ), 
        .QN(n15342) );
  DFF_X1 \registers_reg[8][16]  ( .D(n9037), .CK(clk), .Q(net227199), .QN(
        n15225) );
  DFF_X1 \registers_reg[9][16]  ( .D(n9036), .CK(clk), .Q(\registers[9][16] ), 
        .QN(n14344) );
  DFF_X1 \registers_reg[10][16]  ( .D(n9035), .CK(clk), .Q(\registers[10][16] ), .QN(n14743) );
  DFF_X1 \registers_reg[11][16]  ( .D(n9034), .CK(clk), .Q(\registers[11][16] ), .QN(n14455) );
  DFF_X1 \registers_reg[12][16]  ( .D(n9033), .CK(clk), .Q(\registers[12][16] ), .QN(n15684) );
  DFF_X1 \registers_reg[13][16]  ( .D(n9032), .CK(clk), .Q(net227198), .QN(
        n15101) );
  DFF_X1 \registers_reg[14][16]  ( .D(n9031), .CK(clk), .QN(n11896) );
  DFF_X1 \registers_reg[15][16]  ( .D(n9030), .CK(clk), .Q(\registers[15][16] ), .QN(n15307) );
  DFF_X1 \registers_reg[16][16]  ( .D(n9029), .CK(clk), .Q(\registers[16][16] ), .QN(n15714) );
  DFF_X1 \registers_reg[17][16]  ( .D(n9028), .CK(clk), .Q(\registers[17][16] ), .QN(n14620) );
  DFF_X1 \registers_reg[18][16]  ( .D(n9027), .CK(clk), .Q(\registers[18][16] ), .QN(n14392) );
  DFF_X1 \registers_reg[19][16]  ( .D(n9026), .CK(clk), .Q(\registers[19][16] ), .QN(n15831) );
  DFF_X1 \registers_reg[20][16]  ( .D(n9025), .CK(clk), .QN(n14846) );
  DFF_X1 \registers_reg[21][16]  ( .D(n9024), .CK(clk), .QN(n12257) );
  DFF_X1 \registers_reg[22][16]  ( .D(n9023), .CK(clk), .Q(\registers[22][16] ), .QN(n15387) );
  DFF_X1 \registers_reg[23][16]  ( .D(n9022), .CK(clk), .Q(\registers[23][16] ), .QN(n15897) );
  DFF_X1 \registers_reg[24][16]  ( .D(n9021), .CK(clk), .Q(net227197), .QN(
        n15195) );
  DFF_X1 \registers_reg[25][16]  ( .D(n9020), .CK(clk), .Q(\registers[25][16] ), .QN(n14314) );
  DFF_X1 \registers_reg[26][16]  ( .D(n9019), .CK(clk), .QN(n14035) );
  DFF_X1 \registers_reg[27][16]  ( .D(n9018), .CK(clk), .QN(n12033) );
  DFF_X1 \registers_reg[28][16]  ( .D(n9017), .CK(clk), .Q(net227196), .QN(
        n15018) );
  DFF_X1 \registers_reg[29][16]  ( .D(n9016), .CK(clk), .Q(\registers[29][16] ), .QN(n15830) );
  DFF_X1 \registers_reg[30][16]  ( .D(n9015), .CK(clk), .Q(\registers[30][16] ), .QN(n14692) );
  DFF_X1 \registers_reg[31][16]  ( .D(n9014), .CK(clk), .Q(net227195), .QN(
        n15750) );
  DFF_X1 \registers_reg[32][16]  ( .D(n9013), .CK(clk), .QN(n12325) );
  DFF_X1 \registers_reg[33][16]  ( .D(n9012), .CK(clk), .QN(n11858) );
  DFF_X1 \registers_reg[34][16]  ( .D(n9011), .CK(clk), .Q(\registers[34][16] ), .QN(n15510) );
  DFF_X1 \registers_reg[35][16]  ( .D(n9010), .CK(clk), .Q(net227194), .QN(
        n15609) );
  DFF_X1 \registers_reg[36][16]  ( .D(n9009), .CK(clk), .Q(\registers[36][16] ), .QN(n15167) );
  DFF_X1 \registers_reg[37][16]  ( .D(n9008), .CK(clk), .Q(\registers[37][16] ), .QN(n14391) );
  DFF_X1 \registers_reg[38][16]  ( .D(n9007), .CK(clk), .Q(\registers[38][16] ), .QN(n15051) );
  DFF_X1 \registers_reg[39][16]  ( .D(n9006), .CK(clk), .QN(n12187) );
  DFF_X1 \registers_reg[40][16]  ( .D(n9005), .CK(clk), .Q(\registers[40][16] ), .QN(n15102) );
  DFF_X1 \registers_reg[41][16]  ( .D(n9004), .CK(clk), .Q(\registers[41][16] ), .QN(n14456) );
  DFF_X1 \registers_reg[42][16]  ( .D(n9003), .CK(clk), .Q(\registers[42][16] ), .QN(n15935) );
  DFF_X1 \registers_reg[43][16]  ( .D(n9002), .CK(clk), .Q(\registers[43][16] ), .QN(n14902) );
  DFF_X1 \registers_reg[44][16]  ( .D(n9001), .CK(clk), .Q(\registers[44][16] ), .QN(n15480) );
  DFF_X1 \registers_reg[45][16]  ( .D(n9000), .CK(clk), .Q(\registers[45][16] ), .QN(n14802) );
  DFF_X1 \registers_reg[46][16]  ( .D(n8999), .CK(clk), .QN(n12008) );
  DFF_X1 \registers_reg[47][16]  ( .D(n8998), .CK(clk), .Q(\registers[47][16] ), .QN(n14561) );
  DFF_X1 \registers_reg[48][16]  ( .D(n8997), .CK(clk), .Q(\registers[48][16] ), .QN(n15566) );
  DFF_X1 \registers_reg[49][16]  ( .D(n8996), .CK(clk), .Q(\registers[49][16] ), .QN(n14498) );
  DFF_X1 \registers_reg[50][16]  ( .D(n8995), .CK(clk), .Q(\registers[50][16] ), .QN(n15984) );
  DFF_X1 \registers_reg[51][16]  ( .D(n8994), .CK(clk), .Q(\registers[51][16] ), .QN(n15413) );
  DFF_X1 \registers_reg[52][16]  ( .D(n8993), .CK(clk), .Q(net227192), .QN(
        n14952) );
  DFF_X1 \registers_reg[53][16]  ( .D(n8992), .CK(clk), .Q(net227191), .QN(
        n15962) );
  DFF_X1 \registers_reg[54][16]  ( .D(n8991), .CK(clk), .Q(\registers[54][16] ), .QN(n14584) );
  DFF_X1 \registers_reg[55][16]  ( .D(n8990), .CK(clk), .Q(\registers[55][16] ), .QN(n12103) );
  DFF_X1 \registers_reg[56][16]  ( .D(n8989), .CK(clk), .Q(\registers[56][16] ), .QN(n16020) );
  DFF_X1 \registers_reg[57][16]  ( .D(n8988), .CK(clk), .Q(net227190), .QN(
        n15256) );
  DFF_X1 \registers_reg[58][16]  ( .D(n8987), .CK(clk), .Q(net227189), .QN(
        n14923) );
  DFF_X1 \registers_reg[59][16]  ( .D(n8986), .CK(clk), .Q(\registers[59][16] ), .QN(n15445) );
  DFF_X1 \registers_reg[60][16]  ( .D(n8985), .CK(clk), .Q(\registers[60][16] ), .QN(n14656) );
  DFF_X1 \registers_reg[61][16]  ( .D(n8984), .CK(clk), .Q(net227188), .QN(
        n15647) );
  DFF_X1 \registers_reg[62][16]  ( .D(n8983), .CK(clk), .Q(\registers[62][16] ), .QN(n15136) );
  DFF_X1 \registers_reg[63][16]  ( .D(n8982), .CK(clk), .Q(\registers[63][16] ), .QN(n14519) );
  DFF_X1 \to_mem_reg[16]  ( .D(n8981), .CK(clk), .QN(n7709) );
  DFF_X1 \registers_reg[64][16]  ( .D(n8980), .CK(clk), .Q(net227187), .QN(
        n16158) );
  DFF_X1 \registers_reg[65][16]  ( .D(n8979), .CK(clk), .Q(net227186), .QN(
        n16107) );
  DFF_X1 \registers_reg[66][16]  ( .D(n8978), .CK(clk), .Q(net227185), .QN(
        n16077) );
  DFF_X1 \registers_reg[67][16]  ( .D(n8977), .CK(clk), .QN(n14255) );
  DFF_X1 \registers_reg[68][16]  ( .D(n8976), .CK(clk), .Q(\registers[68][16] ), .QN(n16195) );
  DFF_X1 \registers_reg[69][16]  ( .D(n8975), .CK(clk), .Q(net227184), .QN(
        n16169) );
  DFF_X1 \registers_reg[70][16]  ( .D(n8974), .CK(clk), .Q(net227183), .QN(
        n16076) );
  DFF_X1 \registers_reg[0][15]  ( .D(n8973), .CK(clk), .Q(\registers[0][15] ), 
        .QN(n15866) );
  DFF_X1 \registers_reg[1][15]  ( .D(n8972), .CK(clk), .Q(\registers[1][15] ), 
        .QN(n15608) );
  DFF_X1 \registers_reg[2][15]  ( .D(n8971), .CK(clk), .Q(\registers[2][15] ), 
        .QN(n14799) );
  DFF_X1 \registers_reg[3][15]  ( .D(n8970), .CK(clk), .Q(net227182), .QN(
        n15773) );
  DFF_X1 \registers_reg[4][15]  ( .D(n8969), .CK(clk), .Q(\registers[4][15] ), 
        .QN(n15536) );
  DFF_X1 \registers_reg[5][15]  ( .D(n8968), .CK(clk), .Q(\registers[5][15] ), 
        .QN(n14740) );
  DFF_X1 \registers_reg[6][15]  ( .D(n8967), .CK(clk), .QN(n14032) );
  DFF_X1 \registers_reg[7][15]  ( .D(n8966), .CK(clk), .Q(\registers[7][15] ), 
        .QN(n15341) );
  DFF_X1 \registers_reg[8][15]  ( .D(n8965), .CK(clk), .Q(net227181), .QN(
        n15224) );
  DFF_X1 \registers_reg[9][15]  ( .D(n8964), .CK(clk), .Q(\registers[9][15] ), 
        .QN(n14343) );
  DFF_X1 \registers_reg[10][15]  ( .D(n8963), .CK(clk), .Q(\registers[10][15] ), .QN(n14741) );
  DFF_X1 \registers_reg[11][15]  ( .D(n8962), .CK(clk), .Q(\registers[11][15] ), .QN(n14453) );
  DFF_X1 \registers_reg[12][15]  ( .D(n8961), .CK(clk), .Q(\registers[12][15] ), .QN(n15683) );
  DFF_X1 \registers_reg[13][15]  ( .D(n8960), .CK(clk), .Q(net227180), .QN(
        n15099) );
  DFF_X1 \registers_reg[14][15]  ( .D(n8959), .CK(clk), .QN(n11895) );
  DFF_X1 \registers_reg[15][15]  ( .D(n8958), .CK(clk), .Q(\registers[15][15] ), .QN(n15306) );
  DFF_X1 \registers_reg[16][15]  ( .D(n8957), .CK(clk), .Q(\registers[16][15] ), .QN(n15713) );
  DFF_X1 \registers_reg[17][15]  ( .D(n8956), .CK(clk), .Q(\registers[17][15] ), .QN(n14619) );
  DFF_X1 \registers_reg[18][15]  ( .D(n8955), .CK(clk), .Q(\registers[18][15] ), .QN(n14390) );
  DFF_X1 \registers_reg[19][15]  ( .D(n8954), .CK(clk), .Q(\registers[19][15] ), .QN(n15829) );
  DFF_X1 \registers_reg[20][15]  ( .D(n8953), .CK(clk), .QN(n14845) );
  DFF_X1 \registers_reg[21][15]  ( .D(n8952), .CK(clk), .QN(n12256) );
  DFF_X1 \registers_reg[22][15]  ( .D(n8951), .CK(clk), .Q(\registers[22][15] ), .QN(n15386) );
  DFF_X1 \registers_reg[23][15]  ( .D(n8950), .CK(clk), .Q(\registers[23][15] ), .QN(n15896) );
  DFF_X1 \registers_reg[24][15]  ( .D(n8949), .CK(clk), .Q(net227179), .QN(
        n15194) );
  DFF_X1 \registers_reg[25][15]  ( .D(n8948), .CK(clk), .Q(\registers[25][15] ), .QN(n14313) );
  DFF_X1 \registers_reg[26][15]  ( .D(n8947), .CK(clk), .QN(n14015) );
  DFF_X1 \registers_reg[27][15]  ( .D(n8946), .CK(clk), .QN(n12032) );
  DFF_X1 \registers_reg[28][15]  ( .D(n8945), .CK(clk), .Q(net227178), .QN(
        n15017) );
  DFF_X1 \registers_reg[29][15]  ( .D(n8944), .CK(clk), .Q(\registers[29][15] ), .QN(n15828) );
  DFF_X1 \registers_reg[30][15]  ( .D(n8943), .CK(clk), .Q(\registers[30][15] ), .QN(n14691) );
  DFF_X1 \registers_reg[31][15]  ( .D(n8942), .CK(clk), .Q(net227177), .QN(
        n15749) );
  DFF_X1 \registers_reg[32][15]  ( .D(n8941), .CK(clk), .QN(n12324) );
  DFF_X1 \registers_reg[33][15]  ( .D(n8940), .CK(clk), .QN(n11857) );
  DFF_X1 \registers_reg[34][15]  ( .D(n8939), .CK(clk), .Q(\registers[34][15] ), .QN(n15509) );
  DFF_X1 \registers_reg[35][15]  ( .D(n8938), .CK(clk), .Q(net227176), .QN(
        n15607) );
  DFF_X1 \registers_reg[36][15]  ( .D(n8937), .CK(clk), .Q(\registers[36][15] ), .QN(n15166) );
  DFF_X1 \registers_reg[37][15]  ( .D(n8936), .CK(clk), .Q(\registers[37][15] ), .QN(n14389) );
  DFF_X1 \registers_reg[38][15]  ( .D(n8935), .CK(clk), .Q(\registers[38][15] ), .QN(n15050) );
  DFF_X1 \registers_reg[39][15]  ( .D(n8934), .CK(clk), .QN(n12186) );
  DFF_X1 \registers_reg[40][15]  ( .D(n8933), .CK(clk), .Q(\registers[40][15] ), .QN(n15100) );
  DFF_X1 \registers_reg[41][15]  ( .D(n8932), .CK(clk), .Q(\registers[41][15] ), .QN(n14454) );
  DFF_X1 \registers_reg[42][15]  ( .D(n8931), .CK(clk), .Q(\registers[42][15] ), .QN(n15934) );
  DFF_X1 \registers_reg[43][15]  ( .D(n8930), .CK(clk), .Q(\registers[43][15] ), .QN(n14901) );
  DFF_X1 \registers_reg[44][15]  ( .D(n8929), .CK(clk), .Q(\registers[44][15] ), .QN(n15479) );
  DFF_X1 \registers_reg[45][15]  ( .D(n8928), .CK(clk), .Q(\registers[45][15] ), .QN(n14800) );
  DFF_X1 \registers_reg[46][15]  ( .D(n8927), .CK(clk), .QN(n12007) );
  DFF_X1 \registers_reg[47][15]  ( .D(n8926), .CK(clk), .Q(\registers[47][15] ), .QN(n14560) );
  DFF_X1 \registers_reg[48][15]  ( .D(n8925), .CK(clk), .Q(\registers[48][15] ), .QN(n15565) );
  DFF_X1 \registers_reg[49][15]  ( .D(n8924), .CK(clk), .Q(\registers[49][15] ), .QN(n14497) );
  DFF_X1 \registers_reg[50][15]  ( .D(n8923), .CK(clk), .Q(\registers[50][15] ), .QN(n15983) );
  DFF_X1 \registers_reg[51][15]  ( .D(n8922), .CK(clk), .Q(\registers[51][15] ), .QN(n15412) );
  DFF_X1 \registers_reg[52][15]  ( .D(n8921), .CK(clk), .Q(net227174), .QN(
        n14951) );
  DFF_X1 \registers_reg[53][15]  ( .D(n8920), .CK(clk), .Q(net227173), .QN(
        n15961) );
  DFF_X1 \registers_reg[54][15]  ( .D(n8919), .CK(clk), .Q(\registers[54][15] ), .QN(n14583) );
  DFF_X1 \registers_reg[55][15]  ( .D(n8918), .CK(clk), .Q(\registers[55][15] ), .QN(n12102) );
  DFF_X1 \registers_reg[56][15]  ( .D(n8917), .CK(clk), .Q(\registers[56][15] ), .QN(n16019) );
  DFF_X1 \registers_reg[57][15]  ( .D(n8916), .CK(clk), .Q(net227172), .QN(
        n15255) );
  DFF_X1 \registers_reg[58][15]  ( .D(n8915), .CK(clk), .Q(net227171), .QN(
        n14922) );
  DFF_X1 \registers_reg[59][15]  ( .D(n8914), .CK(clk), .Q(\registers[59][15] ), .QN(n15444) );
  DFF_X1 \registers_reg[60][15]  ( .D(n8913), .CK(clk), .Q(\registers[60][15] ), .QN(n14655) );
  DFF_X1 \registers_reg[61][15]  ( .D(n8912), .CK(clk), .Q(net227170), .QN(
        n15646) );
  DFF_X1 \registers_reg[62][15]  ( .D(n8911), .CK(clk), .Q(\registers[62][15] ), .QN(n15135) );
  DFF_X1 \registers_reg[63][15]  ( .D(n8910), .CK(clk), .Q(\registers[63][15] ), .QN(n14518) );
  DFF_X1 \to_mem_reg[15]  ( .D(n8909), .CK(clk), .QN(n7710) );
  DFF_X1 \registers_reg[64][15]  ( .D(n8908), .CK(clk), .Q(net227169), .QN(
        n16157) );
  DFF_X1 \registers_reg[65][15]  ( .D(n8907), .CK(clk), .Q(net227168), .QN(
        n16106) );
  DFF_X1 \registers_reg[66][15]  ( .D(n8906), .CK(clk), .Q(net227167), .QN(
        n16075) );
  DFF_X1 \registers_reg[67][15]  ( .D(n8905), .CK(clk), .QN(n14246) );
  DFF_X1 \registers_reg[68][15]  ( .D(n8904), .CK(clk), .Q(\registers[68][15] ), .QN(n16194) );
  DFF_X1 \registers_reg[69][15]  ( .D(n8903), .CK(clk), .Q(net227166), .QN(
        n16168) );
  DFF_X1 \registers_reg[70][15]  ( .D(n8902), .CK(clk), .Q(net227165), .QN(
        n16074) );
  DFF_X1 \registers_reg[0][14]  ( .D(n8901), .CK(clk), .Q(\registers[0][14] ), 
        .QN(n15865) );
  DFF_X1 \registers_reg[1][14]  ( .D(n8900), .CK(clk), .Q(\registers[1][14] ), 
        .QN(n15606) );
  DFF_X1 \registers_reg[2][14]  ( .D(n8899), .CK(clk), .Q(\registers[2][14] ), 
        .QN(n14797) );
  DFF_X1 \registers_reg[3][14]  ( .D(n8898), .CK(clk), .Q(net227164), .QN(
        n15772) );
  DFF_X1 \registers_reg[4][14]  ( .D(n8897), .CK(clk), .Q(\registers[4][14] ), 
        .QN(n15535) );
  DFF_X1 \registers_reg[5][14]  ( .D(n8896), .CK(clk), .Q(\registers[5][14] ), 
        .QN(n14738) );
  DFF_X1 \registers_reg[6][14]  ( .D(n8895), .CK(clk), .QN(n14014) );
  DFF_X1 \registers_reg[7][14]  ( .D(n8894), .CK(clk), .Q(\registers[7][14] ), 
        .QN(n15340) );
  DFF_X1 \registers_reg[8][14]  ( .D(n8893), .CK(clk), .Q(net227163), .QN(
        n15223) );
  DFF_X1 \registers_reg[9][14]  ( .D(n8892), .CK(clk), .Q(\registers[9][14] ), 
        .QN(n14342) );
  DFF_X1 \registers_reg[10][14]  ( .D(n8891), .CK(clk), .Q(\registers[10][14] ), .QN(n14739) );
  DFF_X1 \registers_reg[11][14]  ( .D(n8890), .CK(clk), .Q(\registers[11][14] ), .QN(n14451) );
  DFF_X1 \registers_reg[12][14]  ( .D(n8889), .CK(clk), .Q(\registers[12][14] ), .QN(n15682) );
  DFF_X1 \registers_reg[13][14]  ( .D(n8888), .CK(clk), .Q(net227162), .QN(
        n15097) );
  DFF_X1 \registers_reg[14][14]  ( .D(n8887), .CK(clk), .QN(n11894) );
  DFF_X1 \registers_reg[15][14]  ( .D(n8886), .CK(clk), .Q(\registers[15][14] ), .QN(n15305) );
  DFF_X1 \registers_reg[16][14]  ( .D(n8885), .CK(clk), .Q(\registers[16][14] ), .QN(n15712) );
  DFF_X1 \registers_reg[17][14]  ( .D(n8884), .CK(clk), .Q(\registers[17][14] ), .QN(n14618) );
  DFF_X1 \registers_reg[18][14]  ( .D(n8883), .CK(clk), .Q(\registers[18][14] ), .QN(n14388) );
  DFF_X1 \registers_reg[19][14]  ( .D(n8882), .CK(clk), .Q(\registers[19][14] ), .QN(n15827) );
  DFF_X1 \registers_reg[20][14]  ( .D(n8881), .CK(clk), .QN(n14844) );
  DFF_X1 \registers_reg[21][14]  ( .D(n8880), .CK(clk), .QN(n12255) );
  DFF_X1 \registers_reg[22][14]  ( .D(n8879), .CK(clk), .Q(\registers[22][14] ), .QN(n15385) );
  DFF_X1 \registers_reg[23][14]  ( .D(n8878), .CK(clk), .Q(\registers[23][14] ), .QN(n15895) );
  DFF_X1 \registers_reg[24][14]  ( .D(n8877), .CK(clk), .Q(net227161), .QN(
        n15193) );
  DFF_X1 \registers_reg[25][14]  ( .D(n8876), .CK(clk), .Q(\registers[25][14] ), .QN(n14312) );
  DFF_X1 \registers_reg[26][14]  ( .D(n8875), .CK(clk), .QN(n14008) );
  DFF_X1 \registers_reg[27][14]  ( .D(n8874), .CK(clk), .QN(n12031) );
  DFF_X1 \registers_reg[28][14]  ( .D(n8873), .CK(clk), .Q(net227160), .QN(
        n15016) );
  DFF_X1 \registers_reg[29][14]  ( .D(n8872), .CK(clk), .Q(\registers[29][14] ), .QN(n15826) );
  DFF_X1 \registers_reg[30][14]  ( .D(n8871), .CK(clk), .Q(\registers[30][14] ), .QN(n14690) );
  DFF_X1 \registers_reg[31][14]  ( .D(n8870), .CK(clk), .Q(net227159), .QN(
        n15748) );
  DFF_X1 \registers_reg[32][14]  ( .D(n8869), .CK(clk), .QN(n12323) );
  DFF_X1 \registers_reg[33][14]  ( .D(n8868), .CK(clk), .QN(n11856) );
  DFF_X1 \registers_reg[34][14]  ( .D(n8867), .CK(clk), .Q(\registers[34][14] ), .QN(n15508) );
  DFF_X1 \registers_reg[35][14]  ( .D(n8866), .CK(clk), .Q(net227158), .QN(
        n15605) );
  DFF_X1 \registers_reg[36][14]  ( .D(n8865), .CK(clk), .Q(\registers[36][14] ), .QN(n15165) );
  DFF_X1 \registers_reg[37][14]  ( .D(n8864), .CK(clk), .Q(\registers[37][14] ), .QN(n14387) );
  DFF_X1 \registers_reg[38][14]  ( .D(n8863), .CK(clk), .Q(\registers[38][14] ), .QN(n15049) );
  DFF_X1 \registers_reg[39][14]  ( .D(n8862), .CK(clk), .QN(n12185) );
  DFF_X1 \registers_reg[40][14]  ( .D(n8861), .CK(clk), .Q(\registers[40][14] ), .QN(n15098) );
  DFF_X1 \registers_reg[41][14]  ( .D(n8860), .CK(clk), .Q(\registers[41][14] ), .QN(n14452) );
  DFF_X1 \registers_reg[42][14]  ( .D(n8859), .CK(clk), .Q(\registers[42][14] ), .QN(n15933) );
  DFF_X1 \registers_reg[43][14]  ( .D(n8858), .CK(clk), .Q(\registers[43][14] ), .QN(n14900) );
  DFF_X1 \registers_reg[44][14]  ( .D(n8857), .CK(clk), .Q(\registers[44][14] ), .QN(n15478) );
  DFF_X1 \registers_reg[45][14]  ( .D(n8856), .CK(clk), .Q(\registers[45][14] ), .QN(n14798) );
  DFF_X1 \registers_reg[46][14]  ( .D(n8855), .CK(clk), .QN(n12006) );
  DFF_X1 \registers_reg[47][14]  ( .D(n8854), .CK(clk), .Q(\registers[47][14] ), .QN(n14559) );
  DFF_X1 \registers_reg[48][14]  ( .D(n8853), .CK(clk), .Q(\registers[48][14] ), .QN(n15564) );
  DFF_X1 \registers_reg[49][14]  ( .D(n8852), .CK(clk), .Q(\registers[49][14] ), .QN(n14496) );
  DFF_X1 \registers_reg[50][14]  ( .D(n8851), .CK(clk), .Q(\registers[50][14] ), .QN(n15982) );
  DFF_X1 \registers_reg[51][14]  ( .D(n8850), .CK(clk), .Q(\registers[51][14] ), .QN(n15411) );
  DFF_X1 \registers_reg[52][14]  ( .D(n8849), .CK(clk), .Q(net227156), .QN(
        n14950) );
  DFF_X1 \registers_reg[53][14]  ( .D(n8848), .CK(clk), .Q(net227155), .QN(
        n15960) );
  DFF_X1 \registers_reg[54][14]  ( .D(n8847), .CK(clk), .Q(\registers[54][14] ), .QN(n14582) );
  DFF_X1 \registers_reg[55][14]  ( .D(n8846), .CK(clk), .Q(\registers[55][14] ), .QN(n12101) );
  DFF_X1 \registers_reg[56][14]  ( .D(n8845), .CK(clk), .Q(\registers[56][14] ), .QN(n16018) );
  DFF_X1 \registers_reg[57][14]  ( .D(n8844), .CK(clk), .Q(net227154), .QN(
        n15254) );
  DFF_X1 \registers_reg[58][14]  ( .D(n8843), .CK(clk), .Q(net227153), .QN(
        n14921) );
  DFF_X1 \registers_reg[59][14]  ( .D(n8842), .CK(clk), .Q(\registers[59][14] ), .QN(n15443) );
  DFF_X1 \registers_reg[60][14]  ( .D(n8841), .CK(clk), .Q(\registers[60][14] ), .QN(n14654) );
  DFF_X1 \registers_reg[61][14]  ( .D(n8840), .CK(clk), .Q(net227152), .QN(
        n15645) );
  DFF_X1 \registers_reg[62][14]  ( .D(n8839), .CK(clk), .Q(\registers[62][14] ), .QN(n15134) );
  DFF_X1 \registers_reg[63][14]  ( .D(n8838), .CK(clk), .Q(\registers[63][14] ), .QN(n14517) );
  DFF_X1 \to_mem_reg[14]  ( .D(n8837), .CK(clk), .QN(n7711) );
  DFF_X1 \registers_reg[64][14]  ( .D(n8836), .CK(clk), .Q(net227151), .QN(
        n16156) );
  DFF_X1 \registers_reg[65][14]  ( .D(n8835), .CK(clk), .Q(net227150), .QN(
        n16105) );
  DFF_X1 \registers_reg[66][14]  ( .D(n8834), .CK(clk), .Q(net227149), .QN(
        n16073) );
  DFF_X1 \registers_reg[67][14]  ( .D(n8833), .CK(clk), .QN(n14243) );
  DFF_X1 \registers_reg[68][14]  ( .D(n8832), .CK(clk), .Q(\registers[68][14] ), .QN(n16193) );
  DFF_X1 \registers_reg[69][14]  ( .D(n8831), .CK(clk), .Q(net227148), .QN(
        n16167) );
  DFF_X1 \registers_reg[70][14]  ( .D(n8830), .CK(clk), .Q(net227147), .QN(
        n16072) );
  DFF_X1 \registers_reg[0][13]  ( .D(n8829), .CK(clk), .Q(\registers[0][13] ), 
        .QN(n15864) );
  DFF_X1 \registers_reg[1][13]  ( .D(n8828), .CK(clk), .Q(\registers[1][13] ), 
        .QN(n15604) );
  DFF_X1 \registers_reg[2][13]  ( .D(n8827), .CK(clk), .Q(\registers[2][13] ), 
        .QN(n14795) );
  DFF_X1 \registers_reg[3][13]  ( .D(n8826), .CK(clk), .Q(net227146), .QN(
        n15771) );
  DFF_X1 \registers_reg[4][13]  ( .D(n8825), .CK(clk), .Q(\registers[4][13] ), 
        .QN(n15534) );
  DFF_X1 \registers_reg[5][13]  ( .D(n8824), .CK(clk), .Q(\registers[5][13] ), 
        .QN(n14736) );
  DFF_X1 \registers_reg[6][13]  ( .D(n8823), .CK(clk), .QN(n13999) );
  DFF_X1 \registers_reg[7][13]  ( .D(n8822), .CK(clk), .Q(\registers[7][13] ), 
        .QN(n15339) );
  DFF_X1 \registers_reg[8][13]  ( .D(n8821), .CK(clk), .Q(net227145), .QN(
        n15222) );
  DFF_X1 \registers_reg[9][13]  ( .D(n8820), .CK(clk), .Q(\registers[9][13] ), 
        .QN(n14341) );
  DFF_X1 \registers_reg[10][13]  ( .D(n8819), .CK(clk), .Q(\registers[10][13] ), .QN(n14737) );
  DFF_X1 \registers_reg[11][13]  ( .D(n8818), .CK(clk), .Q(\registers[11][13] ), .QN(n14449) );
  DFF_X1 \registers_reg[12][13]  ( .D(n8817), .CK(clk), .Q(\registers[12][13] ), .QN(n15681) );
  DFF_X1 \registers_reg[13][13]  ( .D(n8816), .CK(clk), .Q(net227144), .QN(
        n15095) );
  DFF_X1 \registers_reg[14][13]  ( .D(n8815), .CK(clk), .QN(n11893) );
  DFF_X1 \registers_reg[15][13]  ( .D(n8814), .CK(clk), .Q(\registers[15][13] ), .QN(n15304) );
  DFF_X1 \registers_reg[16][13]  ( .D(n8813), .CK(clk), .Q(\registers[16][13] ), .QN(n15711) );
  DFF_X1 \registers_reg[17][13]  ( .D(n8812), .CK(clk), .Q(\registers[17][13] ), .QN(n14617) );
  DFF_X1 \registers_reg[18][13]  ( .D(n8811), .CK(clk), .Q(\registers[18][13] ), .QN(n14386) );
  DFF_X1 \registers_reg[19][13]  ( .D(n8810), .CK(clk), .Q(\registers[19][13] ), .QN(n15825) );
  DFF_X1 \registers_reg[20][13]  ( .D(n8809), .CK(clk), .QN(n14843) );
  DFF_X1 \registers_reg[21][13]  ( .D(n8808), .CK(clk), .QN(n12254) );
  DFF_X1 \registers_reg[22][13]  ( .D(n8807), .CK(clk), .Q(\registers[22][13] ), .QN(n15384) );
  DFF_X1 \registers_reg[23][13]  ( .D(n8806), .CK(clk), .Q(\registers[23][13] ), .QN(n15894) );
  DFF_X1 \registers_reg[24][13]  ( .D(n8805), .CK(clk), .Q(net227143), .QN(
        n15192) );
  DFF_X1 \registers_reg[25][13]  ( .D(n8804), .CK(clk), .Q(\registers[25][13] ), .QN(n14311) );
  DFF_X1 \registers_reg[26][13]  ( .D(n8803), .CK(clk), .QN(n13996) );
  DFF_X1 \registers_reg[27][13]  ( .D(n8802), .CK(clk), .QN(n12030) );
  DFF_X1 \registers_reg[28][13]  ( .D(n8801), .CK(clk), .Q(net227142), .QN(
        n15015) );
  DFF_X1 \registers_reg[29][13]  ( .D(n8800), .CK(clk), .Q(\registers[29][13] ), .QN(n15824) );
  DFF_X1 \registers_reg[30][13]  ( .D(n8799), .CK(clk), .Q(\registers[30][13] ), .QN(n14689) );
  DFF_X1 \registers_reg[31][13]  ( .D(n8798), .CK(clk), .Q(net227141), .QN(
        n15747) );
  DFF_X1 \registers_reg[32][13]  ( .D(n8797), .CK(clk), .QN(n12322) );
  DFF_X1 \registers_reg[33][13]  ( .D(n8796), .CK(clk), .QN(n11855) );
  DFF_X1 \registers_reg[34][13]  ( .D(n8795), .CK(clk), .Q(\registers[34][13] ), .QN(n15507) );
  DFF_X1 \registers_reg[35][13]  ( .D(n8794), .CK(clk), .Q(net227140), .QN(
        n15603) );
  DFF_X1 \registers_reg[36][13]  ( .D(n8793), .CK(clk), .Q(\registers[36][13] ), .QN(n15164) );
  DFF_X1 \registers_reg[37][13]  ( .D(n8792), .CK(clk), .Q(\registers[37][13] ), .QN(n14385) );
  DFF_X1 \registers_reg[38][13]  ( .D(n8791), .CK(clk), .Q(\registers[38][13] ), .QN(n15048) );
  DFF_X1 \registers_reg[39][13]  ( .D(n8790), .CK(clk), .QN(n12183) );
  DFF_X1 \registers_reg[40][13]  ( .D(n8789), .CK(clk), .Q(\registers[40][13] ), .QN(n15096) );
  DFF_X1 \registers_reg[41][13]  ( .D(n8788), .CK(clk), .Q(\registers[41][13] ), .QN(n14450) );
  DFF_X1 \registers_reg[42][13]  ( .D(n8787), .CK(clk), .Q(\registers[42][13] ), .QN(n15932) );
  DFF_X1 \registers_reg[43][13]  ( .D(n8786), .CK(clk), .Q(\registers[43][13] ), .QN(n14899) );
  DFF_X1 \registers_reg[44][13]  ( .D(n8785), .CK(clk), .Q(\registers[44][13] ), .QN(n15477) );
  DFF_X1 \registers_reg[45][13]  ( .D(n8784), .CK(clk), .Q(\registers[45][13] ), .QN(n14796) );
  DFF_X1 \registers_reg[46][13]  ( .D(n8783), .CK(clk), .QN(n12005) );
  DFF_X1 \registers_reg[47][13]  ( .D(n8782), .CK(clk), .Q(\registers[47][13] ), .QN(n14558) );
  DFF_X1 \registers_reg[48][13]  ( .D(n8781), .CK(clk), .Q(\registers[48][13] ), .QN(n15563) );
  DFF_X1 \registers_reg[49][13]  ( .D(n8780), .CK(clk), .Q(\registers[49][13] ), .QN(n14495) );
  DFF_X1 \registers_reg[50][13]  ( .D(n8779), .CK(clk), .Q(\registers[50][13] ), .QN(n15981) );
  DFF_X1 \registers_reg[51][13]  ( .D(n8778), .CK(clk), .Q(\registers[51][13] ), .QN(n15410) );
  DFF_X1 \registers_reg[52][13]  ( .D(n8777), .CK(clk), .Q(net227138), .QN(
        n14949) );
  DFF_X1 \registers_reg[53][13]  ( .D(n8776), .CK(clk), .Q(net227137), .QN(
        n15959) );
  DFF_X1 \registers_reg[54][13]  ( .D(n8775), .CK(clk), .Q(\registers[54][13] ), .QN(n14581) );
  DFF_X1 \registers_reg[55][13]  ( .D(n8774), .CK(clk), .Q(\registers[55][13] ), .QN(n12100) );
  DFF_X1 \registers_reg[56][13]  ( .D(n8773), .CK(clk), .Q(\registers[56][13] ), .QN(n16017) );
  DFF_X1 \registers_reg[57][13]  ( .D(n8772), .CK(clk), .Q(net227136), .QN(
        n15253) );
  DFF_X1 \registers_reg[58][13]  ( .D(n8771), .CK(clk), .Q(net227135), .QN(
        n14920) );
  DFF_X1 \registers_reg[59][13]  ( .D(n8770), .CK(clk), .Q(\registers[59][13] ), .QN(n15442) );
  DFF_X1 \registers_reg[60][13]  ( .D(n8769), .CK(clk), .Q(\registers[60][13] ), .QN(n14653) );
  DFF_X1 \registers_reg[61][13]  ( .D(n8768), .CK(clk), .Q(net227134), .QN(
        n15644) );
  DFF_X1 \registers_reg[62][13]  ( .D(n8767), .CK(clk), .Q(\registers[62][13] ), .QN(n15133) );
  DFF_X1 \registers_reg[63][13]  ( .D(n8766), .CK(clk), .Q(\registers[63][13] ), .QN(n14516) );
  DFF_X1 \to_mem_reg[13]  ( .D(n8765), .CK(clk), .QN(n7712) );
  DFF_X1 \registers_reg[64][13]  ( .D(n8764), .CK(clk), .Q(net227133), .QN(
        n16155) );
  DFF_X1 \registers_reg[65][13]  ( .D(n8763), .CK(clk), .Q(net227132), .QN(
        n16104) );
  DFF_X1 \registers_reg[66][13]  ( .D(n8762), .CK(clk), .Q(net227131), .QN(
        n16071) );
  DFF_X1 \registers_reg[67][13]  ( .D(n8761), .CK(clk), .QN(n14242) );
  DFF_X1 \registers_reg[68][13]  ( .D(n8760), .CK(clk), .Q(\registers[68][13] ), .QN(n16192) );
  DFF_X1 \registers_reg[69][13]  ( .D(n8759), .CK(clk), .Q(net227130), .QN(
        n16166) );
  DFF_X1 \registers_reg[70][13]  ( .D(n8758), .CK(clk), .Q(net227129), .QN(
        n16070) );
  DFF_X1 \registers_reg[0][12]  ( .D(n8757), .CK(clk), .Q(\registers[0][12] ), 
        .QN(n15863) );
  DFF_X1 \registers_reg[1][12]  ( .D(n8756), .CK(clk), .Q(\registers[1][12] ), 
        .QN(n15602) );
  DFF_X1 \registers_reg[2][12]  ( .D(n8755), .CK(clk), .Q(\registers[2][12] ), 
        .QN(n14793) );
  DFF_X1 \registers_reg[3][12]  ( .D(n8754), .CK(clk), .Q(net227128), .QN(
        n15770) );
  DFF_X1 \registers_reg[4][12]  ( .D(n8753), .CK(clk), .Q(\registers[4][12] ), 
        .QN(n15533) );
  DFF_X1 \registers_reg[5][12]  ( .D(n8752), .CK(clk), .Q(\registers[5][12] ), 
        .QN(n14734) );
  DFF_X1 \registers_reg[6][12]  ( .D(n8751), .CK(clk), .QN(n12669) );
  DFF_X1 \registers_reg[7][12]  ( .D(n8750), .CK(clk), .Q(\registers[7][12] ), 
        .QN(n15338) );
  DFF_X1 \registers_reg[8][12]  ( .D(n8749), .CK(clk), .Q(net227127), .QN(
        n15221) );
  DFF_X1 \registers_reg[9][12]  ( .D(n8748), .CK(clk), .Q(\registers[9][12] ), 
        .QN(n14340) );
  DFF_X1 \registers_reg[10][12]  ( .D(n8747), .CK(clk), .Q(\registers[10][12] ), .QN(n14735) );
  DFF_X1 \registers_reg[11][12]  ( .D(n8746), .CK(clk), .Q(\registers[11][12] ), .QN(n14447) );
  DFF_X1 \registers_reg[12][12]  ( .D(n8745), .CK(clk), .Q(\registers[12][12] ), .QN(n15680) );
  DFF_X1 \registers_reg[13][12]  ( .D(n8744), .CK(clk), .Q(net227126), .QN(
        n15093) );
  DFF_X1 \registers_reg[14][12]  ( .D(n8743), .CK(clk), .QN(n11892) );
  DFF_X1 \registers_reg[15][12]  ( .D(n8742), .CK(clk), .Q(\registers[15][12] ), .QN(n15303) );
  DFF_X1 \registers_reg[16][12]  ( .D(n8741), .CK(clk), .Q(\registers[16][12] ), .QN(n15710) );
  DFF_X1 \registers_reg[17][12]  ( .D(n8740), .CK(clk), .Q(\registers[17][12] ), .QN(n14616) );
  DFF_X1 \registers_reg[18][12]  ( .D(n8739), .CK(clk), .Q(\registers[18][12] ), .QN(n14384) );
  DFF_X1 \registers_reg[19][12]  ( .D(n8738), .CK(clk), .Q(\registers[19][12] ), .QN(n15823) );
  DFF_X1 \registers_reg[20][12]  ( .D(n8737), .CK(clk), .QN(n14842) );
  DFF_X1 \registers_reg[21][12]  ( .D(n8736), .CK(clk), .QN(n12253) );
  DFF_X1 \registers_reg[22][12]  ( .D(n8735), .CK(clk), .Q(\registers[22][12] ), .QN(n15383) );
  DFF_X1 \registers_reg[23][12]  ( .D(n8734), .CK(clk), .Q(\registers[23][12] ), .QN(n15893) );
  DFF_X1 \registers_reg[24][12]  ( .D(n8733), .CK(clk), .Q(net227125), .QN(
        n15191) );
  DFF_X1 \registers_reg[25][12]  ( .D(n8732), .CK(clk), .Q(\registers[25][12] ), .QN(n14310) );
  DFF_X1 \registers_reg[26][12]  ( .D(n8731), .CK(clk), .QN(n12652) );
  DFF_X1 \registers_reg[27][12]  ( .D(n8730), .CK(clk), .QN(n12028) );
  DFF_X1 \registers_reg[28][12]  ( .D(n8729), .CK(clk), .Q(net227124), .QN(
        n15014) );
  DFF_X1 \registers_reg[29][12]  ( .D(n8728), .CK(clk), .Q(\registers[29][12] ), .QN(n15822) );
  DFF_X1 \registers_reg[30][12]  ( .D(n8727), .CK(clk), .Q(\registers[30][12] ), .QN(n14688) );
  DFF_X1 \registers_reg[31][12]  ( .D(n8726), .CK(clk), .Q(net227123), .QN(
        n15746) );
  DFF_X1 \registers_reg[32][12]  ( .D(n8725), .CK(clk), .QN(n12321) );
  DFF_X1 \registers_reg[33][12]  ( .D(n8724), .CK(clk), .QN(n11854) );
  DFF_X1 \registers_reg[34][12]  ( .D(n8723), .CK(clk), .Q(\registers[34][12] ), .QN(n15506) );
  DFF_X1 \registers_reg[35][12]  ( .D(n8722), .CK(clk), .Q(net227122), .QN(
        n15601) );
  DFF_X1 \registers_reg[36][12]  ( .D(n8721), .CK(clk), .Q(\registers[36][12] ), .QN(n15163) );
  DFF_X1 \registers_reg[37][12]  ( .D(n8720), .CK(clk), .Q(\registers[37][12] ), .QN(n14383) );
  DFF_X1 \registers_reg[38][12]  ( .D(n8719), .CK(clk), .Q(\registers[38][12] ), .QN(n15047) );
  DFF_X1 \registers_reg[39][12]  ( .D(n8718), .CK(clk), .QN(n12182) );
  DFF_X1 \registers_reg[40][12]  ( .D(n8717), .CK(clk), .Q(\registers[40][12] ), .QN(n15094) );
  DFF_X1 \registers_reg[41][12]  ( .D(n8716), .CK(clk), .Q(\registers[41][12] ), .QN(n14448) );
  DFF_X1 \registers_reg[42][12]  ( .D(n8715), .CK(clk), .Q(\registers[42][12] ), .QN(n15931) );
  DFF_X1 \registers_reg[43][12]  ( .D(n8714), .CK(clk), .Q(\registers[43][12] ), .QN(n14898) );
  DFF_X1 \registers_reg[44][12]  ( .D(n8713), .CK(clk), .Q(\registers[44][12] ), .QN(n15476) );
  DFF_X1 \registers_reg[45][12]  ( .D(n8712), .CK(clk), .Q(\registers[45][12] ), .QN(n14794) );
  DFF_X1 \registers_reg[46][12]  ( .D(n8711), .CK(clk), .QN(n12004) );
  DFF_X1 \registers_reg[47][12]  ( .D(n8710), .CK(clk), .Q(\registers[47][12] ), .QN(n14557) );
  DFF_X1 \registers_reg[48][12]  ( .D(n8709), .CK(clk), .Q(\registers[48][12] ), .QN(n15562) );
  DFF_X1 \registers_reg[49][12]  ( .D(n8708), .CK(clk), .Q(\registers[49][12] ), .QN(n14494) );
  DFF_X1 \registers_reg[50][12]  ( .D(n8707), .CK(clk), .Q(\registers[50][12] ), .QN(n15980) );
  DFF_X1 \registers_reg[51][12]  ( .D(n8706), .CK(clk), .Q(\registers[51][12] ), .QN(n15409) );
  DFF_X1 \registers_reg[52][12]  ( .D(n8705), .CK(clk), .Q(net227120), .QN(
        n14948) );
  DFF_X1 \registers_reg[53][12]  ( .D(n8704), .CK(clk), .Q(net227119), .QN(
        n15958) );
  DFF_X1 \registers_reg[54][12]  ( .D(n8703), .CK(clk), .Q(\registers[54][12] ), .QN(n14580) );
  DFF_X1 \registers_reg[55][12]  ( .D(n8702), .CK(clk), .Q(\registers[55][12] ), .QN(n12099) );
  DFF_X1 \registers_reg[56][12]  ( .D(n8701), .CK(clk), .Q(\registers[56][12] ), .QN(n16016) );
  DFF_X1 \registers_reg[57][12]  ( .D(n8700), .CK(clk), .Q(net227118), .QN(
        n15252) );
  DFF_X1 \registers_reg[58][12]  ( .D(n8699), .CK(clk), .Q(net227117), .QN(
        n14919) );
  DFF_X1 \registers_reg[59][12]  ( .D(n8698), .CK(clk), .Q(\registers[59][12] ), .QN(n15441) );
  DFF_X1 \registers_reg[60][12]  ( .D(n8697), .CK(clk), .Q(\registers[60][12] ), .QN(n14652) );
  DFF_X1 \registers_reg[61][12]  ( .D(n8696), .CK(clk), .Q(net227116), .QN(
        n15643) );
  DFF_X1 \registers_reg[62][12]  ( .D(n8695), .CK(clk), .Q(\registers[62][12] ), .QN(n15132) );
  DFF_X1 \registers_reg[63][12]  ( .D(n8694), .CK(clk), .Q(\registers[63][12] ), .QN(n14515) );
  DFF_X1 \to_mem_reg[12]  ( .D(n8693), .CK(clk), .QN(n7713) );
  DFF_X1 \registers_reg[64][12]  ( .D(n8692), .CK(clk), .Q(net227115), .QN(
        n16154) );
  DFF_X1 \registers_reg[65][12]  ( .D(n8691), .CK(clk), .Q(net227114), .QN(
        n16103) );
  DFF_X1 \registers_reg[66][12]  ( .D(n8690), .CK(clk), .Q(net227113), .QN(
        n16069) );
  DFF_X1 \registers_reg[67][12]  ( .D(n8689), .CK(clk), .QN(n14235) );
  DFF_X1 \registers_reg[68][12]  ( .D(n8688), .CK(clk), .Q(\registers[68][12] ), .QN(n16191) );
  DFF_X1 \registers_reg[69][12]  ( .D(n8687), .CK(clk), .Q(net227112), .QN(
        n16165) );
  DFF_X1 \registers_reg[70][12]  ( .D(n8686), .CK(clk), .Q(net227111), .QN(
        n16068) );
  DFF_X1 \registers_reg[0][11]  ( .D(n8685), .CK(clk), .Q(\registers[0][11] ), 
        .QN(n15862) );
  DFF_X1 \registers_reg[1][11]  ( .D(n8684), .CK(clk), .Q(\registers[1][11] ), 
        .QN(n15600) );
  DFF_X1 \registers_reg[2][11]  ( .D(n8683), .CK(clk), .Q(\registers[2][11] ), 
        .QN(n14791) );
  DFF_X1 \registers_reg[3][11]  ( .D(n8682), .CK(clk), .Q(net227110), .QN(
        n15769) );
  DFF_X1 \registers_reg[4][11]  ( .D(n8681), .CK(clk), .Q(\registers[4][11] ), 
        .QN(n15532) );
  DFF_X1 \registers_reg[5][11]  ( .D(n8680), .CK(clk), .Q(\registers[5][11] ), 
        .QN(n14732) );
  DFF_X1 \registers_reg[6][11]  ( .D(n8679), .CK(clk), .QN(n12602) );
  DFF_X1 \registers_reg[7][11]  ( .D(n8678), .CK(clk), .Q(\registers[7][11] ), 
        .QN(n15337) );
  DFF_X1 \registers_reg[8][11]  ( .D(n8677), .CK(clk), .Q(net227109), .QN(
        n15220) );
  DFF_X1 \registers_reg[9][11]  ( .D(n8676), .CK(clk), .Q(\registers[9][11] ), 
        .QN(n14339) );
  DFF_X1 \registers_reg[10][11]  ( .D(n8675), .CK(clk), .Q(\registers[10][11] ), .QN(n14733) );
  DFF_X1 \registers_reg[11][11]  ( .D(n8674), .CK(clk), .Q(\registers[11][11] ), .QN(n14445) );
  DFF_X1 \registers_reg[12][11]  ( .D(n8673), .CK(clk), .Q(\registers[12][11] ), .QN(n15679) );
  DFF_X1 \registers_reg[13][11]  ( .D(n8672), .CK(clk), .Q(net227108), .QN(
        n15091) );
  DFF_X1 \registers_reg[14][11]  ( .D(n8671), .CK(clk), .QN(n11891) );
  DFF_X1 \registers_reg[15][11]  ( .D(n8670), .CK(clk), .Q(\registers[15][11] ), .QN(n15302) );
  DFF_X1 \registers_reg[16][11]  ( .D(n8669), .CK(clk), .Q(\registers[16][11] ), .QN(n15709) );
  DFF_X1 \registers_reg[17][11]  ( .D(n8668), .CK(clk), .Q(\registers[17][11] ), .QN(n14615) );
  DFF_X1 \registers_reg[18][11]  ( .D(n8667), .CK(clk), .Q(\registers[18][11] ), .QN(n14382) );
  DFF_X1 \registers_reg[19][11]  ( .D(n8666), .CK(clk), .Q(\registers[19][11] ), .QN(n15821) );
  DFF_X1 \registers_reg[20][11]  ( .D(n8665), .CK(clk), .QN(n14841) );
  DFF_X1 \registers_reg[21][11]  ( .D(n8664), .CK(clk), .QN(n12215) );
  DFF_X1 \registers_reg[22][11]  ( .D(n8663), .CK(clk), .Q(\registers[22][11] ), .QN(n15382) );
  DFF_X1 \registers_reg[23][11]  ( .D(n8662), .CK(clk), .Q(\registers[23][11] ), .QN(n15892) );
  DFF_X1 \registers_reg[24][11]  ( .D(n8661), .CK(clk), .Q(net227107), .QN(
        n15190) );
  DFF_X1 \registers_reg[25][11]  ( .D(n8660), .CK(clk), .Q(\registers[25][11] ), .QN(n14309) );
  DFF_X1 \registers_reg[26][11]  ( .D(n8659), .CK(clk), .QN(n12600) );
  DFF_X1 \registers_reg[27][11]  ( .D(n8658), .CK(clk), .QN(n12027) );
  DFF_X1 \registers_reg[28][11]  ( .D(n8657), .CK(clk), .Q(net227106), .QN(
        n15013) );
  DFF_X1 \registers_reg[29][11]  ( .D(n8656), .CK(clk), .Q(\registers[29][11] ), .QN(n15820) );
  DFF_X1 \registers_reg[30][11]  ( .D(n8655), .CK(clk), .Q(\registers[30][11] ), .QN(n14687) );
  DFF_X1 \registers_reg[31][11]  ( .D(n8654), .CK(clk), .Q(net227105), .QN(
        n15745) );
  DFF_X1 \registers_reg[32][11]  ( .D(n8653), .CK(clk), .QN(n12320) );
  DFF_X1 \registers_reg[33][11]  ( .D(n8652), .CK(clk), .QN(n11852) );
  DFF_X1 \registers_reg[34][11]  ( .D(n8651), .CK(clk), .Q(\registers[34][11] ), .QN(n15505) );
  DFF_X1 \registers_reg[35][11]  ( .D(n8650), .CK(clk), .Q(net227104), .QN(
        n15599) );
  DFF_X1 \registers_reg[36][11]  ( .D(n8649), .CK(clk), .Q(\registers[36][11] ), .QN(n15162) );
  DFF_X1 \registers_reg[37][11]  ( .D(n8648), .CK(clk), .Q(\registers[37][11] ), .QN(n14381) );
  DFF_X1 \registers_reg[38][11]  ( .D(n8647), .CK(clk), .Q(\registers[38][11] ), .QN(n15046) );
  DFF_X1 \registers_reg[39][11]  ( .D(n8646), .CK(clk), .QN(n12181) );
  DFF_X1 \registers_reg[40][11]  ( .D(n8645), .CK(clk), .Q(\registers[40][11] ), .QN(n15092) );
  DFF_X1 \registers_reg[41][11]  ( .D(n8644), .CK(clk), .Q(\registers[41][11] ), .QN(n14446) );
  DFF_X1 \registers_reg[42][11]  ( .D(n8643), .CK(clk), .Q(\registers[42][11] ), .QN(n15930) );
  DFF_X1 \registers_reg[43][11]  ( .D(n8642), .CK(clk), .Q(\registers[43][11] ), .QN(n14897) );
  DFF_X1 \registers_reg[44][11]  ( .D(n8641), .CK(clk), .Q(\registers[44][11] ), .QN(n15475) );
  DFF_X1 \registers_reg[45][11]  ( .D(n8640), .CK(clk), .Q(\registers[45][11] ), .QN(n14792) );
  DFF_X1 \registers_reg[46][11]  ( .D(n8639), .CK(clk), .QN(n12003) );
  DFF_X1 \registers_reg[47][11]  ( .D(n8638), .CK(clk), .Q(\registers[47][11] ), .QN(n14556) );
  DFF_X1 \registers_reg[48][11]  ( .D(n8637), .CK(clk), .Q(\registers[48][11] ), .QN(n15561) );
  DFF_X1 \registers_reg[49][11]  ( .D(n8636), .CK(clk), .Q(\registers[49][11] ), .QN(n14493) );
  DFF_X1 \registers_reg[50][11]  ( .D(n8635), .CK(clk), .Q(\registers[50][11] ), .QN(n15979) );
  DFF_X1 \registers_reg[51][11]  ( .D(n8634), .CK(clk), .Q(\registers[51][11] ), .QN(n15408) );
  DFF_X1 \registers_reg[52][11]  ( .D(n8633), .CK(clk), .Q(net227102), .QN(
        n14947) );
  DFF_X1 \registers_reg[53][11]  ( .D(n8632), .CK(clk), .Q(net227101), .QN(
        n15957) );
  DFF_X1 \registers_reg[54][11]  ( .D(n8631), .CK(clk), .Q(\registers[54][11] ), .QN(n14579) );
  DFF_X1 \registers_reg[55][11]  ( .D(n8630), .CK(clk), .Q(\registers[55][11] ), .QN(n12098) );
  DFF_X1 \registers_reg[56][11]  ( .D(n8629), .CK(clk), .Q(\registers[56][11] ), .QN(n16015) );
  DFF_X1 \registers_reg[57][11]  ( .D(n8628), .CK(clk), .Q(net227100), .QN(
        n15251) );
  DFF_X1 \registers_reg[58][11]  ( .D(n8627), .CK(clk), .Q(net227099), .QN(
        n14918) );
  DFF_X1 \registers_reg[59][11]  ( .D(n8626), .CK(clk), .Q(\registers[59][11] ), .QN(n15440) );
  DFF_X1 \registers_reg[60][11]  ( .D(n8625), .CK(clk), .Q(\registers[60][11] ), .QN(n14651) );
  DFF_X1 \registers_reg[61][11]  ( .D(n8624), .CK(clk), .Q(net227098), .QN(
        n15642) );
  DFF_X1 \registers_reg[62][11]  ( .D(n8623), .CK(clk), .Q(\registers[62][11] ), .QN(n15131) );
  DFF_X1 \registers_reg[63][11]  ( .D(n8622), .CK(clk), .Q(\registers[63][11] ), .QN(n14514) );
  DFF_X1 \to_mem_reg[11]  ( .D(n8621), .CK(clk), .QN(n7714) );
  DFF_X1 \registers_reg[64][11]  ( .D(n8620), .CK(clk), .Q(net227097), .QN(
        n16153) );
  DFF_X1 \registers_reg[65][11]  ( .D(n8619), .CK(clk), .Q(net227096), .QN(
        n16102) );
  DFF_X1 \registers_reg[66][11]  ( .D(n8618), .CK(clk), .Q(net227095), .QN(
        n16067) );
  DFF_X1 \registers_reg[67][11]  ( .D(n8617), .CK(clk), .QN(n14230) );
  DFF_X1 \registers_reg[68][11]  ( .D(n8616), .CK(clk), .Q(\registers[68][11] ), .QN(n16190) );
  DFF_X1 \registers_reg[69][11]  ( .D(n8615), .CK(clk), .Q(net227094), .QN(
        n16164) );
  DFF_X1 \registers_reg[70][11]  ( .D(n8614), .CK(clk), .Q(net227093), .QN(
        n16066) );
  DFF_X1 \registers_reg[0][10]  ( .D(n8613), .CK(clk), .Q(\registers[0][10] ), 
        .QN(n15861) );
  DFF_X1 \registers_reg[1][10]  ( .D(n8612), .CK(clk), .Q(\registers[1][10] ), 
        .QN(n15598) );
  DFF_X1 \registers_reg[2][10]  ( .D(n8611), .CK(clk), .Q(\registers[2][10] ), 
        .QN(n14789) );
  DFF_X1 \registers_reg[3][10]  ( .D(n8610), .CK(clk), .Q(net227092), .QN(
        n15768) );
  DFF_X1 \registers_reg[4][10]  ( .D(n8609), .CK(clk), .Q(\registers[4][10] ), 
        .QN(n15531) );
  DFF_X1 \registers_reg[5][10]  ( .D(n8608), .CK(clk), .Q(\registers[5][10] ), 
        .QN(n14730) );
  DFF_X1 \registers_reg[6][10]  ( .D(n8607), .CK(clk), .QN(n12551) );
  DFF_X1 \registers_reg[7][10]  ( .D(n8606), .CK(clk), .Q(\registers[7][10] ), 
        .QN(n15336) );
  DFF_X1 \registers_reg[8][10]  ( .D(n8605), .CK(clk), .Q(net227091), .QN(
        n15219) );
  DFF_X1 \registers_reg[9][10]  ( .D(n8604), .CK(clk), .Q(\registers[9][10] ), 
        .QN(n14338) );
  DFF_X1 \registers_reg[10][10]  ( .D(n8603), .CK(clk), .Q(\registers[10][10] ), .QN(n14731) );
  DFF_X1 \registers_reg[11][10]  ( .D(n8602), .CK(clk), .Q(\registers[11][10] ), .QN(n14443) );
  DFF_X1 \registers_reg[12][10]  ( .D(n8601), .CK(clk), .Q(\registers[12][10] ), .QN(n15678) );
  DFF_X1 \registers_reg[13][10]  ( .D(n8600), .CK(clk), .Q(net227090), .QN(
        n15089) );
  DFF_X1 \registers_reg[14][10]  ( .D(n8599), .CK(clk), .QN(n11890) );
  DFF_X1 \registers_reg[15][10]  ( .D(n8598), .CK(clk), .Q(\registers[15][10] ), .QN(n15301) );
  DFF_X1 \registers_reg[16][10]  ( .D(n8597), .CK(clk), .Q(\registers[16][10] ), .QN(n15708) );
  DFF_X1 \registers_reg[17][10]  ( .D(n8596), .CK(clk), .Q(\registers[17][10] ), .QN(n14614) );
  DFF_X1 \registers_reg[18][10]  ( .D(n8595), .CK(clk), .Q(\registers[18][10] ), .QN(n14380) );
  DFF_X1 \registers_reg[19][10]  ( .D(n8594), .CK(clk), .Q(\registers[19][10] ), .QN(n15819) );
  DFF_X1 \registers_reg[20][10]  ( .D(n8593), .CK(clk), .QN(n14840) );
  DFF_X1 \registers_reg[21][10]  ( .D(n8592), .CK(clk), .QN(n12214) );
  DFF_X1 \registers_reg[22][10]  ( .D(n8591), .CK(clk), .Q(\registers[22][10] ), .QN(n15381) );
  DFF_X1 \registers_reg[23][10]  ( .D(n8590), .CK(clk), .Q(\registers[23][10] ), .QN(n15891) );
  DFF_X1 \registers_reg[24][10]  ( .D(n8589), .CK(clk), .Q(net227089), .QN(
        n15189) );
  DFF_X1 \registers_reg[25][10]  ( .D(n8588), .CK(clk), .Q(\registers[25][10] ), .QN(n14308) );
  DFF_X1 \registers_reg[26][10]  ( .D(n8587), .CK(clk), .QN(n12411) );
  DFF_X1 \registers_reg[27][10]  ( .D(n8586), .CK(clk), .QN(n12026) );
  DFF_X1 \registers_reg[28][10]  ( .D(n8585), .CK(clk), .Q(net227088), .QN(
        n15012) );
  DFF_X1 \registers_reg[29][10]  ( .D(n8584), .CK(clk), .Q(\registers[29][10] ), .QN(n15818) );
  DFF_X1 \registers_reg[30][10]  ( .D(n8583), .CK(clk), .Q(\registers[30][10] ), .QN(n14686) );
  DFF_X1 \registers_reg[31][10]  ( .D(n8582), .CK(clk), .Q(net227087), .QN(
        n15744) );
  DFF_X1 \registers_reg[32][10]  ( .D(n8581), .CK(clk), .QN(n12319) );
  DFF_X1 \registers_reg[33][10]  ( .D(n8580), .CK(clk), .QN(n11851) );
  DFF_X1 \registers_reg[34][10]  ( .D(n8579), .CK(clk), .Q(\registers[34][10] ), .QN(n15504) );
  DFF_X1 \registers_reg[35][10]  ( .D(n8578), .CK(clk), .Q(net227086), .QN(
        n15597) );
  DFF_X1 \registers_reg[36][10]  ( .D(n8577), .CK(clk), .Q(\registers[36][10] ), .QN(n15161) );
  DFF_X1 \registers_reg[37][10]  ( .D(n8576), .CK(clk), .Q(\registers[37][10] ), .QN(n14379) );
  DFF_X1 \registers_reg[38][10]  ( .D(n8575), .CK(clk), .Q(\registers[38][10] ), .QN(n15045) );
  DFF_X1 \registers_reg[39][10]  ( .D(n8574), .CK(clk), .QN(n12180) );
  DFF_X1 \registers_reg[40][10]  ( .D(n8573), .CK(clk), .Q(\registers[40][10] ), .QN(n15090) );
  DFF_X1 \registers_reg[41][10]  ( .D(n8572), .CK(clk), .Q(\registers[41][10] ), .QN(n14444) );
  DFF_X1 \registers_reg[42][10]  ( .D(n8571), .CK(clk), .Q(\registers[42][10] ), .QN(n15929) );
  DFF_X1 \registers_reg[43][10]  ( .D(n8570), .CK(clk), .Q(\registers[43][10] ), .QN(n14896) );
  DFF_X1 \registers_reg[44][10]  ( .D(n8569), .CK(clk), .Q(\registers[44][10] ), .QN(n15474) );
  DFF_X1 \registers_reg[45][10]  ( .D(n8568), .CK(clk), .Q(\registers[45][10] ), .QN(n14790) );
  DFF_X1 \registers_reg[46][10]  ( .D(n8567), .CK(clk), .QN(n12002) );
  DFF_X1 \registers_reg[47][10]  ( .D(n8566), .CK(clk), .Q(\registers[47][10] ), .QN(n14555) );
  DFF_X1 \registers_reg[48][10]  ( .D(n8565), .CK(clk), .Q(\registers[48][10] ), .QN(n15560) );
  DFF_X1 \registers_reg[49][10]  ( .D(n8564), .CK(clk), .Q(\registers[49][10] ), .QN(n14492) );
  DFF_X1 \registers_reg[50][10]  ( .D(n8563), .CK(clk), .Q(\registers[50][10] ), .QN(n15978) );
  DFF_X1 \registers_reg[51][10]  ( .D(n8562), .CK(clk), .Q(\registers[51][10] ), .QN(n15407) );
  DFF_X1 \registers_reg[52][10]  ( .D(n8561), .CK(clk), .Q(net227084), .QN(
        n14946) );
  DFF_X1 \registers_reg[53][10]  ( .D(n8560), .CK(clk), .Q(net227083), .QN(
        n15956) );
  DFF_X1 \registers_reg[54][10]  ( .D(n8559), .CK(clk), .Q(\registers[54][10] ), .QN(n14578) );
  DFF_X1 \registers_reg[55][10]  ( .D(n8558), .CK(clk), .Q(\registers[55][10] ), .QN(n12060) );
  DFF_X1 \registers_reg[56][10]  ( .D(n8557), .CK(clk), .Q(\registers[56][10] ), .QN(n16014) );
  DFF_X1 \registers_reg[57][10]  ( .D(n8556), .CK(clk), .Q(net227082), .QN(
        n15250) );
  DFF_X1 \registers_reg[58][10]  ( .D(n8555), .CK(clk), .Q(net227081), .QN(
        n14917) );
  DFF_X1 \registers_reg[59][10]  ( .D(n8554), .CK(clk), .Q(\registers[59][10] ), .QN(n15439) );
  DFF_X1 \registers_reg[60][10]  ( .D(n8553), .CK(clk), .Q(\registers[60][10] ), .QN(n14650) );
  DFF_X1 \registers_reg[61][10]  ( .D(n8552), .CK(clk), .Q(net227080), .QN(
        n15641) );
  DFF_X1 \registers_reg[62][10]  ( .D(n8551), .CK(clk), .Q(\registers[62][10] ), .QN(n15130) );
  DFF_X1 \registers_reg[63][10]  ( .D(n8550), .CK(clk), .Q(\registers[63][10] ), .QN(n14513) );
  DFF_X1 \to_mem_reg[10]  ( .D(n8549), .CK(clk), .QN(n7715) );
  DFF_X1 \registers_reg[64][10]  ( .D(n8548), .CK(clk), .Q(net227079), .QN(
        n16152) );
  DFF_X1 \registers_reg[65][10]  ( .D(n8547), .CK(clk), .Q(net227078), .QN(
        n16101) );
  DFF_X1 \registers_reg[66][10]  ( .D(n8546), .CK(clk), .Q(net227077), .QN(
        n16065) );
  DFF_X1 \registers_reg[67][10]  ( .D(n8545), .CK(clk), .QN(n14227) );
  DFF_X1 \registers_reg[68][10]  ( .D(n8544), .CK(clk), .Q(\registers[68][10] ), .QN(n16189) );
  DFF_X1 \registers_reg[69][10]  ( .D(n8543), .CK(clk), .Q(net227076), .QN(
        n16163) );
  DFF_X1 \registers_reg[70][10]  ( .D(n8542), .CK(clk), .Q(net227075), .QN(
        n16064) );
  DFF_X1 \registers_reg[0][9]  ( .D(n8541), .CK(clk), .Q(\registers[0][9] ), 
        .QN(n15860) );
  DFF_X1 \registers_reg[1][9]  ( .D(n8540), .CK(clk), .Q(\registers[1][9] ), 
        .QN(n15596) );
  DFF_X1 \registers_reg[2][9]  ( .D(n8539), .CK(clk), .Q(\registers[2][9] ), 
        .QN(n14787) );
  DFF_X1 \registers_reg[3][9]  ( .D(n8538), .CK(clk), .Q(net227074), .QN(
        n15767) );
  DFF_X1 \registers_reg[4][9]  ( .D(n8537), .CK(clk), .Q(\registers[4][9] ), 
        .QN(n15530) );
  DFF_X1 \registers_reg[5][9]  ( .D(n8536), .CK(clk), .Q(\registers[5][9] ), 
        .QN(n14728) );
  DFF_X1 \registers_reg[6][9]  ( .D(n8535), .CK(clk), .QN(n12410) );
  DFF_X1 \registers_reg[7][9]  ( .D(n8534), .CK(clk), .Q(\registers[7][9] ), 
        .QN(n15335) );
  DFF_X1 \registers_reg[8][9]  ( .D(n8533), .CK(clk), .Q(net227073), .QN(
        n15218) );
  DFF_X1 \registers_reg[9][9]  ( .D(n8532), .CK(clk), .Q(\registers[9][9] ), 
        .QN(n14337) );
  DFF_X1 \registers_reg[10][9]  ( .D(n8531), .CK(clk), .Q(\registers[10][9] ), 
        .QN(n14729) );
  DFF_X1 \registers_reg[11][9]  ( .D(n8530), .CK(clk), .Q(\registers[11][9] ), 
        .QN(n14441) );
  DFF_X1 \registers_reg[12][9]  ( .D(n8529), .CK(clk), .Q(\registers[12][9] ), 
        .QN(n15677) );
  DFF_X1 \registers_reg[13][9]  ( .D(n8528), .CK(clk), .Q(net227072), .QN(
        n15087) );
  DFF_X1 \registers_reg[14][9]  ( .D(n8527), .CK(clk), .QN(n11889) );
  DFF_X1 \registers_reg[15][9]  ( .D(n8526), .CK(clk), .Q(\registers[15][9] ), 
        .QN(n15300) );
  DFF_X1 \registers_reg[16][9]  ( .D(n8525), .CK(clk), .Q(\registers[16][9] ), 
        .QN(n15707) );
  DFF_X1 \registers_reg[17][9]  ( .D(n8524), .CK(clk), .Q(\registers[17][9] ), 
        .QN(n14613) );
  DFF_X1 \registers_reg[18][9]  ( .D(n8523), .CK(clk), .Q(\registers[18][9] ), 
        .QN(n14378) );
  DFF_X1 \registers_reg[19][9]  ( .D(n8522), .CK(clk), .Q(\registers[19][9] ), 
        .QN(n15817) );
  DFF_X1 \registers_reg[20][9]  ( .D(n8521), .CK(clk), .QN(n14839) );
  DFF_X1 \registers_reg[21][9]  ( .D(n8520), .CK(clk), .QN(n12213) );
  DFF_X1 \registers_reg[22][9]  ( .D(n8519), .CK(clk), .Q(\registers[22][9] ), 
        .QN(n15380) );
  DFF_X1 \registers_reg[23][9]  ( .D(n8518), .CK(clk), .Q(\registers[23][9] ), 
        .QN(n15890) );
  DFF_X1 \registers_reg[24][9]  ( .D(n8517), .CK(clk), .Q(net227071), .QN(
        n15188) );
  DFF_X1 \registers_reg[25][9]  ( .D(n8516), .CK(clk), .Q(\registers[25][9] ), 
        .QN(n14307) );
  DFF_X1 \registers_reg[26][9]  ( .D(n8515), .CK(clk), .QN(n12409) );
  DFF_X1 \registers_reg[27][9]  ( .D(n8514), .CK(clk), .QN(n12025) );
  DFF_X1 \registers_reg[28][9]  ( .D(n8513), .CK(clk), .Q(net227070), .QN(
        n15011) );
  DFF_X1 \registers_reg[29][9]  ( .D(n8512), .CK(clk), .Q(\registers[29][9] ), 
        .QN(n15816) );
  DFF_X1 \registers_reg[30][9]  ( .D(n8511), .CK(clk), .Q(\registers[30][9] ), 
        .QN(n14685) );
  DFF_X1 \registers_reg[31][9]  ( .D(n8510), .CK(clk), .Q(net227069), .QN(
        n15743) );
  DFF_X1 \registers_reg[32][9]  ( .D(n8509), .CK(clk), .QN(n12318) );
  DFF_X1 \registers_reg[33][9]  ( .D(n8508), .CK(clk), .QN(n11850) );
  DFF_X1 \registers_reg[34][9]  ( .D(n8507), .CK(clk), .Q(\registers[34][9] ), 
        .QN(n15503) );
  DFF_X1 \registers_reg[35][9]  ( .D(n8506), .CK(clk), .Q(net227068), .QN(
        n15595) );
  DFF_X1 \registers_reg[36][9]  ( .D(n8505), .CK(clk), .Q(\registers[36][9] ), 
        .QN(n15160) );
  DFF_X1 \registers_reg[37][9]  ( .D(n8504), .CK(clk), .Q(\registers[37][9] ), 
        .QN(n14377) );
  DFF_X1 \registers_reg[38][9]  ( .D(n8503), .CK(clk), .Q(\registers[38][9] ), 
        .QN(n15044) );
  DFF_X1 \registers_reg[39][9]  ( .D(n8502), .CK(clk), .QN(n12179) );
  DFF_X1 \registers_reg[40][9]  ( .D(n8501), .CK(clk), .Q(\registers[40][9] ), 
        .QN(n15088) );
  DFF_X1 \registers_reg[41][9]  ( .D(n8500), .CK(clk), .Q(\registers[41][9] ), 
        .QN(n14442) );
  DFF_X1 \registers_reg[42][9]  ( .D(n8499), .CK(clk), .Q(\registers[42][9] ), 
        .QN(n15928) );
  DFF_X1 \registers_reg[43][9]  ( .D(n8498), .CK(clk), .Q(\registers[43][9] ), 
        .QN(n14895) );
  DFF_X1 \registers_reg[44][9]  ( .D(n8497), .CK(clk), .Q(\registers[44][9] ), 
        .QN(n15473) );
  DFF_X1 \registers_reg[45][9]  ( .D(n8496), .CK(clk), .Q(\registers[45][9] ), 
        .QN(n14788) );
  DFF_X1 \registers_reg[46][9]  ( .D(n8495), .CK(clk), .QN(n12001) );
  DFF_X1 \registers_reg[47][9]  ( .D(n8494), .CK(clk), .Q(\registers[47][9] ), 
        .QN(n14554) );
  DFF_X1 \registers_reg[48][9]  ( .D(n8493), .CK(clk), .Q(\registers[48][9] ), 
        .QN(n15559) );
  DFF_X1 \registers_reg[49][9]  ( .D(n8492), .CK(clk), .Q(\registers[49][9] ), 
        .QN(n14491) );
  DFF_X1 \registers_reg[50][9]  ( .D(n8491), .CK(clk), .Q(\registers[50][9] ), 
        .QN(n15977) );
  DFF_X1 \registers_reg[51][9]  ( .D(n8490), .CK(clk), .Q(\registers[51][9] ), 
        .QN(n15406) );
  DFF_X1 \registers_reg[52][9]  ( .D(n8489), .CK(clk), .Q(net227066), .QN(
        n14945) );
  DFF_X1 \registers_reg[53][9]  ( .D(n8488), .CK(clk), .Q(net227065), .QN(
        n15919) );
  DFF_X1 \registers_reg[54][9]  ( .D(n8487), .CK(clk), .Q(\registers[54][9] ), 
        .QN(n14577) );
  DFF_X1 \registers_reg[55][9]  ( .D(n8486), .CK(clk), .Q(\registers[55][9] ), 
        .QN(n12059) );
  DFF_X1 \registers_reg[56][9]  ( .D(n8485), .CK(clk), .Q(\registers[56][9] ), 
        .QN(n16003) );
  DFF_X1 \registers_reg[57][9]  ( .D(n8484), .CK(clk), .Q(net227064), .QN(
        n15249) );
  DFF_X1 \registers_reg[58][9]  ( .D(n8483), .CK(clk), .Q(net227063), .QN(
        n14916) );
  DFF_X1 \registers_reg[59][9]  ( .D(n8482), .CK(clk), .Q(\registers[59][9] ), 
        .QN(n15438) );
  DFF_X1 \registers_reg[60][9]  ( .D(n8481), .CK(clk), .Q(\registers[60][9] ), 
        .QN(n14649) );
  DFF_X1 \registers_reg[61][9]  ( .D(n8480), .CK(clk), .Q(net227062), .QN(
        n15640) );
  DFF_X1 \registers_reg[62][9]  ( .D(n8479), .CK(clk), .Q(\registers[62][9] ), 
        .QN(n15129) );
  DFF_X1 \registers_reg[63][9]  ( .D(n8478), .CK(clk), .Q(\registers[63][9] ), 
        .QN(n14512) );
  DFF_X1 \to_mem_reg[9]  ( .D(n8477), .CK(clk), .QN(n7716) );
  DFF_X1 \registers_reg[64][9]  ( .D(n8476), .CK(clk), .Q(net227061), .QN(
        n16151) );
  DFF_X1 \registers_reg[65][9]  ( .D(n8475), .CK(clk), .Q(net227060), .QN(
        n16100) );
  DFF_X1 \registers_reg[66][9]  ( .D(n8474), .CK(clk), .Q(net227059), .QN(
        n16063) );
  DFF_X1 \registers_reg[67][9]  ( .D(n8473), .CK(clk), .QN(n14225) );
  DFF_X1 \registers_reg[68][9]  ( .D(n8472), .CK(clk), .Q(\registers[68][9] ), 
        .QN(n16188) );
  DFF_X1 \registers_reg[69][9]  ( .D(n8471), .CK(clk), .Q(net227058), .QN(
        n16162) );
  DFF_X1 \registers_reg[70][9]  ( .D(n8470), .CK(clk), .Q(net227057), .QN(
        n16062) );
  DFF_X1 \registers_reg[0][8]  ( .D(n8469), .CK(clk), .Q(\registers[0][8] ), 
        .QN(n15859) );
  DFF_X1 \registers_reg[1][8]  ( .D(n8468), .CK(clk), .Q(\registers[1][8] ), 
        .QN(n15594) );
  DFF_X1 \registers_reg[2][8]  ( .D(n8467), .CK(clk), .Q(\registers[2][8] ), 
        .QN(n14785) );
  DFF_X1 \registers_reg[3][8]  ( .D(n8466), .CK(clk), .Q(net227056), .QN(
        n15766) );
  DFF_X1 \registers_reg[4][8]  ( .D(n8465), .CK(clk), .Q(\registers[4][8] ), 
        .QN(n15529) );
  DFF_X1 \registers_reg[5][8]  ( .D(n8464), .CK(clk), .Q(\registers[5][8] ), 
        .QN(n14726) );
  DFF_X1 \registers_reg[6][8]  ( .D(n8463), .CK(clk), .QN(n12408) );
  DFF_X1 \registers_reg[7][8]  ( .D(n8462), .CK(clk), .Q(\registers[7][8] ), 
        .QN(n15334) );
  DFF_X1 \registers_reg[8][8]  ( .D(n8461), .CK(clk), .Q(net227055), .QN(
        n15217) );
  DFF_X1 \registers_reg[9][8]  ( .D(n8460), .CK(clk), .Q(\registers[9][8] ), 
        .QN(n14336) );
  DFF_X1 \registers_reg[10][8]  ( .D(n8459), .CK(clk), .Q(\registers[10][8] ), 
        .QN(n14727) );
  DFF_X1 \registers_reg[11][8]  ( .D(n8458), .CK(clk), .Q(\registers[11][8] ), 
        .QN(n14439) );
  DFF_X1 \registers_reg[12][8]  ( .D(n8457), .CK(clk), .Q(\registers[12][8] ), 
        .QN(n15676) );
  DFF_X1 \registers_reg[13][8]  ( .D(n8456), .CK(clk), .Q(net227054), .QN(
        n15085) );
  DFF_X1 \registers_reg[14][8]  ( .D(n8455), .CK(clk), .QN(n11888) );
  DFF_X1 \registers_reg[15][8]  ( .D(n8454), .CK(clk), .Q(\registers[15][8] ), 
        .QN(n15299) );
  DFF_X1 \registers_reg[16][8]  ( .D(n8453), .CK(clk), .Q(\registers[16][8] ), 
        .QN(n15706) );
  DFF_X1 \registers_reg[17][8]  ( .D(n8452), .CK(clk), .Q(\registers[17][8] ), 
        .QN(n14612) );
  DFF_X1 \registers_reg[18][8]  ( .D(n8451), .CK(clk), .Q(\registers[18][8] ), 
        .QN(n14376) );
  DFF_X1 \registers_reg[19][8]  ( .D(n8450), .CK(clk), .Q(\registers[19][8] ), 
        .QN(n15815) );
  DFF_X1 \registers_reg[20][8]  ( .D(n8449), .CK(clk), .QN(n14838) );
  DFF_X1 \registers_reg[21][8]  ( .D(n8448), .CK(clk), .QN(n12212) );
  DFF_X1 \registers_reg[22][8]  ( .D(n8447), .CK(clk), .Q(\registers[22][8] ), 
        .QN(n15379) );
  DFF_X1 \registers_reg[23][8]  ( .D(n8446), .CK(clk), .Q(\registers[23][8] ), 
        .QN(n15888) );
  DFF_X1 \registers_reg[24][8]  ( .D(n8445), .CK(clk), .Q(net227053), .QN(
        n15187) );
  DFF_X1 \registers_reg[25][8]  ( .D(n8444), .CK(clk), .Q(\registers[25][8] ), 
        .QN(n14306) );
  DFF_X1 \registers_reg[26][8]  ( .D(n8443), .CK(clk), .QN(n12407) );
  DFF_X1 \registers_reg[27][8]  ( .D(n8442), .CK(clk), .QN(n12024) );
  DFF_X1 \registers_reg[28][8]  ( .D(n8441), .CK(clk), .Q(net227052), .QN(
        n15010) );
  DFF_X1 \registers_reg[29][8]  ( .D(n8440), .CK(clk), .Q(\registers[29][8] ), 
        .QN(n15812) );
  DFF_X1 \registers_reg[30][8]  ( .D(n8439), .CK(clk), .Q(\registers[30][8] ), 
        .QN(n14684) );
  DFF_X1 \registers_reg[31][8]  ( .D(n8438), .CK(clk), .Q(net227051), .QN(
        n15742) );
  DFF_X1 \registers_reg[32][8]  ( .D(n8437), .CK(clk), .QN(n12317) );
  DFF_X1 \registers_reg[33][8]  ( .D(n8436), .CK(clk), .QN(n11849) );
  DFF_X1 \registers_reg[34][8]  ( .D(n8435), .CK(clk), .Q(\registers[34][8] ), 
        .QN(n15502) );
  DFF_X1 \registers_reg[35][8]  ( .D(n8434), .CK(clk), .Q(net227050), .QN(
        n15593) );
  DFF_X1 \registers_reg[36][8]  ( .D(n8433), .CK(clk), .Q(\registers[36][8] ), 
        .QN(n15159) );
  DFF_X1 \registers_reg[37][8]  ( .D(n8432), .CK(clk), .Q(\registers[37][8] ), 
        .QN(n14375) );
  DFF_X1 \registers_reg[38][8]  ( .D(n8431), .CK(clk), .Q(\registers[38][8] ), 
        .QN(n15043) );
  DFF_X1 \registers_reg[39][8]  ( .D(n8430), .CK(clk), .QN(n12178) );
  DFF_X1 \registers_reg[40][8]  ( .D(n8429), .CK(clk), .Q(\registers[40][8] ), 
        .QN(n15086) );
  DFF_X1 \registers_reg[41][8]  ( .D(n8428), .CK(clk), .Q(\registers[41][8] ), 
        .QN(n14440) );
  DFF_X1 \registers_reg[42][8]  ( .D(n8427), .CK(clk), .Q(\registers[42][8] ), 
        .QN(n15927) );
  DFF_X1 \registers_reg[43][8]  ( .D(n8426), .CK(clk), .Q(\registers[43][8] ), 
        .QN(n14894) );
  DFF_X1 \registers_reg[44][8]  ( .D(n8425), .CK(clk), .Q(\registers[44][8] ), 
        .QN(n15472) );
  DFF_X1 \registers_reg[45][8]  ( .D(n8424), .CK(clk), .Q(\registers[45][8] ), 
        .QN(n14786) );
  DFF_X1 \registers_reg[46][8]  ( .D(n8423), .CK(clk), .QN(n12000) );
  DFF_X1 \registers_reg[47][8]  ( .D(n8422), .CK(clk), .Q(\registers[47][8] ), 
        .QN(n14553) );
  DFF_X1 \registers_reg[48][8]  ( .D(n8421), .CK(clk), .Q(\registers[48][8] ), 
        .QN(n15558) );
  DFF_X1 \registers_reg[49][8]  ( .D(n8420), .CK(clk), .Q(\registers[49][8] ), 
        .QN(n14490) );
  DFF_X1 \registers_reg[50][8]  ( .D(n8419), .CK(clk), .Q(\registers[50][8] ), 
        .QN(n15976) );
  DFF_X1 \registers_reg[51][8]  ( .D(n8418), .CK(clk), .Q(\registers[51][8] ), 
        .QN(n15405) );
  DFF_X1 \registers_reg[52][8]  ( .D(n8417), .CK(clk), .Q(net227048), .QN(
        n14944) );
  DFF_X1 \registers_reg[53][8]  ( .D(n8416), .CK(clk), .Q(net227047), .QN(
        n15918) );
  DFF_X1 \registers_reg[54][8]  ( .D(n8415), .CK(clk), .Q(\registers[54][8] ), 
        .QN(n14576) );
  DFF_X1 \registers_reg[55][8]  ( .D(n8414), .CK(clk), .Q(\registers[55][8] ), 
        .QN(n12058) );
  DFF_X1 \registers_reg[56][8]  ( .D(n8413), .CK(clk), .Q(\registers[56][8] ), 
        .QN(n16013) );
  DFF_X1 \registers_reg[57][8]  ( .D(n8412), .CK(clk), .Q(net227046), .QN(
        n15248) );
  DFF_X1 \registers_reg[58][8]  ( .D(n8411), .CK(clk), .Q(net227045), .QN(
        n14915) );
  DFF_X1 \registers_reg[59][8]  ( .D(n8410), .CK(clk), .Q(\registers[59][8] ), 
        .QN(n15437) );
  DFF_X1 \registers_reg[60][8]  ( .D(n8409), .CK(clk), .Q(\registers[60][8] ), 
        .QN(n14648) );
  DFF_X1 \registers_reg[61][8]  ( .D(n8408), .CK(clk), .Q(net227044), .QN(
        n15639) );
  DFF_X1 \registers_reg[62][8]  ( .D(n8407), .CK(clk), .Q(\registers[62][8] ), 
        .QN(n15128) );
  DFF_X1 \registers_reg[63][8]  ( .D(n8406), .CK(clk), .Q(\registers[63][8] ), 
        .QN(n14511) );
  DFF_X1 \to_mem_reg[8]  ( .D(n8405), .CK(clk), .QN(n7717) );
  DFF_X1 \registers_reg[64][8]  ( .D(n8404), .CK(clk), .Q(net227043), .QN(
        n16150) );
  DFF_X1 \registers_reg[65][8]  ( .D(n8403), .CK(clk), .Q(net227042), .QN(
        n16099) );
  DFF_X1 \registers_reg[66][8]  ( .D(n8402), .CK(clk), .Q(net227041), .QN(
        n16061) );
  DFF_X1 \registers_reg[67][8]  ( .D(n8401), .CK(clk), .QN(n14219) );
  DFF_X1 \registers_reg[68][8]  ( .D(n8400), .CK(clk), .Q(\registers[68][8] ), 
        .QN(n16187) );
  DFF_X1 \registers_reg[69][8]  ( .D(n8399), .CK(clk), .Q(net227040), .QN(
        n16161) );
  DFF_X1 \registers_reg[70][8]  ( .D(n8398), .CK(clk), .Q(net227039), .QN(
        n16039) );
  DFF_X1 \registers_reg[0][7]  ( .D(n8397), .CK(clk), .Q(\registers[0][7] ), 
        .QN(n15858) );
  DFF_X1 \registers_reg[1][7]  ( .D(n8396), .CK(clk), .Q(\registers[1][7] ), 
        .QN(n15592) );
  DFF_X1 \registers_reg[2][7]  ( .D(n8395), .CK(clk), .Q(\registers[2][7] ), 
        .QN(n14783) );
  DFF_X1 \registers_reg[3][7]  ( .D(n8394), .CK(clk), .Q(net227038), .QN(
        n15765) );
  DFF_X1 \registers_reg[4][7]  ( .D(n8393), .CK(clk), .Q(\registers[4][7] ), 
        .QN(n15528) );
  DFF_X1 \registers_reg[5][7]  ( .D(n8392), .CK(clk), .Q(\registers[5][7] ), 
        .QN(n14724) );
  DFF_X1 \registers_reg[6][7]  ( .D(n8391), .CK(clk), .QN(n12369) );
  DFF_X1 \registers_reg[7][7]  ( .D(n8390), .CK(clk), .Q(\registers[7][7] ), 
        .QN(n15333) );
  DFF_X1 \registers_reg[8][7]  ( .D(n8389), .CK(clk), .Q(net227037), .QN(
        n15216) );
  DFF_X1 \registers_reg[9][7]  ( .D(n8388), .CK(clk), .Q(\registers[9][7] ), 
        .QN(n14335) );
  DFF_X1 \registers_reg[10][7]  ( .D(n8387), .CK(clk), .Q(\registers[10][7] ), 
        .QN(n14725) );
  DFF_X1 \registers_reg[11][7]  ( .D(n8386), .CK(clk), .Q(\registers[11][7] ), 
        .QN(n14437) );
  DFF_X1 \registers_reg[12][7]  ( .D(n8385), .CK(clk), .Q(\registers[12][7] ), 
        .QN(n15675) );
  DFF_X1 \registers_reg[13][7]  ( .D(n8384), .CK(clk), .Q(net227036), .QN(
        n15083) );
  DFF_X1 \registers_reg[14][7]  ( .D(n8383), .CK(clk), .QN(n11887) );
  DFF_X1 \registers_reg[15][7]  ( .D(n8382), .CK(clk), .Q(\registers[15][7] ), 
        .QN(n15298) );
  DFF_X1 \registers_reg[16][7]  ( .D(n8381), .CK(clk), .Q(\registers[16][7] ), 
        .QN(n15705) );
  DFF_X1 \registers_reg[17][7]  ( .D(n8380), .CK(clk), .Q(\registers[17][7] ), 
        .QN(n14611) );
  DFF_X1 \registers_reg[18][7]  ( .D(n8379), .CK(clk), .Q(\registers[18][7] ), 
        .QN(n14374) );
  DFF_X1 \registers_reg[19][7]  ( .D(n8378), .CK(clk), .Q(\registers[19][7] ), 
        .QN(n15811) );
  DFF_X1 \registers_reg[20][7]  ( .D(n8377), .CK(clk), .QN(n14837) );
  DFF_X1 \registers_reg[21][7]  ( .D(n8376), .CK(clk), .QN(n12211) );
  DFF_X1 \registers_reg[22][7]  ( .D(n8375), .CK(clk), .Q(\registers[22][7] ), 
        .QN(n15378) );
  DFF_X1 \registers_reg[23][7]  ( .D(n8374), .CK(clk), .Q(\registers[23][7] ), 
        .QN(n15887) );
  DFF_X1 \registers_reg[24][7]  ( .D(n8373), .CK(clk), .Q(net227035), .QN(
        n15186) );
  DFF_X1 \registers_reg[25][7]  ( .D(n8372), .CK(clk), .Q(\registers[25][7] ), 
        .QN(n14305) );
  DFF_X1 \registers_reg[26][7]  ( .D(n8371), .CK(clk), .QN(n12368) );
  DFF_X1 \registers_reg[27][7]  ( .D(n8370), .CK(clk), .QN(n12023) );
  DFF_X1 \registers_reg[28][7]  ( .D(n8369), .CK(clk), .Q(net227034), .QN(
        n15009) );
  DFF_X1 \registers_reg[29][7]  ( .D(n8368), .CK(clk), .Q(\registers[29][7] ), 
        .QN(n15810) );
  DFF_X1 \registers_reg[30][7]  ( .D(n8367), .CK(clk), .Q(\registers[30][7] ), 
        .QN(n14683) );
  DFF_X1 \registers_reg[31][7]  ( .D(n8366), .CK(clk), .Q(net227033), .QN(
        n15741) );
  DFF_X1 \registers_reg[32][7]  ( .D(n8365), .CK(clk), .QN(n12316) );
  DFF_X1 \registers_reg[33][7]  ( .D(n8364), .CK(clk), .QN(n11847) );
  DFF_X1 \registers_reg[34][7]  ( .D(n8363), .CK(clk), .Q(\registers[34][7] ), 
        .QN(n15501) );
  DFF_X1 \registers_reg[35][7]  ( .D(n8362), .CK(clk), .Q(net227032), .QN(
        n15591) );
  DFF_X1 \registers_reg[36][7]  ( .D(n8361), .CK(clk), .Q(\registers[36][7] ), 
        .QN(n15158) );
  DFF_X1 \registers_reg[37][7]  ( .D(n8360), .CK(clk), .Q(\registers[37][7] ), 
        .QN(n14373) );
  DFF_X1 \registers_reg[38][7]  ( .D(n8359), .CK(clk), .Q(\registers[38][7] ), 
        .QN(n15042) );
  DFF_X1 \registers_reg[39][7]  ( .D(n8358), .CK(clk), .QN(n12177) );
  DFF_X1 \registers_reg[40][7]  ( .D(n8357), .CK(clk), .Q(\registers[40][7] ), 
        .QN(n15084) );
  DFF_X1 \registers_reg[41][7]  ( .D(n8356), .CK(clk), .Q(\registers[41][7] ), 
        .QN(n14438) );
  DFF_X1 \registers_reg[42][7]  ( .D(n8355), .CK(clk), .Q(\registers[42][7] ), 
        .QN(n15925) );
  DFF_X1 \registers_reg[43][7]  ( .D(n8354), .CK(clk), .Q(\registers[43][7] ), 
        .QN(n14893) );
  DFF_X1 \registers_reg[44][7]  ( .D(n8353), .CK(clk), .Q(\registers[44][7] ), 
        .QN(n15471) );
  DFF_X1 \registers_reg[45][7]  ( .D(n8352), .CK(clk), .Q(\registers[45][7] ), 
        .QN(n14784) );
  DFF_X1 \registers_reg[46][7]  ( .D(n8351), .CK(clk), .QN(n11999) );
  DFF_X1 \registers_reg[47][7]  ( .D(n8350), .CK(clk), .Q(\registers[47][7] ), 
        .QN(n14552) );
  DFF_X1 \registers_reg[48][7]  ( .D(n8349), .CK(clk), .Q(\registers[48][7] ), 
        .QN(n15557) );
  DFF_X1 \registers_reg[49][7]  ( .D(n8348), .CK(clk), .Q(\registers[49][7] ), 
        .QN(n14489) );
  DFF_X1 \registers_reg[50][7]  ( .D(n8347), .CK(clk), .Q(\registers[50][7] ), 
        .QN(n15974) );
  DFF_X1 \registers_reg[51][7]  ( .D(n8346), .CK(clk), .Q(\registers[51][7] ), 
        .QN(n15404) );
  DFF_X1 \registers_reg[52][7]  ( .D(n8345), .CK(clk), .Q(net227030), .QN(
        n14943) );
  DFF_X1 \registers_reg[53][7]  ( .D(n8344), .CK(clk), .Q(net227029), .QN(
        n15917) );
  DFF_X1 \registers_reg[54][7]  ( .D(n8343), .CK(clk), .Q(\registers[54][7] ), 
        .QN(n14575) );
  DFF_X1 \registers_reg[55][7]  ( .D(n8342), .CK(clk), .Q(\registers[55][7] ), 
        .QN(n12057) );
  DFF_X1 \registers_reg[56][7]  ( .D(n8341), .CK(clk), .Q(\registers[56][7] ), 
        .QN(n16002) );
  DFF_X1 \registers_reg[57][7]  ( .D(n8340), .CK(clk), .Q(net227028), .QN(
        n15247) );
  DFF_X1 \registers_reg[58][7]  ( .D(n8339), .CK(clk), .Q(net227027), .QN(
        n14914) );
  DFF_X1 \registers_reg[59][7]  ( .D(n8338), .CK(clk), .Q(\registers[59][7] ), 
        .QN(n15436) );
  DFF_X1 \registers_reg[60][7]  ( .D(n8337), .CK(clk), .Q(\registers[60][7] ), 
        .QN(n14647) );
  DFF_X1 \registers_reg[61][7]  ( .D(n8336), .CK(clk), .Q(net227026), .QN(
        n15638) );
  DFF_X1 \registers_reg[62][7]  ( .D(n8335), .CK(clk), .Q(\registers[62][7] ), 
        .QN(n15127) );
  DFF_X1 \registers_reg[63][7]  ( .D(n8334), .CK(clk), .Q(\registers[63][7] ), 
        .QN(n14510) );
  DFF_X1 \to_mem_reg[7]  ( .D(n8333), .CK(clk), .QN(n7718) );
  DFF_X1 \registers_reg[64][7]  ( .D(n8332), .CK(clk), .Q(net227025), .QN(
        n16149) );
  DFF_X1 \registers_reg[65][7]  ( .D(n8331), .CK(clk), .Q(net227024), .QN(
        n16098) );
  DFF_X1 \registers_reg[66][7]  ( .D(n8330), .CK(clk), .Q(net227023), .QN(
        n16060) );
  DFF_X1 \registers_reg[67][7]  ( .D(n8329), .CK(clk), .QN(n14216) );
  DFF_X1 \registers_reg[68][7]  ( .D(n8328), .CK(clk), .Q(\registers[68][7] ), 
        .QN(n16186) );
  DFF_X1 \registers_reg[69][7]  ( .D(n8327), .CK(clk), .Q(net227022), .QN(
        n16128) );
  DFF_X1 \registers_reg[70][7]  ( .D(n8326), .CK(clk), .Q(net227021), .QN(
        n16038) );
  DFF_X1 \registers_reg[0][6]  ( .D(n8325), .CK(clk), .Q(\registers[0][6] ), 
        .QN(n15802) );
  DFF_X1 \registers_reg[1][6]  ( .D(n8324), .CK(clk), .Q(\registers[1][6] ), 
        .QN(n15579) );
  DFF_X1 \registers_reg[2][6]  ( .D(n8323), .CK(clk), .Q(\registers[2][6] ), 
        .QN(n14781) );
  DFF_X1 \registers_reg[3][6]  ( .D(n8322), .CK(clk), .Q(net227020), .QN(
        n15764) );
  DFF_X1 \registers_reg[4][6]  ( .D(n8321), .CK(clk), .Q(\registers[4][6] ), 
        .QN(n15527) );
  DFF_X1 \registers_reg[5][6]  ( .D(n8320), .CK(clk), .Q(\registers[5][6] ), 
        .QN(n14722) );
  DFF_X1 \registers_reg[6][6]  ( .D(n8319), .CK(clk), .QN(n12367) );
  DFF_X1 \registers_reg[7][6]  ( .D(n8318), .CK(clk), .Q(\registers[7][6] ), 
        .QN(n15332) );
  DFF_X1 \registers_reg[8][6]  ( .D(n8317), .CK(clk), .Q(net227019), .QN(
        n15215) );
  DFF_X1 \registers_reg[9][6]  ( .D(n8316), .CK(clk), .Q(\registers[9][6] ), 
        .QN(n14334) );
  DFF_X1 \registers_reg[10][6]  ( .D(n8315), .CK(clk), .Q(\registers[10][6] ), 
        .QN(n14723) );
  DFF_X1 \registers_reg[11][6]  ( .D(n8314), .CK(clk), .Q(\registers[11][6] ), 
        .QN(n14435) );
  DFF_X1 \registers_reg[12][6]  ( .D(n8313), .CK(clk), .Q(\registers[12][6] ), 
        .QN(n15674) );
  DFF_X1 \registers_reg[13][6]  ( .D(n8312), .CK(clk), .Q(net227018), .QN(
        n15081) );
  DFF_X1 \registers_reg[14][6]  ( .D(n8311), .CK(clk), .QN(n11886) );
  DFF_X1 \registers_reg[15][6]  ( .D(n8310), .CK(clk), .Q(\registers[15][6] ), 
        .QN(n15297) );
  DFF_X1 \registers_reg[16][6]  ( .D(n8309), .CK(clk), .Q(\registers[16][6] ), 
        .QN(n15704) );
  DFF_X1 \registers_reg[17][6]  ( .D(n8308), .CK(clk), .Q(\registers[17][6] ), 
        .QN(n14610) );
  DFF_X1 \registers_reg[18][6]  ( .D(n8307), .CK(clk), .Q(\registers[18][6] ), 
        .QN(n14372) );
  DFF_X1 \registers_reg[19][6]  ( .D(n8306), .CK(clk), .Q(\registers[19][6] ), 
        .QN(n15809) );
  DFF_X1 \registers_reg[20][6]  ( .D(n8305), .CK(clk), .QN(n14836) );
  DFF_X1 \registers_reg[21][6]  ( .D(n8304), .CK(clk), .QN(n12210) );
  DFF_X1 \registers_reg[22][6]  ( .D(n8303), .CK(clk), .Q(\registers[22][6] ), 
        .QN(n15376) );
  DFF_X1 \registers_reg[23][6]  ( .D(n8302), .CK(clk), .Q(\registers[23][6] ), 
        .QN(n15886) );
  DFF_X1 \registers_reg[24][6]  ( .D(n8301), .CK(clk), .Q(net227017), .QN(
        n15185) );
  DFF_X1 \registers_reg[25][6]  ( .D(n8300), .CK(clk), .Q(\registers[25][6] ), 
        .QN(n14304) );
  DFF_X1 \registers_reg[26][6]  ( .D(n8299), .CK(clk), .QN(n12366) );
  DFF_X1 \registers_reg[27][6]  ( .D(n8298), .CK(clk), .QN(n12022) );
  DFF_X1 \registers_reg[28][6]  ( .D(n8297), .CK(clk), .Q(net227016), .QN(
        n15008) );
  DFF_X1 \registers_reg[29][6]  ( .D(n8296), .CK(clk), .Q(\registers[29][6] ), 
        .QN(n15808) );
  DFF_X1 \registers_reg[30][6]  ( .D(n8295), .CK(clk), .Q(\registers[30][6] ), 
        .QN(n14682) );
  DFF_X1 \registers_reg[31][6]  ( .D(n8294), .CK(clk), .Q(net227015), .QN(
        n15740) );
  DFF_X1 \registers_reg[32][6]  ( .D(n8293), .CK(clk), .QN(n12315) );
  DFF_X1 \registers_reg[33][6]  ( .D(n8292), .CK(clk), .QN(n11846) );
  DFF_X1 \registers_reg[34][6]  ( .D(n8291), .CK(clk), .Q(\registers[34][6] ), 
        .QN(n15500) );
  DFF_X1 \registers_reg[35][6]  ( .D(n8290), .CK(clk), .Q(net227014), .QN(
        n15589) );
  DFF_X1 \registers_reg[36][6]  ( .D(n8289), .CK(clk), .Q(\registers[36][6] ), 
        .QN(n15157) );
  DFF_X1 \registers_reg[37][6]  ( .D(n8288), .CK(clk), .Q(\registers[37][6] ), 
        .QN(n14369) );
  DFF_X1 \registers_reg[38][6]  ( .D(n8287), .CK(clk), .Q(\registers[38][6] ), 
        .QN(n15040) );
  DFF_X1 \registers_reg[39][6]  ( .D(n8286), .CK(clk), .QN(n12176) );
  DFF_X1 \registers_reg[40][6]  ( .D(n8285), .CK(clk), .Q(\registers[40][6] ), 
        .QN(n15082) );
  DFF_X1 \registers_reg[41][6]  ( .D(n8284), .CK(clk), .Q(\registers[41][6] ), 
        .QN(n14436) );
  DFF_X1 \registers_reg[42][6]  ( .D(n8283), .CK(clk), .Q(\registers[42][6] ), 
        .QN(n15924) );
  DFF_X1 \registers_reg[43][6]  ( .D(n8282), .CK(clk), .Q(\registers[43][6] ), 
        .QN(n14892) );
  DFF_X1 \registers_reg[44][6]  ( .D(n8281), .CK(clk), .Q(\registers[44][6] ), 
        .QN(n15470) );
  DFF_X1 \registers_reg[45][6]  ( .D(n8280), .CK(clk), .Q(\registers[45][6] ), 
        .QN(n14782) );
  DFF_X1 \registers_reg[46][6]  ( .D(n8279), .CK(clk), .QN(n11998) );
  DFF_X1 \registers_reg[47][6]  ( .D(n8278), .CK(clk), .Q(\registers[47][6] ), 
        .QN(n14551) );
  DFF_X1 \registers_reg[48][6]  ( .D(n8277), .CK(clk), .Q(\registers[48][6] ), 
        .QN(n15556) );
  DFF_X1 \registers_reg[49][6]  ( .D(n8276), .CK(clk), .Q(\registers[49][6] ), 
        .QN(n14488) );
  DFF_X1 \registers_reg[50][6]  ( .D(n8275), .CK(clk), .Q(\registers[50][6] ), 
        .QN(n15973) );
  DFF_X1 \registers_reg[51][6]  ( .D(n8274), .CK(clk), .Q(\registers[51][6] ), 
        .QN(n15403) );
  DFF_X1 \registers_reg[52][6]  ( .D(n8273), .CK(clk), .Q(net227012), .QN(
        n14942) );
  DFF_X1 \registers_reg[53][6]  ( .D(n8272), .CK(clk), .Q(net227011), .QN(
        n15916) );
  DFF_X1 \registers_reg[54][6]  ( .D(n8271), .CK(clk), .Q(\registers[54][6] ), 
        .QN(n14574) );
  DFF_X1 \registers_reg[55][6]  ( .D(n8270), .CK(clk), .Q(\registers[55][6] ), 
        .QN(n12056) );
  DFF_X1 \registers_reg[56][6]  ( .D(n8269), .CK(clk), .Q(\registers[56][6] ), 
        .QN(n16001) );
  DFF_X1 \registers_reg[57][6]  ( .D(n8268), .CK(clk), .Q(net227010), .QN(
        n15246) );
  DFF_X1 \registers_reg[58][6]  ( .D(n8267), .CK(clk), .Q(net227009), .QN(
        n14913) );
  DFF_X1 \registers_reg[59][6]  ( .D(n8266), .CK(clk), .Q(\registers[59][6] ), 
        .QN(n15435) );
  DFF_X1 \registers_reg[60][6]  ( .D(n8265), .CK(clk), .Q(\registers[60][6] ), 
        .QN(n14646) );
  DFF_X1 \registers_reg[61][6]  ( .D(n8264), .CK(clk), .Q(net227008), .QN(
        n15637) );
  DFF_X1 \registers_reg[62][6]  ( .D(n8263), .CK(clk), .Q(\registers[62][6] ), 
        .QN(n15126) );
  DFF_X1 \registers_reg[63][6]  ( .D(n8262), .CK(clk), .Q(\registers[63][6] ), 
        .QN(n14509) );
  DFF_X1 \to_mem_reg[6]  ( .D(n8261), .CK(clk), .QN(n7719) );
  DFF_X1 \registers_reg[64][6]  ( .D(n8260), .CK(clk), .Q(net227007) );
  DFF_X1 \registers_reg[65][6]  ( .D(n8259), .CK(clk), .Q(net227006) );
  DFF_X1 \registers_reg[66][6]  ( .D(n8258), .CK(clk), .Q(net227005) );
  DFF_X1 \registers_reg[67][6]  ( .D(n8257), .CK(clk), .QN(n14053) );
  DFF_X1 \registers_reg[68][6]  ( .D(n8256), .CK(clk), .Q(\registers[68][6] )
         );
  DFF_X1 \registers_reg[69][6]  ( .D(n8255), .CK(clk), .Q(net227004) );
  DFF_X1 \registers_reg[70][6]  ( .D(n8254), .CK(clk), .Q(net227003) );
  DFF_X1 \registers_reg[40][5]  ( .D(n8253), .CK(clk), .Q(\registers[40][5] ), 
        .QN(n14996) );
  DFF_X1 \registers_reg[41][5]  ( .D(n8252), .CK(clk), .Q(\registers[41][5] ), 
        .QN(n14293) );
  DFF_X1 \registers_reg[42][5]  ( .D(n8251), .CK(clk), .Q(\registers[42][5] )
         );
  DFF_X1 \registers_reg[43][5]  ( .D(n8250), .CK(clk), .Q(\registers[43][5] ), 
        .QN(n14862) );
  DFF_X1 \registers_reg[44][5]  ( .D(n8249), .CK(clk), .Q(\registers[44][5] ), 
        .QN(n15357) );
  DFF_X1 \registers_reg[45][5]  ( .D(n8248), .CK(clk), .Q(\registers[45][5] ), 
        .QN(n14642) );
  DFF_X1 \registers_reg[46][5]  ( .D(n8247), .CK(clk), .QN(n11906) );
  DFF_X1 \registers_reg[47][5]  ( .D(n8246), .CK(clk), .Q(\registers[47][5] ), 
        .QN(n14537) );
  DFF_X1 \registers_reg[48][5]  ( .D(n8245), .CK(clk), .Q(\registers[48][5] ), 
        .QN(n15360) );
  DFF_X1 \registers_reg[49][5]  ( .D(n8244), .CK(clk), .Q(\registers[49][5] ), 
        .QN(n14295) );
  DFF_X1 \registers_reg[50][5]  ( .D(n8243), .CK(clk), .Q(\registers[50][5] )
         );
  DFF_X1 \registers_reg[51][5]  ( .D(n8242), .CK(clk), .Q(\registers[51][5] ), 
        .QN(n15352) );
  DFF_X1 \registers_reg[52][5]  ( .D(n8241), .CK(clk), .Q(net227001), .QN(
        n14867) );
  DFF_X1 \registers_reg[53][5]  ( .D(n8240), .CK(clk), .Q(net227000) );
  DFF_X1 \registers_reg[54][5]  ( .D(n8239), .CK(clk), .Q(\registers[54][5] ), 
        .QN(n14539) );
  DFF_X1 \registers_reg[55][5]  ( .D(n8238), .CK(clk), .Q(\registers[55][5] ), 
        .QN(n12051) );
  DFF_X1 \registers_reg[56][5]  ( .D(n8237), .CK(clk), .Q(\registers[56][5] )
         );
  DFF_X1 \registers_reg[57][5]  ( .D(n8236), .CK(clk), .Q(net226999), .QN(
        n15242) );
  DFF_X1 \registers_reg[58][5]  ( .D(n8235), .CK(clk), .Q(net226998), .QN(
        n14865) );
  DFF_X1 \registers_reg[59][5]  ( .D(n8234), .CK(clk), .Q(\registers[59][5] ), 
        .QN(n15355) );
  DFF_X1 \registers_reg[60][5]  ( .D(n8233), .CK(clk), .Q(\registers[60][5] ), 
        .QN(n14637) );
  DFF_X1 \registers_reg[61][5]  ( .D(n8232), .CK(clk), .Q(net226997), .QN(
        n15364) );
  DFF_X1 \registers_reg[62][5]  ( .D(n8231), .CK(clk), .Q(\registers[62][5] ), 
        .QN(n14999) );
  DFF_X1 \registers_reg[63][5]  ( .D(n8230), .CK(clk), .Q(\registers[63][5] ), 
        .QN(n14298) );
  DFF_X1 \registers_reg[0][5]  ( .D(n8229), .CK(clk), .Q(\registers[0][5] ), 
        .QN(n15800) );
  DFF_X1 \registers_reg[1][5]  ( .D(n8228), .CK(clk), .Q(\registers[1][5] ), 
        .QN(n15584) );
  DFF_X1 \registers_reg[2][5]  ( .D(n8227), .CK(clk), .Q(\registers[2][5] ), 
        .QN(n14780) );
  DFF_X1 \registers_reg[3][5]  ( .D(n8226), .CK(clk), .Q(net226996), .QN(
        n15763) );
  DFF_X1 \registers_reg[4][5]  ( .D(n8225), .CK(clk), .Q(\registers[4][5] ), 
        .QN(n15526) );
  DFF_X1 \registers_reg[5][5]  ( .D(n8224), .CK(clk), .Q(\registers[5][5] ), 
        .QN(n14720) );
  DFF_X1 \registers_reg[6][5]  ( .D(n8223), .CK(clk), .QN(n12365) );
  DFF_X1 \registers_reg[7][5]  ( .D(n8222), .CK(clk), .Q(\registers[7][5] ), 
        .QN(n15331) );
  DFF_X1 \registers_reg[8][5]  ( .D(n8221), .CK(clk), .Q(net226995), .QN(
        n15214) );
  DFF_X1 \registers_reg[9][5]  ( .D(n8220), .CK(clk), .Q(\registers[9][5] ), 
        .QN(n14333) );
  DFF_X1 \registers_reg[10][5]  ( .D(n8219), .CK(clk), .Q(\registers[10][5] ), 
        .QN(n14721) );
  DFF_X1 \registers_reg[11][5]  ( .D(n8218), .CK(clk), .Q(\registers[11][5] ), 
        .QN(n14434) );
  DFF_X1 \registers_reg[12][5]  ( .D(n8217), .CK(clk), .Q(\registers[12][5] ), 
        .QN(n15673) );
  DFF_X1 \registers_reg[13][5]  ( .D(n8216), .CK(clk), .Q(net226994), .QN(
        n15080) );
  DFF_X1 \registers_reg[14][5]  ( .D(n8215), .CK(clk), .QN(n11885) );
  DFF_X1 \registers_reg[15][5]  ( .D(n8214), .CK(clk), .Q(\registers[15][5] ), 
        .QN(n15296) );
  DFF_X1 \registers_reg[16][5]  ( .D(n8213), .CK(clk), .Q(\registers[16][5] ), 
        .QN(n15703) );
  DFF_X1 \registers_reg[17][5]  ( .D(n8212), .CK(clk), .Q(\registers[17][5] ), 
        .QN(n14609) );
  DFF_X1 \registers_reg[18][5]  ( .D(n8211), .CK(clk), .Q(\registers[18][5] ), 
        .QN(n14368) );
  DFF_X1 \registers_reg[19][5]  ( .D(n8210), .CK(clk), .Q(\registers[19][5] ), 
        .QN(n15807) );
  DFF_X1 \registers_reg[20][5]  ( .D(n8209), .CK(clk), .QN(n14835) );
  DFF_X1 \registers_reg[21][5]  ( .D(n8208), .CK(clk), .QN(n12209) );
  DFF_X1 \registers_reg[22][5]  ( .D(n8207), .CK(clk), .Q(\registers[22][5] ), 
        .QN(n15375) );
  DFF_X1 \registers_reg[23][5]  ( .D(n8206), .CK(clk), .Q(\registers[23][5] ), 
        .QN(n15885) );
  DFF_X1 \registers_reg[24][5]  ( .D(n8205), .CK(clk), .Q(net226993), .QN(
        n15184) );
  DFF_X1 \registers_reg[25][5]  ( .D(n8204), .CK(clk), .Q(\registers[25][5] ), 
        .QN(n14303) );
  DFF_X1 \registers_reg[26][5]  ( .D(n8203), .CK(clk), .QN(n12364) );
  DFF_X1 \registers_reg[27][5]  ( .D(n8202), .CK(clk), .QN(n12021) );
  DFF_X1 \registers_reg[28][5]  ( .D(n8201), .CK(clk), .Q(net226992), .QN(
        n15007) );
  DFF_X1 \registers_reg[29][5]  ( .D(n8200), .CK(clk), .Q(\registers[29][5] ), 
        .QN(n15806) );
  DFF_X1 \registers_reg[30][5]  ( .D(n8199), .CK(clk), .Q(\registers[30][5] ), 
        .QN(n14681) );
  DFF_X1 \registers_reg[31][5]  ( .D(n8198), .CK(clk), .Q(net226991), .QN(
        n15739) );
  DFF_X1 \registers_reg[32][5]  ( .D(n8197), .CK(clk), .QN(n12308) );
  DFF_X1 \registers_reg[33][5]  ( .D(n8196), .CK(clk), .QN(n11584) );
  DFF_X1 \registers_reg[34][5]  ( .D(n8195), .CK(clk), .Q(\registers[34][5] ), 
        .QN(n15358) );
  DFF_X1 \registers_reg[35][5]  ( .D(n8194), .CK(clk), .Q(net226990), .QN(
        n15363) );
  DFF_X1 \registers_reg[36][5]  ( .D(n8193), .CK(clk), .Q(\registers[36][5] ), 
        .QN(n15000) );
  DFF_X1 \registers_reg[37][5]  ( .D(n8192), .CK(clk), .Q(\registers[37][5] ), 
        .QN(n14290) );
  DFF_X1 \registers_reg[38][5]  ( .D(n8191), .CK(clk), .Q(\registers[38][5] ), 
        .QN(n14993) );
  DFF_X1 \registers_reg[39][5]  ( .D(n8190), .CK(clk), .QN(n12162) );
  DFF_X1 \to_mem_reg[5]  ( .D(n8189), .CK(clk), .QN(n7720) );
  DFF_X1 \registers_reg[64][5]  ( .D(n8188), .CK(clk), .Q(net226989), .QN(
        n16125) );
  DFF_X1 \registers_reg[65][5]  ( .D(n8187), .CK(clk), .Q(net226988), .QN(
        n16087) );
  DFF_X1 \registers_reg[66][5]  ( .D(n8186), .CK(clk), .Q(net226987), .QN(
        n16041) );
  DFF_X1 \registers_reg[67][5]  ( .D(n8185), .CK(clk), .QN(n14212) );
  DFF_X1 \registers_reg[68][5]  ( .D(n8184), .CK(clk), .Q(\registers[68][5] ), 
        .QN(n16175) );
  DFF_X1 \registers_reg[69][5]  ( .D(n8183), .CK(clk), .Q(net226986), .QN(
        n16127) );
  DFF_X1 \registers_reg[70][5]  ( .D(n8182), .CK(clk), .Q(net226985), .QN(
        n16037) );
  DFF_X1 \registers_reg[24][4]  ( .D(n8181), .CK(clk), .Q(net226984), .QN(
        n15002) );
  DFF_X1 \registers_reg[25][4]  ( .D(n8180), .CK(clk), .Q(\registers[25][4] ), 
        .QN(n14283) );
  DFF_X1 \registers_reg[26][4]  ( .D(n8179), .CK(clk), .QN(n12341) );
  DFF_X1 \registers_reg[27][4]  ( .D(n8178), .CK(clk), .QN(n12017) );
  DFF_X1 \registers_reg[28][4]  ( .D(n8177), .CK(clk), .Q(net226983), .QN(
        n14990) );
  DFF_X1 \registers_reg[29][4]  ( .D(n8176), .CK(clk), .Q(\registers[29][4] )
         );
  DFF_X1 \registers_reg[30][4]  ( .D(n8175), .CK(clk), .Q(\registers[30][4] ), 
        .QN(n14639) );
  DFF_X1 \registers_reg[31][4]  ( .D(n8174), .CK(clk), .Q(net226982), .QN(
        n15368) );
  DFF_X1 \registers_reg[48][4]  ( .D(n8173), .CK(clk), .Q(\registers[48][4] ), 
        .QN(n15359) );
  DFF_X1 \registers_reg[49][4]  ( .D(n8172), .CK(clk), .Q(\registers[49][4] ), 
        .QN(n14294) );
  DFF_X1 \registers_reg[50][4]  ( .D(n8171), .CK(clk), .Q(\registers[50][4] )
         );
  DFF_X1 \registers_reg[51][4]  ( .D(n8170), .CK(clk), .Q(\registers[51][4] ), 
        .QN(n15351) );
  DFF_X1 \registers_reg[52][4]  ( .D(n8169), .CK(clk), .Q(net226981), .QN(
        n14866) );
  DFF_X1 \registers_reg[53][4]  ( .D(n8168), .CK(clk), .Q(net226980) );
  DFF_X1 \registers_reg[54][4]  ( .D(n8167), .CK(clk), .Q(\registers[54][4] ), 
        .QN(n14538) );
  DFF_X1 \registers_reg[55][4]  ( .D(n8166), .CK(clk), .Q(\registers[55][4] ), 
        .QN(n12050) );
  DFF_X1 \registers_reg[56][4]  ( .D(n8165), .CK(clk), .Q(\registers[56][4] )
         );
  DFF_X1 \registers_reg[57][4]  ( .D(n8164), .CK(clk), .Q(net226979), .QN(
        n15241) );
  DFF_X1 \registers_reg[58][4]  ( .D(n8163), .CK(clk), .Q(net226978), .QN(
        n14864) );
  DFF_X1 \registers_reg[59][4]  ( .D(n8162), .CK(clk), .Q(\registers[59][4] ), 
        .QN(n15354) );
  DFF_X1 \registers_reg[60][4]  ( .D(n8161), .CK(clk), .Q(\registers[60][4] ), 
        .QN(n14636) );
  DFF_X1 \registers_reg[61][4]  ( .D(n8160), .CK(clk), .Q(net226977), .QN(
        n15362) );
  DFF_X1 \registers_reg[62][4]  ( .D(n8159), .CK(clk), .Q(\registers[62][4] ), 
        .QN(n14998) );
  DFF_X1 \registers_reg[63][4]  ( .D(n8158), .CK(clk), .Q(\registers[63][4] ), 
        .QN(n14297) );
  DFF_X1 \registers_reg[0][4]  ( .D(n8157), .CK(clk), .Q(\registers[0][4] ), 
        .QN(n15799) );
  DFF_X1 \registers_reg[1][4]  ( .D(n8156), .CK(clk), .Q(\registers[1][4] ), 
        .QN(n15583) );
  DFF_X1 \registers_reg[2][4]  ( .D(n8155), .CK(clk), .Q(\registers[2][4] ), 
        .QN(n14778) );
  DFF_X1 \registers_reg[3][4]  ( .D(n8154), .CK(clk), .Q(net226976), .QN(
        n15762) );
  DFF_X1 \registers_reg[4][4]  ( .D(n8153), .CK(clk), .Q(\registers[4][4] ), 
        .QN(n15525) );
  DFF_X1 \registers_reg[5][4]  ( .D(n8152), .CK(clk), .Q(\registers[5][4] ), 
        .QN(n14718) );
  DFF_X1 \registers_reg[6][4]  ( .D(n8151), .CK(clk), .QN(n12363) );
  DFF_X1 \registers_reg[7][4]  ( .D(n8150), .CK(clk), .Q(\registers[7][4] ), 
        .QN(n15330) );
  DFF_X1 \registers_reg[8][4]  ( .D(n8149), .CK(clk), .Q(net226975), .QN(
        n15213) );
  DFF_X1 \registers_reg[9][4]  ( .D(n8148), .CK(clk), .Q(\registers[9][4] ), 
        .QN(n14332) );
  DFF_X1 \registers_reg[10][4]  ( .D(n8147), .CK(clk), .Q(\registers[10][4] ), 
        .QN(n14719) );
  DFF_X1 \registers_reg[11][4]  ( .D(n8146), .CK(clk), .Q(\registers[11][4] ), 
        .QN(n14432) );
  DFF_X1 \registers_reg[12][4]  ( .D(n8145), .CK(clk), .Q(\registers[12][4] ), 
        .QN(n15672) );
  DFF_X1 \registers_reg[13][4]  ( .D(n8144), .CK(clk), .Q(net226974), .QN(
        n15078) );
  DFF_X1 \registers_reg[14][4]  ( .D(n8143), .CK(clk), .QN(n11884) );
  DFF_X1 \registers_reg[15][4]  ( .D(n8142), .CK(clk), .Q(\registers[15][4] ), 
        .QN(n15295) );
  DFF_X1 \registers_reg[16][4]  ( .D(n8141), .CK(clk), .Q(\registers[16][4] ), 
        .QN(n15366) );
  DFF_X1 \registers_reg[17][4]  ( .D(n8140), .CK(clk), .Q(\registers[17][4] ), 
        .QN(n14569) );
  DFF_X1 \registers_reg[18][4]  ( .D(n8139), .CK(clk), .Q(\registers[18][4] ), 
        .QN(n14289) );
  DFF_X1 \registers_reg[19][4]  ( .D(n8138), .CK(clk), .Q(\registers[19][4] )
         );
  DFF_X1 \registers_reg[20][4]  ( .D(n8137), .CK(clk), .QN(n14823) );
  DFF_X1 \registers_reg[21][4]  ( .D(n8136), .CK(clk), .QN(n12195) );
  DFF_X1 \registers_reg[22][4]  ( .D(n8135), .CK(clk), .Q(\registers[22][4] ), 
        .QN(n15350) );
  DFF_X1 \registers_reg[23][4]  ( .D(n8134), .CK(clk), .Q(\registers[23][4] )
         );
  DFF_X1 \registers_reg[32][4]  ( .D(n8133), .CK(clk), .QN(n12313) );
  DFF_X1 \registers_reg[33][4]  ( .D(n8132), .CK(clk), .QN(n11844) );
  DFF_X1 \registers_reg[34][4]  ( .D(n8131), .CK(clk), .Q(\registers[34][4] ), 
        .QN(n15499) );
  DFF_X1 \registers_reg[35][4]  ( .D(n8130), .CK(clk), .Q(net226973), .QN(
        n15588) );
  DFF_X1 \registers_reg[36][4]  ( .D(n8129), .CK(clk), .Q(\registers[36][4] ), 
        .QN(n15155) );
  DFF_X1 \registers_reg[37][4]  ( .D(n8128), .CK(clk), .Q(\registers[37][4] ), 
        .QN(n14367) );
  DFF_X1 \registers_reg[38][4]  ( .D(n8127), .CK(clk), .Q(\registers[38][4] ), 
        .QN(n15039) );
  DFF_X1 \registers_reg[39][4]  ( .D(n8126), .CK(clk), .QN(n12175) );
  DFF_X1 \registers_reg[40][4]  ( .D(n8125), .CK(clk), .Q(\registers[40][4] ), 
        .QN(n15079) );
  DFF_X1 \registers_reg[41][4]  ( .D(n8124), .CK(clk), .Q(\registers[41][4] ), 
        .QN(n14433) );
  DFF_X1 \registers_reg[42][4]  ( .D(n8123), .CK(clk), .Q(\registers[42][4] ), 
        .QN(n15923) );
  DFF_X1 \registers_reg[43][4]  ( .D(n8122), .CK(clk), .Q(\registers[43][4] ), 
        .QN(n14891) );
  DFF_X1 \registers_reg[44][4]  ( .D(n8121), .CK(clk), .Q(\registers[44][4] ), 
        .QN(n15469) );
  DFF_X1 \registers_reg[45][4]  ( .D(n8120), .CK(clk), .Q(\registers[45][4] ), 
        .QN(n14779) );
  DFF_X1 \registers_reg[46][4]  ( .D(n8119), .CK(clk), .QN(n11997) );
  DFF_X1 \registers_reg[47][4]  ( .D(n8118), .CK(clk), .Q(\registers[47][4] ), 
        .QN(n14550) );
  DFF_X1 \to_mem_reg[4]  ( .D(n8117), .CK(clk), .QN(n7721) );
  DFF_X1 \registers_reg[64][4]  ( .D(n8116), .CK(clk), .Q(net226971), .QN(
        n16124) );
  DFF_X1 \registers_reg[65][4]  ( .D(n8115), .CK(clk), .Q(net226970), .QN(
        n16086) );
  DFF_X1 \registers_reg[66][4]  ( .D(n8114), .CK(clk), .Q(net226969), .QN(
        n16040) );
  DFF_X1 \registers_reg[67][4]  ( .D(n8113), .CK(clk), .QN(n14071) );
  DFF_X1 \registers_reg[68][4]  ( .D(n8112), .CK(clk), .Q(\registers[68][4] ), 
        .QN(n16174) );
  DFF_X1 \registers_reg[69][4]  ( .D(n8111), .CK(clk), .Q(net226968), .QN(
        n16126) );
  DFF_X1 \registers_reg[70][4]  ( .D(n8110), .CK(clk), .Q(net226967), .QN(
        n16036) );
  DFF_X1 \registers_reg[71][31]  ( .D(n8109), .CK(clk), .QN(n14051) );
  DFF_X1 \out1_reg[31]  ( .D(n8108), .CK(clk), .Q(out1[31]), .QN(net226965) );
  DFF_X1 \registers_reg[71][30]  ( .D(n8107), .CK(clk), .QN(n14860) );
  DFF_X1 \out1_reg[30]  ( .D(n8106), .CK(clk), .Q(out1[30]), .QN(net226963) );
  DFF_X1 \registers_reg[71][29]  ( .D(n8105), .CK(clk), .QN(n14988) );
  DFF_X1 \out1_reg[29]  ( .D(n8104), .CK(clk), .Q(out1[29]), .QN(net226961) );
  DFF_X1 \registers_reg[71][28]  ( .D(n8103), .CK(clk), .QN(n14987) );
  DFF_X1 \out1_reg[28]  ( .D(n8102), .CK(clk), .Q(out1[28]), .QN(net226959) );
  DFF_X1 \registers_reg[71][27]  ( .D(n8101), .CK(clk), .QN(n14986) );
  DFF_X1 \out1_reg[27]  ( .D(n8100), .CK(clk), .Q(out1[27]), .QN(net226957) );
  DFF_X1 \registers_reg[71][26]  ( .D(n8099), .CK(clk), .QN(n14985) );
  DFF_X1 \out1_reg[26]  ( .D(n8098), .CK(clk), .Q(out1[26]), .QN(net226955) );
  DFF_X1 \registers_reg[71][25]  ( .D(n8097), .CK(clk), .QN(n14984) );
  DFF_X1 \out1_reg[25]  ( .D(n8096), .CK(clk), .Q(out1[25]), .QN(net226953) );
  DFF_X1 \registers_reg[71][24]  ( .D(n8095), .CK(clk), .QN(n14983) );
  DFF_X1 \out1_reg[24]  ( .D(n8094), .CK(clk), .Q(out1[24]), .QN(net226951) );
  DFF_X1 \registers_reg[71][23]  ( .D(n8093), .CK(clk), .QN(n14979) );
  DFF_X1 \out1_reg[23]  ( .D(n8092), .CK(clk), .Q(out1[23]), .QN(net226949) );
  DFF_X1 \registers_reg[71][22]  ( .D(n8091), .CK(clk), .QN(n14982) );
  DFF_X1 \out1_reg[22]  ( .D(n8090), .CK(clk), .Q(out1[22]), .QN(net226947) );
  DFF_X1 \registers_reg[71][21]  ( .D(n8089), .CK(clk), .QN(n14981) );
  DFF_X1 \out1_reg[21]  ( .D(n8088), .CK(clk), .Q(out1[21]), .QN(net226945) );
  DFF_X1 \registers_reg[71][20]  ( .D(n8087), .CK(clk), .QN(n14978) );
  DFF_X1 \out1_reg[20]  ( .D(n8086), .CK(clk), .Q(out1[20]), .QN(net226943) );
  DFF_X1 \registers_reg[71][19]  ( .D(n8085), .CK(clk), .QN(n14977) );
  DFF_X1 \out1_reg[19]  ( .D(n8084), .CK(clk), .Q(out1[19]), .QN(net226941) );
  DFF_X1 \registers_reg[71][18]  ( .D(n8083), .CK(clk), .QN(n14976) );
  DFF_X1 \out1_reg[18]  ( .D(n8082), .CK(clk), .Q(out1[18]), .QN(net226939) );
  DFF_X1 \registers_reg[71][17]  ( .D(n8081), .CK(clk), .QN(n14975) );
  DFF_X1 \out1_reg[17]  ( .D(n8080), .CK(clk), .Q(out1[17]), .QN(net226937) );
  DFF_X1 \registers_reg[71][16]  ( .D(n8079), .CK(clk), .QN(n14974) );
  DFF_X1 \out1_reg[16]  ( .D(n8078), .CK(clk), .Q(out1[16]), .QN(net226935) );
  DFF_X1 \registers_reg[71][15]  ( .D(n8077), .CK(clk), .QN(n14973) );
  DFF_X1 \out1_reg[15]  ( .D(n8076), .CK(clk), .Q(out1[15]), .QN(net226933) );
  DFF_X1 \registers_reg[71][14]  ( .D(n8075), .CK(clk), .QN(n14972) );
  DFF_X1 \out1_reg[14]  ( .D(n8074), .CK(clk), .Q(out1[14]), .QN(net226931) );
  DFF_X1 \registers_reg[71][13]  ( .D(n8073), .CK(clk), .QN(n14971) );
  DFF_X1 \out1_reg[13]  ( .D(n8072), .CK(clk), .Q(out1[13]), .QN(net226929) );
  DFF_X1 \registers_reg[71][12]  ( .D(n8071), .CK(clk), .QN(n14970) );
  DFF_X1 \out1_reg[12]  ( .D(n8070), .CK(clk), .Q(out1[12]), .QN(net226927) );
  DFF_X1 \registers_reg[71][11]  ( .D(n8069), .CK(clk), .QN(n14969) );
  DFF_X1 \out1_reg[11]  ( .D(n8068), .CK(clk), .Q(out1[11]), .QN(net226925) );
  DFF_X1 \registers_reg[71][10]  ( .D(n8067), .CK(clk), .QN(n14968) );
  DFF_X1 \out1_reg[10]  ( .D(n8066), .CK(clk), .Q(out1[10]), .QN(net226923) );
  DFF_X1 \registers_reg[71][9]  ( .D(n8065), .CK(clk), .QN(n14967) );
  DFF_X1 \out1_reg[9]  ( .D(n8064), .CK(clk), .Q(out1[9]), .QN(net226921) );
  DFF_X1 \registers_reg[71][8]  ( .D(n8063), .CK(clk), .QN(n14966) );
  DFF_X1 \out1_reg[8]  ( .D(n8062), .CK(clk), .Q(out1[8]), .QN(net226919) );
  DFF_X1 \registers_reg[71][7]  ( .D(n8061), .CK(clk), .QN(n14965) );
  DFF_X1 \out1_reg[7]  ( .D(n8060), .CK(clk), .Q(out1[7]), .QN(net226917) );
  DFF_X1 \registers_reg[71][6]  ( .D(n8059), .CK(clk), .QN(n14868) );
  DFF_X1 \out1_reg[6]  ( .D(n8058), .CK(clk), .Q(out1[6]), .QN(net226915) );
  DFF_X1 \registers_reg[71][5]  ( .D(n8057), .CK(clk), .QN(n14964) );
  DFF_X1 \out1_reg[5]  ( .D(n8056), .CK(clk), .Q(out1[5]), .QN(net226913) );
  DFF_X1 \registers_reg[71][4]  ( .D(n8055), .CK(clk), .QN(n14963) );
  DFF_X1 \out1_reg[4]  ( .D(n8054), .CK(clk), .Q(out1[4]), .QN(net226911) );
  DFF_X1 \registers_reg[24][3]  ( .D(n8053), .CK(clk), .Q(net226910), .QN(
        n15001) );
  DFF_X1 \registers_reg[25][3]  ( .D(n8052), .CK(clk), .Q(\registers[25][3] ), 
        .QN(n14282) );
  DFF_X1 \registers_reg[26][3]  ( .D(n8051), .CK(clk), .QN(n12340) );
  DFF_X1 \registers_reg[27][3]  ( .D(n8050), .CK(clk), .QN(n12016) );
  DFF_X1 \registers_reg[28][3]  ( .D(n8049), .CK(clk), .Q(net226909), .QN(
        n14989) );
  DFF_X1 \registers_reg[29][3]  ( .D(n8048), .CK(clk), .Q(\registers[29][3] )
         );
  DFF_X1 \registers_reg[30][3]  ( .D(n8047), .CK(clk), .Q(\registers[30][3] ), 
        .QN(n14638) );
  DFF_X1 \registers_reg[31][3]  ( .D(n8046), .CK(clk), .Q(net226908), .QN(
        n15367) );
  DFF_X1 \registers_reg[40][3]  ( .D(n8045), .CK(clk), .Q(\registers[40][3] ), 
        .QN(n14995) );
  DFF_X1 \registers_reg[41][3]  ( .D(n8044), .CK(clk), .Q(\registers[41][3] ), 
        .QN(n14292) );
  DFF_X1 \registers_reg[42][3]  ( .D(n8043), .CK(clk), .Q(\registers[42][3] )
         );
  DFF_X1 \registers_reg[43][3]  ( .D(n8042), .CK(clk), .Q(\registers[43][3] ), 
        .QN(n14861) );
  DFF_X1 \registers_reg[44][3]  ( .D(n8041), .CK(clk), .Q(\registers[44][3] ), 
        .QN(n15356) );
  DFF_X1 \registers_reg[45][3]  ( .D(n8040), .CK(clk), .Q(\registers[45][3] ), 
        .QN(n14641) );
  DFF_X1 \registers_reg[46][3]  ( .D(n8039), .CK(clk), .QN(n11905) );
  DFF_X1 \registers_reg[47][3]  ( .D(n8038), .CK(clk), .Q(\registers[47][3] ), 
        .QN(n14536) );
  DFF_X1 \registers_reg[56][3]  ( .D(n8037), .CK(clk), .Q(\registers[56][3] )
         );
  DFF_X1 \registers_reg[57][3]  ( .D(n8036), .CK(clk), .Q(net226906), .QN(
        n15240) );
  DFF_X1 \registers_reg[58][3]  ( .D(n8035), .CK(clk), .Q(net226905), .QN(
        n14863) );
  DFF_X1 \registers_reg[59][3]  ( .D(n8034), .CK(clk), .Q(\registers[59][3] ), 
        .QN(n15353) );
  DFF_X1 \registers_reg[60][3]  ( .D(n8033), .CK(clk), .Q(\registers[60][3] ), 
        .QN(n14635) );
  DFF_X1 \registers_reg[61][3]  ( .D(n8032), .CK(clk), .Q(net226904), .QN(
        n15361) );
  DFF_X1 \registers_reg[62][3]  ( .D(n8031), .CK(clk), .Q(\registers[62][3] ), 
        .QN(n14997) );
  DFF_X1 \registers_reg[63][3]  ( .D(n8030), .CK(clk), .Q(\registers[63][3] ), 
        .QN(n14296) );
  DFF_X1 \registers_reg[0][3]  ( .D(n8029), .CK(clk), .Q(\registers[0][3] ), 
        .QN(n15798) );
  DFF_X1 \registers_reg[1][3]  ( .D(n8028), .CK(clk), .Q(\registers[1][3] ), 
        .QN(n15582) );
  DFF_X1 \registers_reg[2][3]  ( .D(n8027), .CK(clk), .Q(\registers[2][3] ), 
        .QN(n14777) );
  DFF_X1 \registers_reg[3][3]  ( .D(n8026), .CK(clk), .Q(net226903), .QN(
        n15761) );
  DFF_X1 \registers_reg[4][3]  ( .D(n8025), .CK(clk), .Q(\registers[4][3] ), 
        .QN(n15524) );
  DFF_X1 \registers_reg[5][3]  ( .D(n8024), .CK(clk), .Q(\registers[5][3] ), 
        .QN(n14717) );
  DFF_X1 \registers_reg[6][3]  ( .D(n8023), .CK(clk), .QN(n12362) );
  DFF_X1 \registers_reg[7][3]  ( .D(n8022), .CK(clk), .Q(\registers[7][3] ), 
        .QN(n15329) );
  DFF_X1 \registers_reg[8][3]  ( .D(n8021), .CK(clk), .Q(net226902), .QN(
        n15003) );
  DFF_X1 \registers_reg[9][3]  ( .D(n8020), .CK(clk), .Q(\registers[9][3] ), 
        .QN(n14288) );
  DFF_X1 \registers_reg[10][3]  ( .D(n8019), .CK(clk), .Q(\registers[10][3] ), 
        .QN(n14640) );
  DFF_X1 \registers_reg[11][3]  ( .D(n8018), .CK(clk), .Q(\registers[11][3] ), 
        .QN(n14291) );
  DFF_X1 \registers_reg[12][3]  ( .D(n8017), .CK(clk), .Q(\registers[12][3] ), 
        .QN(n15365) );
  DFF_X1 \registers_reg[13][3]  ( .D(n8016), .CK(clk), .Q(net226901), .QN(
        n14994) );
  DFF_X1 \registers_reg[14][3]  ( .D(n8015), .CK(clk), .QN(n11627) );
  DFF_X1 \registers_reg[15][3]  ( .D(n8014), .CK(clk), .Q(\registers[15][3] ), 
        .QN(n15284) );
  DFF_X1 \registers_reg[16][3]  ( .D(n8013), .CK(clk), .Q(\registers[16][3] ), 
        .QN(n15702) );
  DFF_X1 \registers_reg[17][3]  ( .D(n8012), .CK(clk), .Q(\registers[17][3] ), 
        .QN(n14608) );
  DFF_X1 \registers_reg[18][3]  ( .D(n8011), .CK(clk), .Q(\registers[18][3] ), 
        .QN(n14366) );
  DFF_X1 \registers_reg[19][3]  ( .D(n8010), .CK(clk), .Q(\registers[19][3] ), 
        .QN(n15805) );
  DFF_X1 \registers_reg[20][3]  ( .D(n8009), .CK(clk), .QN(n14834) );
  DFF_X1 \registers_reg[21][3]  ( .D(n8008), .CK(clk), .QN(n12208) );
  DFF_X1 \registers_reg[22][3]  ( .D(n8007), .CK(clk), .Q(\registers[22][3] ), 
        .QN(n15374) );
  DFF_X1 \registers_reg[23][3]  ( .D(n8006), .CK(clk), .Q(\registers[23][3] ), 
        .QN(n15884) );
  DFF_X1 \registers_reg[32][3]  ( .D(n8005), .CK(clk), .QN(n12312) );
  DFF_X1 \registers_reg[33][3]  ( .D(n8004), .CK(clk), .QN(n11842) );
  DFF_X1 \registers_reg[34][3]  ( .D(n8003), .CK(clk), .Q(\registers[34][3] ), 
        .QN(n15498) );
  DFF_X1 \registers_reg[35][3]  ( .D(n8002), .CK(clk), .Q(net226900), .QN(
        n15587) );
  DFF_X1 \registers_reg[36][3]  ( .D(n8001), .CK(clk), .Q(\registers[36][3] ), 
        .QN(n15154) );
  DFF_X1 \registers_reg[37][3]  ( .D(n8000), .CK(clk), .Q(\registers[37][3] ), 
        .QN(n14365) );
  DFF_X1 \registers_reg[38][3]  ( .D(n7999), .CK(clk), .Q(\registers[38][3] ), 
        .QN(n15038) );
  DFF_X1 \registers_reg[39][3]  ( .D(n7998), .CK(clk), .QN(n12174) );
  DFF_X1 \registers_reg[48][3]  ( .D(n7997), .CK(clk), .Q(\registers[48][3] ), 
        .QN(n15555) );
  DFF_X1 \registers_reg[49][3]  ( .D(n7996), .CK(clk), .Q(\registers[49][3] ), 
        .QN(n14487) );
  DFF_X1 \registers_reg[50][3]  ( .D(n7995), .CK(clk), .Q(\registers[50][3] ), 
        .QN(n15972) );
  DFF_X1 \registers_reg[51][3]  ( .D(n7994), .CK(clk), .Q(\registers[51][3] ), 
        .QN(n15402) );
  DFF_X1 \registers_reg[52][3]  ( .D(n7993), .CK(clk), .Q(net226899), .QN(
        n14941) );
  DFF_X1 \registers_reg[53][3]  ( .D(n7992), .CK(clk), .Q(net226898), .QN(
        n15915) );
  DFF_X1 \registers_reg[54][3]  ( .D(n7991), .CK(clk), .Q(\registers[54][3] ), 
        .QN(n14572) );
  DFF_X1 \registers_reg[55][3]  ( .D(n7990), .CK(clk), .Q(\registers[55][3] ), 
        .QN(n12054) );
  DFF_X1 \to_mem_reg[3]  ( .D(n7989), .CK(clk), .QN(n7722) );
  DFF_X1 \registers_reg[64][3]  ( .D(n7988), .CK(clk), .Q(net226897), .QN(
        n16204) );
  DFF_X1 \registers_reg[65][3]  ( .D(n7987), .CK(clk), .Q(net226896), .QN(
        n16114) );
  DFF_X1 \registers_reg[66][3]  ( .D(n7986), .CK(clk), .Q(net226895), .QN(
        n16122) );
  DFF_X1 \registers_reg[67][3]  ( .D(n7985), .CK(clk), .QN(n14287) );
  DFF_X1 \registers_reg[68][3]  ( .D(n7984), .CK(clk), .Q(\registers[68][3] ), 
        .QN(n16210) );
  DFF_X1 \registers_reg[69][3]  ( .D(n7983), .CK(clk), .Q(net226894), .QN(
        n16206) );
  DFF_X1 \registers_reg[70][3]  ( .D(n7982), .CK(clk), .Q(net226893), .QN(
        n16119) );
  DFF_X1 \registers_reg[71][3]  ( .D(n7981), .CK(clk), .QN(n14980) );
  DFF_X1 \out1_reg[3]  ( .D(n7980), .CK(clk), .Q(out1[3]), .QN(net226891) );
  DFF_X1 \registers_reg[4][2]  ( .D(n7979), .CK(clk), .Q(\registers[4][2] ), 
        .QN(n15523) );
  DFF_X1 \registers_reg[5][2]  ( .D(n7978), .CK(clk), .Q(\registers[5][2] ), 
        .QN(n14715) );
  DFF_X1 \registers_reg[6][2]  ( .D(n7977), .CK(clk), .QN(n12361) );
  DFF_X1 \registers_reg[7][2]  ( .D(n7976), .CK(clk), .Q(\registers[7][2] ), 
        .QN(n15328) );
  DFF_X1 \registers_reg[12][2]  ( .D(n7975), .CK(clk), .Q(\registers[12][2] ), 
        .QN(n15671) );
  DFF_X1 \registers_reg[13][2]  ( .D(n7974), .CK(clk), .Q(net226890), .QN(
        n15076) );
  DFF_X1 \registers_reg[14][2]  ( .D(n7973), .CK(clk), .QN(n11883) );
  DFF_X1 \registers_reg[15][2]  ( .D(n7972), .CK(clk), .Q(\registers[15][2] ), 
        .QN(n15294) );
  DFF_X1 \registers_reg[20][2]  ( .D(n7971), .CK(clk), .QN(n14833) );
  DFF_X1 \registers_reg[21][2]  ( .D(n7970), .CK(clk), .QN(n12207) );
  DFF_X1 \registers_reg[22][2]  ( .D(n7969), .CK(clk), .Q(\registers[22][2] ), 
        .QN(n15372) );
  DFF_X1 \registers_reg[23][2]  ( .D(n7968), .CK(clk), .Q(\registers[23][2] ), 
        .QN(n15883) );
  DFF_X1 \registers_reg[28][2]  ( .D(n7967), .CK(clk), .Q(net226889), .QN(
        n15006) );
  DFF_X1 \registers_reg[29][2]  ( .D(n7966), .CK(clk), .Q(\registers[29][2] ), 
        .QN(n15794) );
  DFF_X1 \registers_reg[30][2]  ( .D(n7965), .CK(clk), .Q(\registers[30][2] ), 
        .QN(n14680) );
  DFF_X1 \registers_reg[31][2]  ( .D(n7964), .CK(clk), .Q(net226888), .QN(
        n15738) );
  DFF_X1 \registers_reg[36][2]  ( .D(n7963), .CK(clk), .Q(\registers[36][2] ), 
        .QN(n15151) );
  DFF_X1 \registers_reg[37][2]  ( .D(n7962), .CK(clk), .Q(\registers[37][2] ), 
        .QN(n14361) );
  DFF_X1 \registers_reg[38][2]  ( .D(n7961), .CK(clk), .Q(\registers[38][2] ), 
        .QN(n15036) );
  DFF_X1 \registers_reg[39][2]  ( .D(n7960), .CK(clk), .QN(n12173) );
  DFF_X1 \registers_reg[44][2]  ( .D(n7959), .CK(clk), .Q(\registers[44][2] ), 
        .QN(n15468) );
  DFF_X1 \registers_reg[45][2]  ( .D(n7958), .CK(clk), .Q(\registers[45][2] ), 
        .QN(n14776) );
  DFF_X1 \registers_reg[46][2]  ( .D(n7957), .CK(clk), .QN(n11995) );
  DFF_X1 \registers_reg[47][2]  ( .D(n7956), .CK(clk), .Q(\registers[47][2] ), 
        .QN(n14549) );
  DFF_X1 \registers_reg[52][2]  ( .D(n7955), .CK(clk), .Q(net226886), .QN(
        n14940) );
  DFF_X1 \registers_reg[53][2]  ( .D(n7954), .CK(clk), .Q(net226885), .QN(
        n15913) );
  DFF_X1 \registers_reg[54][2]  ( .D(n7953), .CK(clk), .Q(\registers[54][2] ), 
        .QN(n14571) );
  DFF_X1 \registers_reg[55][2]  ( .D(n7952), .CK(clk), .Q(\registers[55][2] ), 
        .QN(n12053) );
  DFF_X1 \registers_reg[60][2]  ( .D(n7951), .CK(clk), .Q(\registers[60][2] ), 
        .QN(n14643) );
  DFF_X1 \registers_reg[61][2]  ( .D(n7950), .CK(clk), .Q(net226884), .QN(
        n15578) );
  DFF_X1 \registers_reg[62][2]  ( .D(n7949), .CK(clk), .Q(\registers[62][2] ), 
        .QN(n15125) );
  DFF_X1 \registers_reg[63][2]  ( .D(n7948), .CK(clk), .Q(\registers[63][2] ), 
        .QN(n14508) );
  DFF_X1 \registers_reg[0][2]  ( .D(n7947), .CK(clk), .Q(\registers[0][2] ), 
        .QN(n15797) );
  DFF_X1 \registers_reg[1][2]  ( .D(n7946), .CK(clk), .Q(\registers[1][2] ), 
        .QN(n15581) );
  DFF_X1 \registers_reg[2][2]  ( .D(n7945), .CK(clk), .Q(\registers[2][2] ), 
        .QN(n14775) );
  DFF_X1 \registers_reg[3][2]  ( .D(n7944), .CK(clk), .Q(net226883), .QN(
        n15760) );
  DFF_X1 \registers_reg[8][2]  ( .D(n7943), .CK(clk), .Q(net226882), .QN(
        n15212) );
  DFF_X1 \registers_reg[9][2]  ( .D(n7942), .CK(clk), .Q(\registers[9][2] ), 
        .QN(n14331) );
  DFF_X1 \registers_reg[10][2]  ( .D(n7941), .CK(clk), .Q(\registers[10][2] ), 
        .QN(n14716) );
  DFF_X1 \registers_reg[11][2]  ( .D(n7940), .CK(clk), .Q(\registers[11][2] ), 
        .QN(n14430) );
  DFF_X1 \registers_reg[16][2]  ( .D(n7939), .CK(clk), .Q(\registers[16][2] ), 
        .QN(n15701) );
  DFF_X1 \registers_reg[17][2]  ( .D(n7938), .CK(clk), .Q(\registers[17][2] ), 
        .QN(n14607) );
  DFF_X1 \registers_reg[18][2]  ( .D(n7937), .CK(clk), .Q(\registers[18][2] ), 
        .QN(n14364) );
  DFF_X1 \registers_reg[19][2]  ( .D(n7936), .CK(clk), .Q(\registers[19][2] ), 
        .QN(n15804) );
  DFF_X1 \registers_reg[24][2]  ( .D(n7935), .CK(clk), .Q(net226881), .QN(
        n15183) );
  DFF_X1 \registers_reg[25][2]  ( .D(n7934), .CK(clk), .Q(\registers[25][2] ), 
        .QN(n14302) );
  DFF_X1 \registers_reg[26][2]  ( .D(n7933), .CK(clk), .QN(n12360) );
  DFF_X1 \registers_reg[27][2]  ( .D(n7932), .CK(clk), .QN(n12020) );
  DFF_X1 \registers_reg[32][2]  ( .D(n7931), .CK(clk), .QN(n12311) );
  DFF_X1 \registers_reg[33][2]  ( .D(n7930), .CK(clk), .QN(n11799) );
  DFF_X1 \registers_reg[34][2]  ( .D(n7929), .CK(clk), .Q(\registers[34][2] ), 
        .QN(n15497) );
  DFF_X1 \registers_reg[35][2]  ( .D(n7928), .CK(clk), .Q(net226880), .QN(
        n15586) );
  DFF_X1 \registers_reg[40][2]  ( .D(n7927), .CK(clk), .Q(\registers[40][2] ), 
        .QN(n15077) );
  DFF_X1 \registers_reg[41][2]  ( .D(n7926), .CK(clk), .Q(\registers[41][2] ), 
        .QN(n14431) );
  DFF_X1 \registers_reg[42][2]  ( .D(n7925), .CK(clk), .Q(\registers[42][2] ), 
        .QN(n15922) );
  DFF_X1 \registers_reg[43][2]  ( .D(n7924), .CK(clk), .Q(\registers[43][2] ), 
        .QN(n14890) );
  DFF_X1 \registers_reg[48][2]  ( .D(n7923), .CK(clk), .Q(\registers[48][2] ), 
        .QN(n15554) );
  DFF_X1 \registers_reg[49][2]  ( .D(n7922), .CK(clk), .Q(\registers[49][2] ), 
        .QN(n14486) );
  DFF_X1 \registers_reg[50][2]  ( .D(n7921), .CK(clk), .Q(\registers[50][2] ), 
        .QN(n15971) );
  DFF_X1 \registers_reg[51][2]  ( .D(n7920), .CK(clk), .Q(\registers[51][2] ), 
        .QN(n15401) );
  DFF_X1 \registers_reg[56][2]  ( .D(n7919), .CK(clk), .Q(\registers[56][2] ), 
        .QN(n16000) );
  DFF_X1 \registers_reg[57][2]  ( .D(n7918), .CK(clk), .Q(net226879), .QN(
        n15244) );
  DFF_X1 \registers_reg[58][2]  ( .D(n7917), .CK(clk), .Q(net226878), .QN(
        n14912) );
  DFF_X1 \registers_reg[59][2]  ( .D(n7916), .CK(clk), .Q(\registers[59][2] ), 
        .QN(n15434) );
  DFF_X1 \to_mem_reg[2]  ( .D(n7915), .CK(clk), .QN(n7723) );
  DFF_X1 \registers_reg[64][2]  ( .D(n7914), .CK(clk), .Q(net226877), .QN(
        n16203) );
  DFF_X1 \registers_reg[65][2]  ( .D(n7913), .CK(clk), .Q(net226876), .QN(
        n16113) );
  DFF_X1 \registers_reg[66][2]  ( .D(n7912), .CK(clk), .Q(net226875), .QN(
        n16121) );
  DFF_X1 \registers_reg[67][2]  ( .D(n7911), .CK(clk), .QN(n14286) );
  DFF_X1 \registers_reg[68][2]  ( .D(n7910), .CK(clk), .Q(\registers[68][2] ), 
        .QN(n16207) );
  DFF_X1 \registers_reg[69][2]  ( .D(n7909), .CK(clk), .Q(net226874), .QN(
        n16200) );
  DFF_X1 \registers_reg[70][2]  ( .D(n7908), .CK(clk), .Q(net226873), .QN(
        n16117) );
  DFF_X1 \registers_reg[71][2]  ( .D(n7907), .CK(clk), .QN(n14962) );
  DFF_X1 \out1_reg[2]  ( .D(n7906), .CK(clk), .Q(out1[2]), .QN(net226871) );
  DFF_X1 \registers_reg[2][1]  ( .D(n7905), .CK(clk), .Q(\registers[2][1] ), 
        .QN(n14773) );
  DFF_X1 \registers_reg[3][1]  ( .D(n7904), .CK(clk), .Q(net226870), .QN(
        n15759) );
  DFF_X1 \registers_reg[6][1]  ( .D(n7903), .CK(clk), .QN(n12359) );
  DFF_X1 \registers_reg[7][1]  ( .D(n7902), .CK(clk), .Q(\registers[7][1] ), 
        .QN(n15327) );
  DFF_X1 \registers_reg[10][1]  ( .D(n7901), .CK(clk), .Q(\registers[10][1] ), 
        .QN(n14714) );
  DFF_X1 \registers_reg[11][1]  ( .D(n7900), .CK(clk), .Q(\registers[11][1] ), 
        .QN(n14428) );
  DFF_X1 \registers_reg[14][1]  ( .D(n7899), .CK(clk), .QN(n11882) );
  DFF_X1 \registers_reg[15][1]  ( .D(n7898), .CK(clk), .Q(\registers[15][1] ), 
        .QN(n15293) );
  DFF_X1 \registers_reg[18][1]  ( .D(n7897), .CK(clk), .Q(\registers[18][1] ), 
        .QN(n14360) );
  DFF_X1 \registers_reg[19][1]  ( .D(n7896), .CK(clk), .Q(\registers[19][1] ), 
        .QN(n15793) );
  DFF_X1 \registers_reg[22][1]  ( .D(n7895), .CK(clk), .Q(\registers[22][1] ), 
        .QN(n15371) );
  DFF_X1 \registers_reg[23][1]  ( .D(n7894), .CK(clk), .Q(\registers[23][1] ), 
        .QN(n15882) );
  DFF_X1 \registers_reg[26][1]  ( .D(n7893), .CK(clk), .QN(n12358) );
  DFF_X1 \registers_reg[27][1]  ( .D(n7892), .CK(clk), .QN(n12019) );
  DFF_X1 \registers_reg[30][1]  ( .D(n7891), .CK(clk), .Q(\registers[30][1] ), 
        .QN(n14679) );
  DFF_X1 \registers_reg[31][1]  ( .D(n7890), .CK(clk), .Q(net226869), .QN(
        n15737) );
  DFF_X1 \registers_reg[34][1]  ( .D(n7889), .CK(clk), .Q(\registers[34][1] ), 
        .QN(n15496) );
  DFF_X1 \registers_reg[35][1]  ( .D(n7888), .CK(clk), .Q(net226868), .QN(
        n15577) );
  DFF_X1 \registers_reg[38][1]  ( .D(n7887), .CK(clk), .Q(\registers[38][1] ), 
        .QN(n15035) );
  DFF_X1 \registers_reg[39][1]  ( .D(n7886), .CK(clk), .QN(n12172) );
  DFF_X1 \registers_reg[42][1]  ( .D(n7885), .CK(clk), .Q(\registers[42][1] ), 
        .QN(n15912) );
  DFF_X1 \registers_reg[43][1]  ( .D(n7884), .CK(clk), .Q(\registers[43][1] ), 
        .QN(n14889) );
  DFF_X1 \registers_reg[46][1]  ( .D(n7883), .CK(clk), .QN(n11952) );
  DFF_X1 \registers_reg[47][1]  ( .D(n7882), .CK(clk), .Q(\registers[47][1] ), 
        .QN(n14548) );
  DFF_X1 \registers_reg[50][1]  ( .D(n7881), .CK(clk), .Q(\registers[50][1] ), 
        .QN(n15969) );
  DFF_X1 \registers_reg[51][1]  ( .D(n7880), .CK(clk), .Q(\registers[51][1] ), 
        .QN(n15370) );
  DFF_X1 \registers_reg[54][1]  ( .D(n7879), .CK(clk), .Q(\registers[54][1] ), 
        .QN(n14570) );
  DFF_X1 \registers_reg[55][1]  ( .D(n7878), .CK(clk), .Q(\registers[55][1] ), 
        .QN(n12052) );
  DFF_X1 \registers_reg[58][1]  ( .D(n7877), .CK(clk), .Q(net226866), .QN(
        n14911) );
  DFF_X1 \registers_reg[59][1]  ( .D(n7876), .CK(clk), .Q(\registers[59][1] ), 
        .QN(n15433) );
  DFF_X1 \registers_reg[62][1]  ( .D(n7875), .CK(clk), .Q(\registers[62][1] ), 
        .QN(n15124) );
  DFF_X1 \registers_reg[63][1]  ( .D(n7874), .CK(clk), .Q(\registers[63][1] ), 
        .QN(n14507) );
  DFF_X1 \registers_reg[66][1]  ( .D(n7873), .CK(clk), .Q(net226865), .QN(
        n16116) );
  DFF_X1 \registers_reg[67][1]  ( .D(n7872), .CK(clk), .QN(n14285) );
  DFF_X1 \registers_reg[0][1]  ( .D(n7871), .CK(clk), .Q(\registers[0][1] ), 
        .QN(n15796) );
  DFF_X1 \registers_reg[1][1]  ( .D(n7870), .CK(clk), .Q(\registers[1][1] ), 
        .QN(n15580) );
  DFF_X1 \registers_reg[4][1]  ( .D(n7869), .CK(clk), .Q(\registers[4][1] ), 
        .QN(n15522) );
  DFF_X1 \registers_reg[5][1]  ( .D(n7868), .CK(clk), .Q(\registers[5][1] ), 
        .QN(n14713) );
  DFF_X1 \registers_reg[8][1]  ( .D(n7867), .CK(clk), .Q(net226864), .QN(
        n15211) );
  DFF_X1 \registers_reg[9][1]  ( .D(n7866), .CK(clk), .Q(\registers[9][1] ), 
        .QN(n14330) );
  DFF_X1 \registers_reg[12][1]  ( .D(n7865), .CK(clk), .Q(\registers[12][1] ), 
        .QN(n15670) );
  DFF_X1 \registers_reg[13][1]  ( .D(n7864), .CK(clk), .Q(net226863), .QN(
        n15074) );
  DFF_X1 \registers_reg[16][1]  ( .D(n7863), .CK(clk), .Q(\registers[16][1] ), 
        .QN(n15700) );
  DFF_X1 \registers_reg[17][1]  ( .D(n7862), .CK(clk), .Q(\registers[17][1] ), 
        .QN(n14606) );
  DFF_X1 \registers_reg[20][1]  ( .D(n7861), .CK(clk), .QN(n14832) );
  DFF_X1 \registers_reg[21][1]  ( .D(n7860), .CK(clk), .QN(n12206) );
  DFF_X1 \registers_reg[24][1]  ( .D(n7859), .CK(clk), .Q(net226862), .QN(
        n15182) );
  DFF_X1 \registers_reg[25][1]  ( .D(n7858), .CK(clk), .Q(\registers[25][1] ), 
        .QN(n14301) );
  DFF_X1 \registers_reg[28][1]  ( .D(n7857), .CK(clk), .Q(net226861), .QN(
        n15005) );
  DFF_X1 \registers_reg[29][1]  ( .D(n7856), .CK(clk), .Q(\registers[29][1] ), 
        .QN(n15803) );
  DFF_X1 \registers_reg[32][1]  ( .D(n7855), .CK(clk), .QN(n12310) );
  DFF_X1 \registers_reg[33][1]  ( .D(n7854), .CK(clk), .QN(n11756) );
  DFF_X1 \registers_reg[36][1]  ( .D(n7853), .CK(clk), .Q(\registers[36][1] ), 
        .QN(n15153) );
  DFF_X1 \registers_reg[37][1]  ( .D(n7852), .CK(clk), .Q(\registers[37][1] ), 
        .QN(n14363) );
  DFF_X1 \registers_reg[40][1]  ( .D(n7851), .CK(clk), .Q(\registers[40][1] ), 
        .QN(n15075) );
  DFF_X1 \registers_reg[41][1]  ( .D(n7850), .CK(clk), .Q(\registers[41][1] ), 
        .QN(n14429) );
  DFF_X1 \registers_reg[44][1]  ( .D(n7849), .CK(clk), .Q(\registers[44][1] ), 
        .QN(n15467) );
  DFF_X1 \registers_reg[45][1]  ( .D(n7848), .CK(clk), .Q(\registers[45][1] ), 
        .QN(n14774) );
  DFF_X1 \registers_reg[48][1]  ( .D(n7847), .CK(clk), .Q(\registers[48][1] ), 
        .QN(n15553) );
  DFF_X1 \registers_reg[49][1]  ( .D(n7846), .CK(clk), .Q(\registers[49][1] ), 
        .QN(n14485) );
  DFF_X1 \registers_reg[52][1]  ( .D(n7845), .CK(clk), .Q(net226860), .QN(
        n14939) );
  DFF_X1 \registers_reg[53][1]  ( .D(n7844), .CK(clk), .Q(net226859), .QN(
        n15914) );
  DFF_X1 \registers_reg[56][1]  ( .D(n7843), .CK(clk), .Q(\registers[56][1] ), 
        .QN(n15999) );
  DFF_X1 \registers_reg[57][1]  ( .D(n7842), .CK(clk), .Q(net226858), .QN(
        n15243) );
  DFF_X1 \registers_reg[60][1]  ( .D(n7841), .CK(clk), .Q(\registers[60][1] ), 
        .QN(n14645) );
  DFF_X1 \registers_reg[61][1]  ( .D(n7840), .CK(clk), .Q(net226857), .QN(
        n15661) );
  DFF_X1 \to_mem_reg[1]  ( .D(n7839), .CK(clk), .QN(n7724) );
  DFF_X1 \registers_reg[64][1]  ( .D(n7838), .CK(clk), .Q(net226856), .QN(
        n16202) );
  DFF_X1 \registers_reg[65][1]  ( .D(n7837), .CK(clk), .Q(net226855), .QN(
        n16112) );
  DFF_X1 \registers_reg[68][1]  ( .D(n7836), .CK(clk), .Q(\registers[68][1] ), 
        .QN(n16209) );
  DFF_X1 \registers_reg[69][1]  ( .D(n7835), .CK(clk), .Q(net226854), .QN(
        n16205) );
  DFF_X1 \registers_reg[70][1]  ( .D(n7834), .CK(clk), .Q(net226853), .QN(
        n16115) );
  DFF_X1 \registers_reg[71][1]  ( .D(n7833), .CK(clk), .QN(n14961) );
  DFF_X1 \out1_reg[1]  ( .D(n7832), .CK(clk), .Q(out1[1]), .QN(net226851) );
  DFF_X1 \registers_reg[1][0]  ( .D(n7831), .CK(clk), .Q(\registers[1][0] ), 
        .QN(n15576) );
  DFF_X1 \registers_reg[3][0]  ( .D(n7830), .CK(clk), .Q(net226850), .QN(
        n15758) );
  DFF_X1 \registers_reg[5][0]  ( .D(n7829), .CK(clk), .Q(\registers[5][0] ), 
        .QN(n14711) );
  DFF_X1 \registers_reg[7][0]  ( .D(n7828), .CK(clk), .Q(\registers[7][0] ), 
        .QN(n15326) );
  DFF_X1 \registers_reg[9][0]  ( .D(n7827), .CK(clk), .Q(\registers[9][0] ), 
        .QN(n14329) );
  DFF_X1 \registers_reg[11][0]  ( .D(n7826), .CK(clk), .Q(\registers[11][0] ), 
        .QN(n14426) );
  DFF_X1 \registers_reg[13][0]  ( .D(n7825), .CK(clk), .Q(net226849), .QN(
        n15072) );
  DFF_X1 \registers_reg[15][0]  ( .D(n7824), .CK(clk), .Q(\registers[15][0] ), 
        .QN(n15292) );
  DFF_X1 \registers_reg[17][0]  ( .D(n7823), .CK(clk), .Q(\registers[17][0] ), 
        .QN(n14605) );
  DFF_X1 \registers_reg[19][0]  ( .D(n7822), .CK(clk), .Q(\registers[19][0] ), 
        .QN(n15792) );
  DFF_X1 \registers_reg[21][0]  ( .D(n7821), .CK(clk), .QN(n12205) );
  DFF_X1 \registers_reg[23][0]  ( .D(n7820), .CK(clk), .Q(\registers[23][0] ), 
        .QN(n15881) );
  DFF_X1 \registers_reg[25][0]  ( .D(n7819), .CK(clk), .Q(\registers[25][0] ), 
        .QN(n14300) );
  DFF_X1 \registers_reg[27][0]  ( .D(n7818), .CK(clk), .QN(n12018) );
  DFF_X1 \registers_reg[29][0]  ( .D(n7817), .CK(clk), .Q(\registers[29][0] ), 
        .QN(n15791) );
  DFF_X1 \registers_reg[31][0]  ( .D(n7816), .CK(clk), .Q(net226848), .QN(
        n15736) );
  DFF_X1 \registers_reg[33][0]  ( .D(n7815), .CK(clk), .QN(n11713) );
  DFF_X1 \registers_reg[35][0]  ( .D(n7814), .CK(clk), .Q(net226847), .QN(
        n15575) );
  DFF_X1 \registers_reg[37][0]  ( .D(n7813), .CK(clk), .Q(\registers[37][0] ), 
        .QN(n14359) );
  DFF_X1 \registers_reg[39][0]  ( .D(n7812), .CK(clk), .QN(n12171) );
  DFF_X1 \registers_reg[41][0]  ( .D(n7811), .CK(clk), .Q(\registers[41][0] ), 
        .QN(n14427) );
  DFF_X1 \registers_reg[43][0]  ( .D(n7810), .CK(clk), .Q(\registers[43][0] ), 
        .QN(n14888) );
  DFF_X1 \registers_reg[45][0]  ( .D(n7809), .CK(clk), .Q(\registers[45][0] ), 
        .QN(n14772) );
  DFF_X1 \registers_reg[47][0]  ( .D(n7808), .CK(clk), .Q(\registers[47][0] ), 
        .QN(n14547) );
  DFF_X1 \registers_reg[49][0]  ( .D(n7807), .CK(clk), .Q(\registers[49][0] ), 
        .QN(n14484) );
  DFF_X1 \registers_reg[51][0]  ( .D(n7806), .CK(clk), .Q(\registers[51][0] ), 
        .QN(n15369) );
  DFF_X1 \registers_reg[53][0]  ( .D(n7805), .CK(clk), .Q(net226846), .QN(
        n15911) );
  DFF_X1 \registers_reg[55][0]  ( .D(n7804), .CK(clk), .Q(\registers[55][0] ), 
        .QN(n12055) );
  DFF_X1 \registers_reg[57][0]  ( .D(n7803), .CK(clk), .Q(net226845), .QN(
        n15245) );
  DFF_X1 \registers_reg[59][0]  ( .D(n7802), .CK(clk), .Q(\registers[59][0] ), 
        .QN(n15432) );
  DFF_X1 \registers_reg[61][0]  ( .D(n7801), .CK(clk), .Q(net226844), .QN(
        n15574) );
  DFF_X1 \registers_reg[63][0]  ( .D(n7800), .CK(clk), .Q(\registers[63][0] ), 
        .QN(n14506) );
  DFF_X1 \registers_reg[65][0]  ( .D(n7799), .CK(clk), .Q(net226843), .QN(
        n16111) );
  DFF_X1 \registers_reg[67][0]  ( .D(n7798), .CK(clk), .QN(n14284) );
  DFF_X1 \registers_reg[69][0]  ( .D(n7797), .CK(clk), .Q(net226842), .QN(
        n16199) );
  DFF_X1 \registers_reg[0][0]  ( .D(n7796), .CK(clk), .Q(\registers[0][0] ), 
        .QN(n15795) );
  DFF_X1 \registers_reg[2][0]  ( .D(n7795), .CK(clk), .Q(\registers[2][0] ), 
        .QN(n14771) );
  DFF_X1 \registers_reg[4][0]  ( .D(n7794), .CK(clk), .Q(\registers[4][0] ), 
        .QN(n15521) );
  DFF_X1 \registers_reg[6][0]  ( .D(n7793), .CK(clk), .QN(n12357) );
  DFF_X1 \registers_reg[8][0]  ( .D(n7792), .CK(clk), .Q(net226841), .QN(
        n15210) );
  DFF_X1 \registers_reg[10][0]  ( .D(n7791), .CK(clk), .Q(\registers[10][0] ), 
        .QN(n14712) );
  DFF_X1 \registers_reg[12][0]  ( .D(n7790), .CK(clk), .Q(\registers[12][0] ), 
        .QN(n15669) );
  DFF_X1 \registers_reg[14][0]  ( .D(n7789), .CK(clk), .QN(n11881) );
  DFF_X1 \registers_reg[16][0]  ( .D(n7788), .CK(clk), .Q(\registers[16][0] ), 
        .QN(n15699) );
  DFF_X1 \registers_reg[18][0]  ( .D(n7787), .CK(clk), .Q(\registers[18][0] ), 
        .QN(n14362) );
  DFF_X1 \registers_reg[20][0]  ( .D(n7786), .CK(clk), .QN(n14831) );
  DFF_X1 \registers_reg[22][0]  ( .D(n7785), .CK(clk), .Q(\registers[22][0] ), 
        .QN(n15373) );
  DFF_X1 \registers_reg[24][0]  ( .D(n7784), .CK(clk), .Q(net226840), .QN(
        n15181) );
  DFF_X1 \registers_reg[26][0]  ( .D(n7783), .CK(clk), .QN(n12356) );
  DFF_X1 \registers_reg[28][0]  ( .D(n7782), .CK(clk), .Q(net226839), .QN(
        n15004) );
  DFF_X1 \registers_reg[30][0]  ( .D(n7781), .CK(clk), .Q(\registers[30][0] ), 
        .QN(n14678) );
  DFF_X1 \registers_reg[32][0]  ( .D(n7780), .CK(clk), .QN(n12309) );
  DFF_X1 \registers_reg[34][0]  ( .D(n7779), .CK(clk), .Q(\registers[34][0] ), 
        .QN(n15495) );
  DFF_X1 \registers_reg[36][0]  ( .D(n7778), .CK(clk), .Q(\registers[36][0] ), 
        .QN(n15152) );
  DFF_X1 \registers_reg[38][0]  ( .D(n7777), .CK(clk), .Q(\registers[38][0] ), 
        .QN(n15037) );
  DFF_X1 \registers_reg[40][0]  ( .D(n7776), .CK(clk), .Q(\registers[40][0] ), 
        .QN(n15073) );
  DFF_X1 \registers_reg[42][0]  ( .D(n7775), .CK(clk), .Q(\registers[42][0] ), 
        .QN(n15921) );
  DFF_X1 \registers_reg[44][0]  ( .D(n7774), .CK(clk), .Q(\registers[44][0] ), 
        .QN(n15466) );
  DFF_X1 \registers_reg[46][0]  ( .D(n7773), .CK(clk), .QN(n11951) );
  DFF_X1 \registers_reg[48][0]  ( .D(n7772), .CK(clk), .Q(\registers[48][0] ), 
        .QN(n15552) );
  DFF_X1 \registers_reg[50][0]  ( .D(n7771), .CK(clk), .Q(\registers[50][0] ), 
        .QN(n15970) );
  DFF_X1 \registers_reg[52][0]  ( .D(n7770), .CK(clk), .Q(net226837), .QN(
        n14938) );
  DFF_X1 \registers_reg[54][0]  ( .D(n7769), .CK(clk), .Q(\registers[54][0] ), 
        .QN(n14573) );
  DFF_X1 \registers_reg[56][0]  ( .D(n7768), .CK(clk), .Q(\registers[56][0] ), 
        .QN(n15998) );
  DFF_X1 \registers_reg[58][0]  ( .D(n7767), .CK(clk), .Q(net226836), .QN(
        n14910) );
  DFF_X1 \registers_reg[60][0]  ( .D(n7766), .CK(clk), .Q(\registers[60][0] ), 
        .QN(n14669) );
  DFF_X1 \registers_reg[62][0]  ( .D(n7765), .CK(clk), .Q(\registers[62][0] ), 
        .QN(n15123) );
  DFF_X1 \to_mem_reg[0]  ( .D(n7764), .CK(clk), .QN(n7725) );
  DFF_X1 \registers_reg[64][0]  ( .D(n7763), .CK(clk), .Q(net226835), .QN(
        n16201) );
  DFF_X1 \registers_reg[66][0]  ( .D(n7762), .CK(clk), .Q(net226834), .QN(
        n16120) );
  DFF_X1 \registers_reg[68][0]  ( .D(n7761), .CK(clk), .Q(\registers[68][0] ), 
        .QN(n16208) );
  DFF_X1 \registers_reg[70][0]  ( .D(n7760), .CK(clk), .Q(net226833), .QN(
        n16118) );
  DFF_X1 \registers_reg[71][0]  ( .D(n7759), .CK(clk), .QN(n14960) );
  DFF_X1 \out1_reg[0]  ( .D(n7758), .CK(clk), .Q(out1[0]), .QN(net226831) );
  DFF_X1 \out2_reg[31]  ( .D(n7757), .CK(clk), .Q(out2[31]), .QN(net226830) );
  DFF_X1 \out2_reg[30]  ( .D(n7756), .CK(clk), .Q(out2[30]), .QN(net226829) );
  DFF_X1 \out2_reg[29]  ( .D(n7755), .CK(clk), .Q(out2[29]), .QN(net226828) );
  DFF_X1 \out2_reg[28]  ( .D(n7754), .CK(clk), .Q(out2[28]), .QN(net226827) );
  DFF_X1 \out2_reg[27]  ( .D(n7753), .CK(clk), .Q(out2[27]), .QN(net226826) );
  DFF_X1 \out2_reg[26]  ( .D(n7752), .CK(clk), .Q(out2[26]), .QN(net226825) );
  DFF_X1 \out2_reg[25]  ( .D(n7751), .CK(clk), .Q(out2[25]), .QN(net226824) );
  DFF_X1 \out2_reg[24]  ( .D(n7750), .CK(clk), .Q(out2[24]), .QN(net226823) );
  DFF_X1 \out2_reg[23]  ( .D(n7749), .CK(clk), .Q(out2[23]), .QN(net226822) );
  DFF_X1 \out2_reg[22]  ( .D(n7748), .CK(clk), .Q(out2[22]), .QN(net226821) );
  DFF_X1 \out2_reg[21]  ( .D(n7747), .CK(clk), .Q(out2[21]), .QN(net226820) );
  DFF_X1 \out2_reg[20]  ( .D(n7746), .CK(clk), .Q(out2[20]), .QN(net226819) );
  DFF_X1 \out2_reg[19]  ( .D(n7745), .CK(clk), .Q(out2[19]), .QN(net226818) );
  DFF_X1 \out2_reg[18]  ( .D(n7744), .CK(clk), .Q(out2[18]), .QN(net226817) );
  DFF_X1 \out2_reg[17]  ( .D(n7743), .CK(clk), .Q(out2[17]), .QN(net226816) );
  DFF_X1 \out2_reg[16]  ( .D(n7742), .CK(clk), .Q(out2[16]), .QN(net226815) );
  DFF_X1 \out2_reg[15]  ( .D(n7741), .CK(clk), .Q(out2[15]), .QN(net226814) );
  DFF_X1 \out2_reg[14]  ( .D(n7740), .CK(clk), .Q(out2[14]), .QN(net226813) );
  DFF_X1 \out2_reg[13]  ( .D(n7739), .CK(clk), .Q(out2[13]), .QN(net226812) );
  DFF_X1 \out2_reg[12]  ( .D(n7738), .CK(clk), .Q(out2[12]), .QN(net226811) );
  DFF_X1 \out2_reg[11]  ( .D(n7737), .CK(clk), .Q(out2[11]), .QN(net226810) );
  DFF_X1 \out2_reg[10]  ( .D(n7736), .CK(clk), .Q(out2[10]), .QN(net226809) );
  DFF_X1 \out2_reg[9]  ( .D(n7735), .CK(clk), .Q(out2[9]), .QN(net226808) );
  DFF_X1 \out2_reg[8]  ( .D(n7734), .CK(clk), .Q(out2[8]), .QN(net226807) );
  DFF_X1 \out2_reg[7]  ( .D(n7733), .CK(clk), .Q(out2[7]), .QN(net226806) );
  DFF_X1 \out2_reg[6]  ( .D(n7732), .CK(clk), .Q(out2[6]), .QN(net226805) );
  DFF_X1 \out2_reg[5]  ( .D(n7731), .CK(clk), .Q(out2[5]), .QN(net226804) );
  DFF_X1 \out2_reg[4]  ( .D(n7730), .CK(clk), .Q(out2[4]), .QN(net226803) );
  DFF_X1 \out2_reg[3]  ( .D(n7729), .CK(clk), .Q(out2[3]), .QN(net226802) );
  DFF_X1 \out2_reg[2]  ( .D(n7728), .CK(clk), .Q(out2[2]), .QN(net226801) );
  DFF_X1 \out2_reg[1]  ( .D(n7727), .CK(clk), .Q(out2[1]), .QN(net226800) );
  DFF_X1 \out2_reg[0]  ( .D(n7726), .CK(clk), .Q(out2[0]), .QN(net226799) );
  FA_X1 \add_73/U1_1  ( .A(N191), .B(\lastcwp[1] ), .CI(\add_73/carry[1] ), 
        .CO(\add_73/carry[2] ), .S(N273) );
  FA_X1 \add_73/U1_2  ( .A(N192), .B(\lastcwp[2] ), .CI(\add_73/carry[2] ), 
        .CO(\add_73/carry[3] ), .S(N274) );
  FA_X1 \add_73/U1_3  ( .A(\sub_71/carry[4] ), .B(\lastcwp[3] ), .CI(
        \add_73/carry[3] ), .CO(\add_73/carry[4] ), .S(N275) );
  FA_X1 \add_73/U1_4  ( .A(add_wr[4]), .B(\lastcwp[4] ), .CI(\add_73/carry[4] ), .CO(\add_73/carry[5] ), .S(N276) );
  DFF_X1 \cwp_reg[3]  ( .D(n10175), .CK(clk), .Q(N9910), .QN(n10187) );
  DFF_X1 \cwp_reg[2]  ( .D(n10177), .CK(clk), .Q(N9909), .QN(n10188) );
  DFF_X1 \cwp_reg[1]  ( .D(n10179), .CK(clk), .Q(N9908), .QN(n10189) );
  DFF_X1 \cwp_reg[0]  ( .D(n10180), .CK(clk), .Q(N9641), .QN(n10190) );
  NOR4_X2 U8886 ( .A1(n14173), .A2(N9924), .A3(N9926), .A4(call), .ZN(n14105)
         );
  NOR4_X2 U8949 ( .A1(N9922), .A2(N9924), .A3(N9926), .A4(call), .ZN(n14095)
         );
  NAND3_X1 U9269 ( .A1(n10513), .A2(n10514), .A3(n10515), .ZN(n8108) );
  NAND3_X1 U9270 ( .A1(n10665), .A2(n10666), .A3(n10667), .ZN(n8106) );
  NAND3_X1 U9271 ( .A1(n10724), .A2(n10725), .A3(n10726), .ZN(n8104) );
  NAND3_X1 U9272 ( .A1(n10767), .A2(n10768), .A3(n10769), .ZN(n8102) );
  NAND3_X1 U9273 ( .A1(n10810), .A2(n10811), .A3(n10812), .ZN(n8100) );
  NAND3_X1 U9274 ( .A1(n10853), .A2(n10854), .A3(n10855), .ZN(n8098) );
  NAND3_X1 U9275 ( .A1(n10896), .A2(n10897), .A3(n10898), .ZN(n8096) );
  NAND3_X1 U9276 ( .A1(n10939), .A2(n10940), .A3(n10941), .ZN(n8094) );
  NAND3_X1 U9277 ( .A1(n10982), .A2(n10983), .A3(n10984), .ZN(n8092) );
  NAND3_X1 U9278 ( .A1(n11025), .A2(n11026), .A3(n11027), .ZN(n8090) );
  NAND3_X1 U9279 ( .A1(n11068), .A2(n11069), .A3(n11070), .ZN(n8088) );
  NAND3_X1 U9280 ( .A1(n11111), .A2(n11112), .A3(n11113), .ZN(n8086) );
  NAND3_X1 U9281 ( .A1(n11154), .A2(n11155), .A3(n11156), .ZN(n8084) );
  NAND3_X1 U9282 ( .A1(n11197), .A2(n11198), .A3(n11199), .ZN(n8082) );
  NAND3_X1 U9283 ( .A1(n11240), .A2(n11241), .A3(n11242), .ZN(n8080) );
  NAND3_X1 U9284 ( .A1(n11283), .A2(n11284), .A3(n11285), .ZN(n8078) );
  NAND3_X1 U9285 ( .A1(n11326), .A2(n11327), .A3(n11328), .ZN(n8076) );
  NAND3_X1 U9286 ( .A1(n11369), .A2(n11370), .A3(n11371), .ZN(n8074) );
  NAND3_X1 U9287 ( .A1(n11412), .A2(n11413), .A3(n11414), .ZN(n8072) );
  NAND3_X1 U9288 ( .A1(n11455), .A2(n11456), .A3(n11457), .ZN(n8070) );
  NAND3_X1 U9289 ( .A1(n11499), .A2(n11500), .A3(n11501), .ZN(n8068) );
  NAND3_X1 U9290 ( .A1(n11542), .A2(n11543), .A3(n11544), .ZN(n8066) );
  NAND3_X1 U9291 ( .A1(n11585), .A2(n11586), .A3(n11587), .ZN(n8064) );
  NAND3_X1 U9292 ( .A1(n11628), .A2(n11629), .A3(n11630), .ZN(n8062) );
  NAND3_X1 U9293 ( .A1(n11671), .A2(n11672), .A3(n11673), .ZN(n8060) );
  NAND3_X1 U9294 ( .A1(n11714), .A2(n11715), .A3(n11716), .ZN(n8058) );
  NAND3_X1 U9295 ( .A1(n11757), .A2(n11758), .A3(n11759), .ZN(n8056) );
  NAND3_X1 U9296 ( .A1(n11800), .A2(n11801), .A3(n11802), .ZN(n8054) );
  NAND3_X1 U9297 ( .A1(n11953), .A2(n11954), .A3(n11955), .ZN(n7980) );
  NAND3_X1 U9298 ( .A1(n12106), .A2(n12107), .A3(n12108), .ZN(n7906) );
  NAND3_X1 U9299 ( .A1(n12259), .A2(n12260), .A3(n12261), .ZN(n7832) );
  NAND3_X1 U9300 ( .A1(n12416), .A2(n12417), .A3(n12418), .ZN(n7758) );
  XOR2_X1 U9301 ( .A(\sub_71/carry[4] ), .B(\sub_132/carry[4] ), .Z(n12515) );
  NAND3_X1 U9302 ( .A1(enable), .A2(n18044), .A3(rd1), .ZN(n10525) );
  NAND3_X1 U9303 ( .A1(n12516), .A2(n12517), .A3(n12518), .ZN(n7757) );
  NAND3_X1 U9304 ( .A1(n12635), .A2(n12636), .A3(n12637), .ZN(n7756) );
  NAND3_X1 U9305 ( .A1(n12679), .A2(n12680), .A3(n12681), .ZN(n7755) );
  NAND3_X1 U9306 ( .A1(n12721), .A2(n12722), .A3(n12723), .ZN(n7754) );
  NAND3_X1 U9307 ( .A1(n12763), .A2(n12764), .A3(n12765), .ZN(n7753) );
  NAND3_X1 U9308 ( .A1(n12805), .A2(n12806), .A3(n12807), .ZN(n7752) );
  NAND3_X1 U9309 ( .A1(n12847), .A2(n12848), .A3(n12849), .ZN(n7751) );
  NAND3_X1 U9310 ( .A1(n12889), .A2(n12890), .A3(n12891), .ZN(n7750) );
  NAND3_X1 U9311 ( .A1(n12931), .A2(n12932), .A3(n12933), .ZN(n7749) );
  NAND3_X1 U9312 ( .A1(n12973), .A2(n12974), .A3(n12975), .ZN(n7748) );
  NAND3_X1 U9313 ( .A1(n13015), .A2(n13016), .A3(n13017), .ZN(n7747) );
  NAND3_X1 U9314 ( .A1(n13057), .A2(n13058), .A3(n13059), .ZN(n7746) );
  NAND3_X1 U9315 ( .A1(n13099), .A2(n13100), .A3(n13101), .ZN(n7745) );
  NAND3_X1 U9316 ( .A1(n13141), .A2(n13142), .A3(n13143), .ZN(n7744) );
  NAND3_X1 U9317 ( .A1(n13183), .A2(n13184), .A3(n13185), .ZN(n7743) );
  NAND3_X1 U9318 ( .A1(n13225), .A2(n13226), .A3(n13227), .ZN(n7742) );
  NAND3_X1 U9319 ( .A1(n13267), .A2(n13268), .A3(n13269), .ZN(n7741) );
  NAND3_X1 U9320 ( .A1(n13309), .A2(n13310), .A3(n13311), .ZN(n7740) );
  NAND3_X1 U9321 ( .A1(n13351), .A2(n13352), .A3(n13353), .ZN(n7739) );
  NAND3_X1 U9322 ( .A1(n13393), .A2(n13394), .A3(n13395), .ZN(n7738) );
  NAND3_X1 U9323 ( .A1(n13435), .A2(n13436), .A3(n13437), .ZN(n7737) );
  NAND3_X1 U9324 ( .A1(n13477), .A2(n13478), .A3(n13479), .ZN(n7736) );
  NAND3_X1 U9325 ( .A1(n13519), .A2(n13520), .A3(n13521), .ZN(n7735) );
  NAND3_X1 U9326 ( .A1(n13561), .A2(n13562), .A3(n13563), .ZN(n7734) );
  NAND3_X1 U9327 ( .A1(n13603), .A2(n13604), .A3(n13605), .ZN(n7733) );
  NAND3_X1 U9328 ( .A1(n13645), .A2(n13646), .A3(n13647), .ZN(n7732) );
  NAND3_X1 U9329 ( .A1(n13687), .A2(n13688), .A3(n13689), .ZN(n7731) );
  NAND3_X1 U9330 ( .A1(n13729), .A2(n13730), .A3(n13731), .ZN(n7730) );
  NAND3_X1 U9331 ( .A1(n13771), .A2(n13772), .A3(n13773), .ZN(n7729) );
  NAND3_X1 U9332 ( .A1(n13813), .A2(n13814), .A3(n13815), .ZN(n7728) );
  NAND3_X1 U9333 ( .A1(n13855), .A2(n13856), .A3(n13857), .ZN(n7727) );
  NAND3_X1 U9334 ( .A1(n13897), .A2(n13898), .A3(n13899), .ZN(n7726) );
  XOR2_X1 U9335 ( .A(\sub_71/carry[4] ), .B(\sub_146/carry[4] ), .Z(n13995) );
  NAND3_X1 U9336 ( .A1(enable), .A2(n18044), .A3(rd2), .ZN(n12527) );
  XOR2_X1 U9337 ( .A(n3043), .B(n14011), .Z(n14010) );
  NAND3_X1 U9338 ( .A1(call), .A2(n14023), .A3(n14024), .ZN(n13997) );
  NAND3_X1 U9339 ( .A1(n14025), .A2(n14024), .A3(ret), .ZN(n13998) );
  XOR2_X1 U9340 ( .A(swp[5]), .B(n3043), .Z(n14023) );
  NAND3_X1 U9341 ( .A1(n14129), .A2(\r590/carry[5] ), .A3(n14147), .ZN(n14101)
         );
  NAND3_X1 U9342 ( .A1(\r590/carry[5] ), .A2(n14133), .A3(n14147), .ZN(n14142)
         );
  NAND3_X1 U9343 ( .A1(N9926), .A2(N9924), .A3(N9922), .ZN(n14183) );
  NAND3_X1 U9344 ( .A1(\r590/carry[5] ), .A2(n14133), .A3(n14178), .ZN(n14185)
         );
  NAND3_X1 U9345 ( .A1(N9924), .A2(n14173), .A3(N9926), .ZN(n14207) );
  NAND3_X1 U9346 ( .A1(n14178), .A2(\r590/carry[5] ), .A3(n14129), .ZN(n14181)
         );
  NAND3_X1 U9347 ( .A1(n14193), .A2(call), .A3(n14179), .ZN(n14211) );
  NAND3_X1 U9348 ( .A1(n14196), .A2(n10189), .A3(n10187), .ZN(n14116) );
  XOR2_X1 U9349 ( .A(n3043), .B(n14820), .Z(n14178) );
  XOR2_X1 U9353 ( .A(n7587), .B(n14229), .Z(n14263) );
  w_reg_file_M8_N8_F4_Nbit32_DW01_add_0 add_148 ( .A({1'b0, add_rd2[4], 
        \sub_146/carry[4] , N46058, N46057, N46056}), .B({N51637, 
        \r590/carry[5] , N9910, N9909, N9908, N9641}), .CI(1'b0), .SUM({N46303, 
        N46302, N46301, N46300, N46299, N46298}) );
  w_reg_file_M8_N8_F4_Nbit32_DW01_add_1 add_134 ( .A({1'b0, add_rd1[4], 
        \sub_132/carry[4] , N45544, N45543, N45542}), .B({N51637, 
        \r590/carry[5] , N9910, N9909, N9908, N9641}), .CI(1'b0), .SUM({N45789, 
        N45788, N45787, N45786, N45785, N45784}) );
  w_reg_file_M8_N8_F4_Nbit32_DW01_inc_0 add_101 ( .A(i[5:0]), .SUM({N9926, 
        N9925, N9924, N9923, N9922, N9921}) );
  DFF_X1 \cwp_reg[4]  ( .D(n10182), .CK(clk), .Q(\r590/carry[5] ), .QN(n14820)
         );
  NOR2_X1 U6 ( .A1(n13979), .A2(N46298), .ZN(n13932) );
  NOR2_X1 U7 ( .A1(n12498), .A2(N45784), .ZN(n12452) );
  TINV_X1 U8 ( .I(n7694), .EN(n6613), .ZN(to_mem[31]) );
  TINV_X1 U9 ( .I(n7695), .EN(n6620), .ZN(to_mem[30]) );
  TINV_X1 U10 ( .I(n7696), .EN(n6621), .ZN(to_mem[29]) );
  TINV_X1 U11 ( .I(n7697), .EN(n6624), .ZN(to_mem[28]) );
  TINV_X1 U12 ( .I(n7698), .EN(n6630), .ZN(to_mem[27]) );
  TINV_X1 U13 ( .I(n7699), .EN(n6632), .ZN(to_mem[26]) );
  TINV_X1 U14 ( .I(n7700), .EN(n6634), .ZN(to_mem[25]) );
  TINV_X1 U15 ( .I(n7701), .EN(n6641), .ZN(to_mem[24]) );
  TINV_X1 U16 ( .I(n7702), .EN(n6642), .ZN(to_mem[23]) );
  TINV_X1 U17 ( .I(n7703), .EN(n6646), .ZN(to_mem[22]) );
  TINV_X1 U18 ( .I(n7704), .EN(n6647), .ZN(to_mem[21]) );
  TINV_X1 U19 ( .I(n7705), .EN(n6648), .ZN(to_mem[20]) );
  TINV_X1 U20 ( .I(n7706), .EN(n6649), .ZN(to_mem[19]) );
  TINV_X1 U21 ( .I(n7707), .EN(n6650), .ZN(to_mem[18]) );
  TINV_X1 U22 ( .I(n7708), .EN(n6651), .ZN(to_mem[17]) );
  TINV_X1 U23 ( .I(n7709), .EN(n6652), .ZN(to_mem[16]) );
  TINV_X1 U24 ( .I(n7710), .EN(n6653), .ZN(to_mem[15]) );
  TINV_X1 U25 ( .I(n7711), .EN(n6654), .ZN(to_mem[14]) );
  TINV_X1 U26 ( .I(n7712), .EN(n6655), .ZN(to_mem[13]) );
  TINV_X1 U27 ( .I(n7713), .EN(n6656), .ZN(to_mem[12]) );
  TINV_X1 U28 ( .I(n7714), .EN(n6657), .ZN(to_mem[11]) );
  TINV_X1 U29 ( .I(n7715), .EN(n6658), .ZN(to_mem[10]) );
  TINV_X1 U30 ( .I(n7716), .EN(n6659), .ZN(to_mem[9]) );
  TINV_X1 U31 ( .I(n7717), .EN(n6660), .ZN(to_mem[8]) );
  TINV_X1 U32 ( .I(n7718), .EN(n6671), .ZN(to_mem[7]) );
  TINV_X1 U33 ( .I(n7719), .EN(n6674), .ZN(to_mem[6]) );
  TINV_X1 U34 ( .I(n7720), .EN(n6676), .ZN(to_mem[5]) );
  TINV_X1 U35 ( .I(n7721), .EN(n6683), .ZN(to_mem[4]) );
  TINV_X1 U36 ( .I(n7722), .EN(n6684), .ZN(to_mem[3]) );
  TINV_X1 U37 ( .I(n7723), .EN(n6687), .ZN(to_mem[2]) );
  TINV_X1 U38 ( .I(n7724), .EN(n6693), .ZN(to_mem[1]) );
  TINV_X1 U39 ( .I(n7725), .EN(n6695), .ZN(to_mem[0]) );
  NOR2_X1 U40 ( .A1(n13979), .A2(n13978), .ZN(n13918) );
  NOR2_X1 U41 ( .A1(n12498), .A2(n12497), .ZN(n12437) );
  NOR2_X1 U42 ( .A1(N45784), .A2(N45785), .ZN(n12451) );
  NOR2_X1 U43 ( .A1(N46298), .A2(N46299), .ZN(n13927) );
  NOR2_X1 U44 ( .A1(n13978), .A2(N46299), .ZN(n13935) );
  NOR2_X1 U45 ( .A1(n12497), .A2(N45785), .ZN(n12454) );
  INV_X1 U46 ( .A(n17984), .ZN(n17965) );
  INV_X1 U47 ( .A(n17324), .ZN(n17321) );
  INV_X1 U48 ( .A(n17337), .ZN(n17334) );
  INV_X1 U49 ( .A(n17350), .ZN(n17347) );
  INV_X1 U50 ( .A(n17363), .ZN(n17360) );
  INV_X1 U51 ( .A(n17402), .ZN(n17399) );
  INV_X1 U52 ( .A(n17428), .ZN(n17425) );
  INV_X1 U53 ( .A(n17441), .ZN(n17438) );
  INV_X1 U54 ( .A(n17454), .ZN(n17450) );
  INV_X1 U55 ( .A(n17467), .ZN(n17464) );
  INV_X1 U56 ( .A(n17480), .ZN(n17477) );
  INV_X1 U57 ( .A(n17493), .ZN(n17490) );
  INV_X1 U58 ( .A(n17506), .ZN(n17503) );
  INV_X1 U59 ( .A(n17984), .ZN(n17966) );
  INV_X1 U60 ( .A(n17323), .ZN(n17320) );
  INV_X1 U61 ( .A(n17427), .ZN(n17424) );
  INV_X1 U62 ( .A(n17336), .ZN(n17333) );
  INV_X1 U63 ( .A(n17349), .ZN(n17346) );
  INV_X1 U64 ( .A(n17440), .ZN(n17437) );
  INV_X1 U65 ( .A(n17479), .ZN(n17476) );
  INV_X1 U66 ( .A(n17999), .ZN(n17989) );
  INV_X1 U67 ( .A(n17362), .ZN(n17359) );
  INV_X1 U68 ( .A(n17401), .ZN(n17398) );
  INV_X1 U69 ( .A(n17466), .ZN(n17463) );
  INV_X1 U70 ( .A(n17492), .ZN(n17489) );
  INV_X1 U71 ( .A(n17505), .ZN(n17502) );
  INV_X1 U72 ( .A(n17525), .ZN(n17522) );
  INV_X1 U73 ( .A(n17999), .ZN(n17990) );
  INV_X1 U74 ( .A(n17414), .ZN(n17411) );
  INV_X1 U75 ( .A(n17415), .ZN(n17412) );
  INV_X1 U76 ( .A(n17524), .ZN(n17521) );
  INV_X1 U77 ( .A(n17018), .ZN(n17009) );
  INV_X1 U78 ( .A(n17211), .ZN(n17202) );
  INV_X1 U79 ( .A(n17855), .ZN(n17836) );
  INV_X1 U80 ( .A(n17877), .ZN(n17858) );
  INV_X1 U81 ( .A(n17899), .ZN(n17880) );
  INV_X1 U82 ( .A(n17921), .ZN(n17902) );
  INV_X1 U83 ( .A(n17942), .ZN(n17923) );
  INV_X1 U84 ( .A(n17963), .ZN(n17944) );
  INV_X1 U85 ( .A(n18007), .ZN(n18004) );
  INV_X1 U86 ( .A(n18020), .ZN(n18017) );
  INV_X1 U87 ( .A(n16904), .ZN(n16901) );
  INV_X1 U88 ( .A(n16938), .ZN(n16935) );
  INV_X1 U89 ( .A(n16993), .ZN(n16990) );
  INV_X1 U90 ( .A(n17027), .ZN(n17024) );
  INV_X1 U91 ( .A(n17040), .ZN(n17037) );
  INV_X1 U92 ( .A(n17053), .ZN(n17050) );
  INV_X1 U93 ( .A(n17066), .ZN(n17063) );
  INV_X1 U94 ( .A(n17079), .ZN(n17076) );
  INV_X1 U95 ( .A(n17092), .ZN(n17089) );
  INV_X1 U96 ( .A(n17105), .ZN(n17102) );
  INV_X1 U97 ( .A(n17131), .ZN(n17128) );
  INV_X1 U98 ( .A(n17154), .ZN(n17151) );
  INV_X1 U99 ( .A(n17220), .ZN(n17217) );
  INV_X1 U100 ( .A(n17233), .ZN(n17230) );
  INV_X1 U101 ( .A(n17246), .ZN(n17243) );
  INV_X1 U102 ( .A(n17259), .ZN(n17256) );
  INV_X1 U103 ( .A(n17272), .ZN(n17269) );
  INV_X1 U104 ( .A(n17285), .ZN(n17282) );
  INV_X1 U105 ( .A(n17298), .ZN(n17295) );
  INV_X1 U106 ( .A(n17376), .ZN(n17373) );
  INV_X1 U107 ( .A(n17389), .ZN(n17386) );
  INV_X1 U108 ( .A(n17855), .ZN(n17837) );
  INV_X1 U109 ( .A(n17877), .ZN(n17859) );
  INV_X1 U110 ( .A(n17899), .ZN(n17881) );
  INV_X1 U111 ( .A(n17921), .ZN(n17903) );
  INV_X1 U112 ( .A(n17942), .ZN(n17924) );
  INV_X1 U113 ( .A(n17963), .ZN(n17945) );
  INV_X1 U114 ( .A(n17219), .ZN(n17216) );
  INV_X1 U115 ( .A(n16937), .ZN(n16934) );
  INV_X1 U116 ( .A(n17026), .ZN(n17023) );
  INV_X1 U117 ( .A(n17130), .ZN(n17127) );
  INV_X1 U118 ( .A(n18006), .ZN(n18003) );
  INV_X1 U119 ( .A(n17153), .ZN(n17150) );
  INV_X1 U120 ( .A(n16876), .ZN(n16866) );
  INV_X1 U121 ( .A(n17271), .ZN(n17268) );
  INV_X1 U122 ( .A(n17039), .ZN(n17036) );
  INV_X1 U123 ( .A(n17052), .ZN(n17049) );
  INV_X1 U124 ( .A(n17078), .ZN(n17075) );
  INV_X1 U125 ( .A(n17232), .ZN(n17229) );
  INV_X1 U126 ( .A(n17245), .ZN(n17242) );
  INV_X1 U127 ( .A(n17375), .ZN(n17372) );
  INV_X1 U128 ( .A(n18019), .ZN(n18016) );
  INV_X1 U129 ( .A(n16903), .ZN(n16900) );
  INV_X1 U130 ( .A(n16992), .ZN(n16989) );
  INV_X1 U131 ( .A(n17065), .ZN(n17062) );
  INV_X1 U132 ( .A(n17091), .ZN(n17088) );
  INV_X1 U133 ( .A(n17104), .ZN(n17101) );
  INV_X1 U134 ( .A(n17258), .ZN(n17255) );
  INV_X1 U135 ( .A(n17284), .ZN(n17281) );
  INV_X1 U136 ( .A(n17297), .ZN(n17294) );
  INV_X1 U137 ( .A(n17388), .ZN(n17385) );
  INV_X1 U138 ( .A(n17117), .ZN(n17114) );
  INV_X1 U139 ( .A(n17310), .ZN(n17307) );
  INV_X1 U140 ( .A(n17118), .ZN(n17115) );
  INV_X1 U141 ( .A(n17311), .ZN(n17308) );
  INV_X1 U142 ( .A(n16929), .ZN(n16920) );
  INV_X1 U143 ( .A(n16876), .ZN(n16867) );
  INV_X1 U144 ( .A(n16954), .ZN(n16945) );
  INV_X1 U145 ( .A(n17180), .ZN(n17171) );
  BUF_X1 U146 ( .A(n17518), .Z(n17525) );
  BUF_X1 U147 ( .A(n17317), .Z(n17323) );
  BUF_X1 U148 ( .A(n17330), .Z(n17336) );
  BUF_X1 U149 ( .A(n17343), .Z(n17349) );
  BUF_X1 U150 ( .A(n17356), .Z(n17362) );
  BUF_X1 U151 ( .A(n17421), .Z(n17427) );
  BUF_X1 U152 ( .A(n17434), .Z(n17440) );
  BUF_X1 U153 ( .A(n17447), .Z(n17453) );
  BUF_X1 U154 ( .A(n17460), .Z(n17466) );
  BUF_X1 U155 ( .A(n17473), .Z(n17479) );
  BUF_X1 U156 ( .A(n17486), .Z(n17492) );
  BUF_X1 U157 ( .A(n17499), .Z(n17505) );
  BUF_X1 U158 ( .A(n17395), .Z(n17401) );
  BUF_X1 U159 ( .A(n17408), .Z(n17414) );
  BUF_X1 U160 ( .A(n17317), .Z(n17324) );
  BUF_X1 U161 ( .A(n17330), .Z(n17337) );
  BUF_X1 U162 ( .A(n17343), .Z(n17350) );
  BUF_X1 U163 ( .A(n17356), .Z(n17363) );
  BUF_X1 U164 ( .A(n17421), .Z(n17428) );
  BUF_X1 U165 ( .A(n17434), .Z(n17441) );
  BUF_X1 U166 ( .A(n17447), .Z(n17454) );
  BUF_X1 U167 ( .A(n17460), .Z(n17467) );
  BUF_X1 U168 ( .A(n17473), .Z(n17480) );
  BUF_X1 U169 ( .A(n17486), .Z(n17493) );
  BUF_X1 U170 ( .A(n17499), .Z(n17506) );
  BUF_X1 U171 ( .A(n17518), .Z(n17524) );
  BUF_X1 U172 ( .A(n17395), .Z(n17402) );
  BUF_X1 U173 ( .A(n17408), .Z(n17415) );
  BUF_X1 U174 ( .A(n17201), .Z(n17200) );
  BUF_X1 U175 ( .A(n17008), .Z(n17007) );
  BUF_X1 U176 ( .A(n17318), .Z(n17325) );
  BUF_X1 U177 ( .A(n17331), .Z(n17338) );
  BUF_X1 U178 ( .A(n17344), .Z(n17351) );
  BUF_X1 U179 ( .A(n17357), .Z(n17364) );
  BUF_X1 U180 ( .A(n17422), .Z(n17429) );
  BUF_X1 U181 ( .A(n17435), .Z(n17442) );
  BUF_X1 U182 ( .A(n17448), .Z(n17455) );
  BUF_X1 U183 ( .A(n17461), .Z(n17468) );
  BUF_X1 U184 ( .A(n17474), .Z(n17481) );
  BUF_X1 U185 ( .A(n17487), .Z(n17494) );
  BUF_X1 U186 ( .A(n17500), .Z(n17507) );
  BUF_X1 U187 ( .A(n17519), .Z(n17526) );
  BUF_X1 U188 ( .A(n17396), .Z(n17403) );
  BUF_X1 U189 ( .A(n17409), .Z(n17416) );
  BUF_X1 U190 ( .A(n17019), .Z(n17018) );
  BUF_X1 U191 ( .A(n17212), .Z(n17211) );
  BUF_X1 U192 ( .A(n17317), .Z(n17322) );
  BUF_X1 U193 ( .A(n17330), .Z(n17335) );
  BUF_X1 U194 ( .A(n17343), .Z(n17348) );
  BUF_X1 U195 ( .A(n17356), .Z(n17361) );
  BUF_X1 U196 ( .A(n17395), .Z(n17400) );
  BUF_X1 U197 ( .A(n17408), .Z(n17413) );
  BUF_X1 U198 ( .A(n17008), .Z(n17000) );
  BUF_X1 U199 ( .A(n17201), .Z(n17193) );
  BUF_X1 U200 ( .A(n17421), .Z(n17426) );
  BUF_X1 U201 ( .A(n17434), .Z(n17439) );
  BUF_X1 U202 ( .A(n17447), .Z(n17452) );
  BUF_X1 U203 ( .A(n17460), .Z(n17465) );
  BUF_X1 U204 ( .A(n17473), .Z(n17478) );
  BUF_X1 U205 ( .A(n17486), .Z(n17491) );
  BUF_X1 U206 ( .A(n17499), .Z(n17504) );
  BUF_X1 U207 ( .A(n17518), .Z(n17523) );
  BUF_X1 U208 ( .A(n17015), .Z(n17016) );
  BUF_X1 U209 ( .A(n17208), .Z(n17209) );
  BUF_X1 U210 ( .A(n17000), .Z(n17006) );
  BUF_X1 U211 ( .A(n17193), .Z(n17199) );
  BUF_X1 U212 ( .A(n17019), .Z(n17015) );
  BUF_X1 U213 ( .A(n17212), .Z(n17208) );
  BUF_X1 U214 ( .A(n17002), .Z(n17005) );
  BUF_X1 U215 ( .A(n17195), .Z(n17198) );
  BUF_X1 U216 ( .A(n17019), .Z(n17013) );
  BUF_X1 U217 ( .A(n17212), .Z(n17206) );
  BUF_X1 U218 ( .A(n17001), .Z(n17003) );
  BUF_X1 U219 ( .A(n17194), .Z(n17196) );
  BUF_X1 U220 ( .A(n17019), .Z(n17012) );
  BUF_X1 U221 ( .A(n17212), .Z(n17205) );
  BUF_X1 U222 ( .A(n17008), .Z(n17002) );
  BUF_X1 U223 ( .A(n17201), .Z(n17195) );
  BUF_X1 U224 ( .A(n17019), .Z(n17011) );
  BUF_X1 U225 ( .A(n17212), .Z(n17204) );
  BUF_X1 U226 ( .A(n17008), .Z(n17001) );
  BUF_X1 U227 ( .A(n17201), .Z(n17194) );
  BUF_X1 U228 ( .A(n17019), .Z(n17010) );
  BUF_X1 U229 ( .A(n17212), .Z(n17203) );
  BUF_X1 U230 ( .A(n17002), .Z(n17004) );
  BUF_X1 U231 ( .A(n17019), .Z(n17014) );
  BUF_X1 U232 ( .A(n17195), .Z(n17197) );
  BUF_X1 U233 ( .A(n17212), .Z(n17207) );
  BUF_X1 U234 ( .A(n17986), .Z(n17991) );
  BUF_X1 U235 ( .A(n17986), .Z(n17992) );
  BUF_X1 U236 ( .A(n17422), .Z(n17431) );
  BUF_X1 U237 ( .A(n17435), .Z(n17444) );
  BUF_X1 U238 ( .A(n17448), .Z(n17457) );
  BUF_X1 U239 ( .A(n17461), .Z(n17470) );
  BUF_X1 U240 ( .A(n17474), .Z(n17483) );
  BUF_X1 U241 ( .A(n17487), .Z(n17496) );
  BUF_X1 U242 ( .A(n17500), .Z(n17509) );
  BUF_X1 U243 ( .A(n17519), .Z(n17528) );
  BUF_X1 U244 ( .A(n17318), .Z(n17327) );
  BUF_X1 U245 ( .A(n17331), .Z(n17340) );
  BUF_X1 U246 ( .A(n17344), .Z(n17353) );
  BUF_X1 U247 ( .A(n17357), .Z(n17366) );
  BUF_X1 U248 ( .A(n17318), .Z(n17326) );
  BUF_X1 U249 ( .A(n17331), .Z(n17339) );
  BUF_X1 U250 ( .A(n17344), .Z(n17352) );
  BUF_X1 U251 ( .A(n17357), .Z(n17365) );
  BUF_X1 U252 ( .A(n17422), .Z(n17430) );
  BUF_X1 U253 ( .A(n17435), .Z(n17443) );
  BUF_X1 U254 ( .A(n17448), .Z(n17456) );
  BUF_X1 U255 ( .A(n17461), .Z(n17469) );
  BUF_X1 U256 ( .A(n17474), .Z(n17482) );
  BUF_X1 U257 ( .A(n17487), .Z(n17495) );
  BUF_X1 U258 ( .A(n17500), .Z(n17508) );
  BUF_X1 U259 ( .A(n17519), .Z(n17527) );
  BUF_X1 U260 ( .A(n17988), .Z(n17998) );
  BUF_X1 U261 ( .A(n17988), .Z(n17997) );
  BUF_X1 U262 ( .A(n17396), .Z(n17405) );
  BUF_X1 U263 ( .A(n17409), .Z(n17418) );
  BUF_X1 U264 ( .A(n17987), .Z(n17996) );
  BUF_X1 U265 ( .A(n17987), .Z(n17994) );
  BUF_X1 U266 ( .A(n17987), .Z(n17995) );
  BUF_X1 U267 ( .A(n17986), .Z(n17993) );
  BUF_X1 U268 ( .A(n17396), .Z(n17404) );
  BUF_X1 U269 ( .A(n17409), .Z(n17417) );
  BUF_X1 U270 ( .A(n17423), .Z(n17432) );
  BUF_X1 U271 ( .A(n17436), .Z(n17445) );
  BUF_X1 U272 ( .A(n17449), .Z(n17458) );
  BUF_X1 U273 ( .A(n17462), .Z(n17471) );
  BUF_X1 U274 ( .A(n17475), .Z(n17484) );
  BUF_X1 U275 ( .A(n17488), .Z(n17497) );
  BUF_X1 U276 ( .A(n17501), .Z(n17510) );
  BUF_X1 U277 ( .A(n17520), .Z(n17529) );
  BUF_X1 U278 ( .A(n17319), .Z(n17328) );
  BUF_X1 U279 ( .A(n17332), .Z(n17341) );
  BUF_X1 U280 ( .A(n17345), .Z(n17354) );
  BUF_X1 U281 ( .A(n17358), .Z(n17367) );
  BUF_X1 U282 ( .A(n17319), .Z(n17329) );
  BUF_X1 U283 ( .A(n17332), .Z(n17342) );
  BUF_X1 U284 ( .A(n17345), .Z(n17355) );
  BUF_X1 U285 ( .A(n17358), .Z(n17368) );
  BUF_X1 U286 ( .A(n17423), .Z(n17433) );
  BUF_X1 U287 ( .A(n17436), .Z(n17446) );
  BUF_X1 U288 ( .A(n17449), .Z(n17459) );
  BUF_X1 U289 ( .A(n17462), .Z(n17472) );
  BUF_X1 U290 ( .A(n17475), .Z(n17485) );
  BUF_X1 U291 ( .A(n17488), .Z(n17498) );
  BUF_X1 U292 ( .A(n17501), .Z(n17511) );
  BUF_X1 U293 ( .A(n17520), .Z(n17530) );
  BUF_X1 U294 ( .A(n17397), .Z(n17406) );
  BUF_X1 U295 ( .A(n17410), .Z(n17419) );
  BUF_X1 U296 ( .A(n17397), .Z(n17407) );
  BUF_X1 U297 ( .A(n17410), .Z(n17420) );
  BUF_X1 U298 ( .A(n17012), .Z(n17017) );
  BUF_X1 U299 ( .A(n17205), .Z(n17210) );
  BUF_X1 U300 ( .A(n17988), .Z(n17999) );
  INV_X1 U301 ( .A(n18052), .ZN(n18039) );
  INV_X1 U302 ( .A(n18051), .ZN(n18035) );
  INV_X1 U303 ( .A(n18051), .ZN(n18036) );
  INV_X1 U304 ( .A(n18052), .ZN(n18041) );
  INV_X1 U305 ( .A(n18052), .ZN(n18040) );
  INV_X1 U306 ( .A(n18052), .ZN(n18038) );
  INV_X1 U307 ( .A(n16695), .ZN(n16691) );
  INV_X1 U308 ( .A(n17580), .ZN(n17576) );
  INV_X1 U309 ( .A(n17834), .ZN(n17824) );
  INV_X1 U310 ( .A(n17558), .ZN(n17548) );
  INV_X1 U311 ( .A(n17544), .ZN(n17534) );
  INV_X1 U312 ( .A(n17572), .ZN(n17562) );
  INV_X1 U313 ( .A(n17599), .ZN(n17589) );
  INV_X1 U314 ( .A(n17613), .ZN(n17603) );
  INV_X1 U315 ( .A(n17627), .ZN(n17617) );
  INV_X1 U316 ( .A(n17627), .ZN(n17618) );
  INV_X1 U317 ( .A(n18053), .ZN(n18044) );
  BUF_X1 U318 ( .A(n12578), .Z(n16322) );
  BUF_X1 U319 ( .A(n12543), .Z(n16394) );
  BUF_X1 U320 ( .A(n12619), .Z(n16247) );
  BUF_X1 U321 ( .A(n12578), .Z(n16323) );
  BUF_X1 U322 ( .A(n12543), .Z(n16395) );
  BUF_X1 U323 ( .A(n12619), .Z(n16248) );
  BUF_X1 U324 ( .A(n10590), .Z(n16574) );
  BUF_X1 U325 ( .A(n10536), .Z(n16658) );
  BUF_X1 U326 ( .A(n10642), .Z(n16499) );
  BUF_X1 U327 ( .A(n10590), .Z(n16575) );
  BUF_X1 U328 ( .A(n10536), .Z(n16659) );
  BUF_X1 U329 ( .A(n10642), .Z(n16500) );
  INV_X1 U330 ( .A(n18053), .ZN(n18043) );
  INV_X1 U331 ( .A(n18053), .ZN(n18042) );
  BUF_X1 U332 ( .A(n12553), .Z(n16373) );
  BUF_X1 U333 ( .A(n12553), .Z(n16374) );
  BUF_X1 U334 ( .A(n10556), .Z(n16625) );
  BUF_X1 U335 ( .A(n10556), .Z(n16626) );
  INV_X1 U336 ( .A(n17544), .ZN(n17535) );
  INV_X1 U337 ( .A(n17558), .ZN(n17549) );
  INV_X1 U338 ( .A(n17572), .ZN(n17563) );
  INV_X1 U339 ( .A(n17599), .ZN(n17590) );
  INV_X1 U340 ( .A(n17613), .ZN(n17604) );
  BUF_X1 U341 ( .A(n12566), .Z(n16352) );
  BUF_X1 U342 ( .A(n12566), .Z(n16353) );
  BUF_X1 U343 ( .A(n10573), .Z(n16604) );
  BUF_X1 U344 ( .A(n10573), .Z(n16605) );
  BUF_X1 U345 ( .A(n12616), .Z(n16256) );
  BUF_X1 U346 ( .A(n12616), .Z(n16257) );
  BUF_X1 U347 ( .A(n10637), .Z(n16508) );
  BUF_X1 U348 ( .A(n10637), .Z(n16509) );
  BUF_X1 U349 ( .A(n12576), .Z(n16328) );
  BUF_X1 U350 ( .A(n12541), .Z(n16400) );
  BUF_X1 U351 ( .A(n12546), .Z(n16388) );
  BUF_X1 U352 ( .A(n12595), .Z(n16292) );
  BUF_X1 U353 ( .A(n12576), .Z(n16329) );
  BUF_X1 U354 ( .A(n12541), .Z(n16401) );
  BUF_X1 U355 ( .A(n12546), .Z(n16389) );
  BUF_X1 U356 ( .A(n12595), .Z(n16293) );
  BUF_X1 U357 ( .A(n10594), .Z(n16568) );
  BUF_X1 U358 ( .A(n10540), .Z(n16652) );
  BUF_X1 U359 ( .A(n10547), .Z(n16640) );
  BUF_X1 U360 ( .A(n10612), .Z(n16544) );
  BUF_X1 U361 ( .A(n10594), .Z(n16569) );
  BUF_X1 U362 ( .A(n10540), .Z(n16653) );
  BUF_X1 U363 ( .A(n10547), .Z(n16641) );
  BUF_X1 U364 ( .A(n10612), .Z(n16545) );
  BUF_X1 U365 ( .A(n4248), .Z(n17629) );
  BUF_X1 U366 ( .A(n4112), .Z(n17809) );
  BUF_X1 U367 ( .A(n4121), .Z(n17797) );
  BUF_X1 U368 ( .A(n4128), .Z(n17785) );
  BUF_X1 U369 ( .A(n4248), .Z(n17628) );
  BUF_X1 U370 ( .A(n4112), .Z(n17808) );
  BUF_X1 U371 ( .A(n4121), .Z(n17796) );
  BUF_X1 U372 ( .A(n4128), .Z(n17784) );
  BUF_X1 U373 ( .A(n12578), .Z(n16324) );
  BUF_X1 U374 ( .A(n12543), .Z(n16396) );
  BUF_X1 U375 ( .A(n12619), .Z(n16249) );
  BUF_X1 U376 ( .A(n10590), .Z(n16576) );
  BUF_X1 U377 ( .A(n10536), .Z(n16660) );
  BUF_X1 U378 ( .A(n10642), .Z(n16501) );
  BUF_X1 U379 ( .A(n12561), .Z(n16364) );
  BUF_X1 U380 ( .A(n12537), .Z(n16409) );
  BUF_X1 U381 ( .A(n12547), .Z(n16385) );
  BUF_X1 U382 ( .A(n12586), .Z(n16313) );
  BUF_X1 U383 ( .A(n12628), .Z(n16226) );
  BUF_X1 U384 ( .A(n12561), .Z(n16365) );
  BUF_X1 U385 ( .A(n12537), .Z(n16410) );
  BUF_X1 U386 ( .A(n12547), .Z(n16386) );
  BUF_X1 U387 ( .A(n12586), .Z(n16314) );
  BUF_X1 U388 ( .A(n12628), .Z(n16227) );
  BUF_X1 U389 ( .A(n10566), .Z(n16616) );
  BUF_X1 U390 ( .A(n10535), .Z(n16661) );
  BUF_X1 U391 ( .A(n10549), .Z(n16637) );
  BUF_X1 U392 ( .A(n10600), .Z(n16565) );
  BUF_X1 U393 ( .A(n10655), .Z(n16478) );
  BUF_X1 U394 ( .A(n10566), .Z(n16617) );
  BUF_X1 U395 ( .A(n10535), .Z(n16662) );
  BUF_X1 U396 ( .A(n10549), .Z(n16638) );
  BUF_X1 U397 ( .A(n10600), .Z(n16566) );
  BUF_X1 U398 ( .A(n10655), .Z(n16479) );
  BUF_X1 U399 ( .A(n12540), .Z(n16403) );
  BUF_X1 U400 ( .A(n12540), .Z(n16404) );
  BUF_X1 U401 ( .A(n10538), .Z(n16655) );
  BUF_X1 U402 ( .A(n10538), .Z(n16656) );
  BUF_X1 U403 ( .A(n4110), .Z(n17812) );
  BUF_X1 U404 ( .A(n4110), .Z(n17811) );
  BUF_X1 U405 ( .A(n12553), .Z(n16375) );
  BUF_X1 U406 ( .A(n10556), .Z(n16627) );
  BUF_X1 U407 ( .A(n12566), .Z(n16354) );
  BUF_X1 U408 ( .A(n10573), .Z(n16606) );
  BUF_X1 U409 ( .A(n12616), .Z(n16258) );
  BUF_X1 U410 ( .A(n10637), .Z(n16510) );
  BUF_X1 U411 ( .A(n12576), .Z(n16330) );
  BUF_X1 U412 ( .A(n12541), .Z(n16402) );
  BUF_X1 U413 ( .A(n12546), .Z(n16390) );
  BUF_X1 U414 ( .A(n12595), .Z(n16294) );
  BUF_X1 U415 ( .A(n10594), .Z(n16570) );
  BUF_X1 U416 ( .A(n10540), .Z(n16654) );
  BUF_X1 U417 ( .A(n10547), .Z(n16642) );
  BUF_X1 U418 ( .A(n10612), .Z(n16546) );
  BUF_X1 U419 ( .A(n4248), .Z(n17630) );
  BUF_X1 U420 ( .A(n4112), .Z(n17810) );
  BUF_X1 U421 ( .A(n4121), .Z(n17798) );
  BUF_X1 U422 ( .A(n4128), .Z(n17786) );
  BUF_X1 U423 ( .A(n12561), .Z(n16366) );
  BUF_X1 U424 ( .A(n12537), .Z(n16411) );
  BUF_X1 U425 ( .A(n12547), .Z(n16387) );
  BUF_X1 U426 ( .A(n12586), .Z(n16315) );
  BUF_X1 U427 ( .A(n12628), .Z(n16228) );
  BUF_X1 U428 ( .A(n10566), .Z(n16618) );
  BUF_X1 U429 ( .A(n10535), .Z(n16663) );
  BUF_X1 U430 ( .A(n10549), .Z(n16639) );
  BUF_X1 U431 ( .A(n10600), .Z(n16567) );
  BUF_X1 U432 ( .A(n10655), .Z(n16480) );
  BUF_X1 U433 ( .A(n12540), .Z(n16405) );
  BUF_X1 U434 ( .A(n10538), .Z(n16657) );
  BUF_X1 U435 ( .A(n4110), .Z(n17813) );
  BUF_X1 U436 ( .A(n18000), .Z(n18007) );
  BUF_X1 U437 ( .A(n18013), .Z(n18020) );
  BUF_X1 U438 ( .A(n16897), .Z(n16903) );
  BUF_X1 U439 ( .A(n16931), .Z(n16937) );
  BUF_X1 U440 ( .A(n18000), .Z(n18006) );
  BUF_X1 U441 ( .A(n16986), .Z(n16992) );
  BUF_X1 U442 ( .A(n17020), .Z(n17026) );
  BUF_X1 U443 ( .A(n17033), .Z(n17039) );
  BUF_X1 U444 ( .A(n17046), .Z(n17052) );
  BUF_X1 U445 ( .A(n17059), .Z(n17065) );
  BUF_X1 U446 ( .A(n17072), .Z(n17078) );
  BUF_X1 U447 ( .A(n17085), .Z(n17091) );
  BUF_X1 U448 ( .A(n17098), .Z(n17104) );
  BUF_X1 U449 ( .A(n17111), .Z(n17117) );
  BUF_X1 U450 ( .A(n17124), .Z(n17130) );
  BUF_X1 U451 ( .A(n17147), .Z(n17153) );
  BUF_X1 U452 ( .A(n17213), .Z(n17219) );
  BUF_X1 U453 ( .A(n17226), .Z(n17232) );
  BUF_X1 U454 ( .A(n17239), .Z(n17245) );
  BUF_X1 U455 ( .A(n17252), .Z(n17258) );
  BUF_X1 U456 ( .A(n17265), .Z(n17271) );
  BUF_X1 U457 ( .A(n17278), .Z(n17284) );
  BUF_X1 U458 ( .A(n17291), .Z(n17297) );
  BUF_X1 U459 ( .A(n17304), .Z(n17310) );
  BUF_X1 U460 ( .A(n17369), .Z(n17375) );
  BUF_X1 U461 ( .A(n17382), .Z(n17388) );
  BUF_X1 U462 ( .A(n18013), .Z(n18019) );
  BUF_X1 U463 ( .A(n16897), .Z(n16904) );
  BUF_X1 U464 ( .A(n16931), .Z(n16938) );
  BUF_X1 U465 ( .A(n16986), .Z(n16993) );
  BUF_X1 U466 ( .A(n17020), .Z(n17027) );
  BUF_X1 U467 ( .A(n17033), .Z(n17040) );
  BUF_X1 U468 ( .A(n17046), .Z(n17053) );
  BUF_X1 U469 ( .A(n17059), .Z(n17066) );
  BUF_X1 U470 ( .A(n17072), .Z(n17079) );
  BUF_X1 U471 ( .A(n17085), .Z(n17092) );
  BUF_X1 U472 ( .A(n17098), .Z(n17105) );
  BUF_X1 U473 ( .A(n17111), .Z(n17118) );
  BUF_X1 U474 ( .A(n17124), .Z(n17131) );
  BUF_X1 U475 ( .A(n17147), .Z(n17154) );
  BUF_X1 U476 ( .A(n17213), .Z(n17220) );
  BUF_X1 U477 ( .A(n17226), .Z(n17233) );
  BUF_X1 U478 ( .A(n17239), .Z(n17246) );
  BUF_X1 U479 ( .A(n17252), .Z(n17259) );
  BUF_X1 U480 ( .A(n17265), .Z(n17272) );
  BUF_X1 U481 ( .A(n17278), .Z(n17285) );
  BUF_X1 U482 ( .A(n17291), .Z(n17298) );
  BUF_X1 U483 ( .A(n17304), .Z(n17311) );
  BUF_X1 U484 ( .A(n17369), .Z(n17376) );
  BUF_X1 U485 ( .A(n17382), .Z(n17389) );
  BUF_X1 U486 ( .A(n17181), .Z(n17179) );
  BUF_X1 U487 ( .A(n17191), .Z(n17190) );
  BUF_X1 U488 ( .A(n16886), .Z(n16885) );
  BUF_X1 U489 ( .A(n16896), .Z(n16895) );
  BUF_X1 U490 ( .A(n16919), .Z(n16918) );
  BUF_X1 U491 ( .A(n16955), .Z(n16953) );
  BUF_X1 U492 ( .A(n16965), .Z(n16964) );
  BUF_X1 U493 ( .A(n16975), .Z(n16974) );
  BUF_X1 U494 ( .A(n16985), .Z(n16984) );
  BUF_X1 U495 ( .A(n17146), .Z(n17145) );
  BUF_X1 U496 ( .A(n17169), .Z(n17168) );
  BUF_X1 U497 ( .A(n18001), .Z(n18008) );
  BUF_X1 U498 ( .A(n18014), .Z(n18021) );
  BUF_X1 U499 ( .A(n16898), .Z(n16905) );
  BUF_X1 U500 ( .A(n16932), .Z(n16939) );
  BUF_X1 U501 ( .A(n17021), .Z(n17028) );
  BUF_X1 U502 ( .A(n17034), .Z(n17041) );
  BUF_X1 U503 ( .A(n17047), .Z(n17054) );
  BUF_X1 U504 ( .A(n17060), .Z(n17067) );
  BUF_X1 U505 ( .A(n17073), .Z(n17080) );
  BUF_X1 U506 ( .A(n17086), .Z(n17093) );
  BUF_X1 U507 ( .A(n17099), .Z(n17106) );
  BUF_X1 U508 ( .A(n17112), .Z(n17119) );
  BUF_X1 U509 ( .A(n17125), .Z(n17132) );
  BUF_X1 U510 ( .A(n17148), .Z(n17155) );
  BUF_X1 U511 ( .A(n17214), .Z(n17221) );
  BUF_X1 U512 ( .A(n17227), .Z(n17234) );
  BUF_X1 U513 ( .A(n17240), .Z(n17247) );
  BUF_X1 U514 ( .A(n17253), .Z(n17260) );
  BUF_X1 U515 ( .A(n17266), .Z(n17273) );
  BUF_X1 U516 ( .A(n17279), .Z(n17286) );
  BUF_X1 U517 ( .A(n17292), .Z(n17299) );
  BUF_X1 U518 ( .A(n17305), .Z(n17312) );
  BUF_X1 U519 ( .A(n16987), .Z(n16994) );
  BUF_X1 U520 ( .A(n17370), .Z(n17377) );
  BUF_X1 U521 ( .A(n17383), .Z(n17390) );
  BUF_X1 U522 ( .A(n16930), .Z(n16929) );
  BUF_X1 U523 ( .A(n16931), .Z(n16936) );
  BUF_X1 U524 ( .A(n17124), .Z(n17129) );
  BUF_X1 U525 ( .A(n18000), .Z(n18005) );
  BUF_X1 U526 ( .A(n18013), .Z(n18018) );
  BUF_X1 U527 ( .A(n17020), .Z(n17025) );
  BUF_X1 U528 ( .A(n17033), .Z(n17038) );
  BUF_X1 U529 ( .A(n17046), .Z(n17051) );
  BUF_X1 U530 ( .A(n17059), .Z(n17064) );
  BUF_X1 U531 ( .A(n17072), .Z(n17077) );
  BUF_X1 U532 ( .A(n17085), .Z(n17090) );
  BUF_X1 U533 ( .A(n17098), .Z(n17103) );
  BUF_X1 U534 ( .A(n17111), .Z(n17116) );
  BUF_X1 U535 ( .A(n17226), .Z(n17231) );
  BUF_X1 U536 ( .A(n17239), .Z(n17244) );
  BUF_X1 U537 ( .A(n17252), .Z(n17257) );
  BUF_X1 U538 ( .A(n17278), .Z(n17283) );
  BUF_X1 U539 ( .A(n17291), .Z(n17296) );
  BUF_X1 U540 ( .A(n17304), .Z(n17309) );
  BUF_X1 U541 ( .A(n17369), .Z(n17374) );
  BUF_X1 U542 ( .A(n17382), .Z(n17387) );
  BUF_X1 U543 ( .A(n16896), .Z(n16888) );
  BUF_X1 U544 ( .A(n16955), .Z(n16946) );
  BUF_X1 U545 ( .A(n16965), .Z(n16957) );
  BUF_X1 U546 ( .A(n16985), .Z(n16977) );
  BUF_X1 U547 ( .A(n17146), .Z(n17138) );
  BUF_X1 U548 ( .A(n17181), .Z(n17172) );
  BUF_X1 U549 ( .A(n16863), .Z(n16868) );
  BUF_X1 U550 ( .A(n16886), .Z(n16878) );
  BUF_X1 U551 ( .A(n16919), .Z(n16911) );
  BUF_X1 U552 ( .A(n16975), .Z(n16967) );
  BUF_X1 U553 ( .A(n17169), .Z(n17161) );
  BUF_X1 U554 ( .A(n17191), .Z(n17183) );
  BUF_X1 U555 ( .A(n16897), .Z(n16902) );
  BUF_X1 U556 ( .A(n17147), .Z(n17152) );
  BUF_X1 U557 ( .A(n16986), .Z(n16991) );
  BUF_X1 U558 ( .A(n17213), .Z(n17218) );
  BUF_X1 U559 ( .A(n17265), .Z(n17270) );
  BUF_X1 U560 ( .A(n16926), .Z(n16927) );
  BUF_X1 U561 ( .A(n16878), .Z(n16884) );
  BUF_X1 U562 ( .A(n16911), .Z(n16917) );
  BUF_X1 U563 ( .A(n16967), .Z(n16973) );
  BUF_X1 U564 ( .A(n17161), .Z(n17167) );
  BUF_X1 U565 ( .A(n17183), .Z(n17189) );
  BUF_X1 U566 ( .A(n16888), .Z(n16894) );
  BUF_X1 U567 ( .A(n16946), .Z(n16952) );
  BUF_X1 U568 ( .A(n16957), .Z(n16963) );
  BUF_X1 U569 ( .A(n16977), .Z(n16983) );
  BUF_X1 U570 ( .A(n17138), .Z(n17144) );
  BUF_X1 U571 ( .A(n17172), .Z(n17178) );
  BUF_X1 U572 ( .A(n16930), .Z(n16926) );
  BUF_X1 U573 ( .A(n16880), .Z(n16883) );
  BUF_X1 U574 ( .A(n16913), .Z(n16916) );
  BUF_X1 U575 ( .A(n16969), .Z(n16972) );
  BUF_X1 U576 ( .A(n17163), .Z(n17166) );
  BUF_X1 U577 ( .A(n17185), .Z(n17188) );
  BUF_X1 U578 ( .A(n16890), .Z(n16893) );
  BUF_X1 U579 ( .A(n16948), .Z(n16951) );
  BUF_X1 U580 ( .A(n16959), .Z(n16962) );
  BUF_X1 U581 ( .A(n16979), .Z(n16982) );
  BUF_X1 U582 ( .A(n17140), .Z(n17143) );
  BUF_X1 U583 ( .A(n17174), .Z(n17177) );
  BUF_X1 U584 ( .A(n16930), .Z(n16924) );
  BUF_X1 U585 ( .A(n16879), .Z(n16881) );
  BUF_X1 U586 ( .A(n16912), .Z(n16914) );
  BUF_X1 U587 ( .A(n16968), .Z(n16970) );
  BUF_X1 U588 ( .A(n17162), .Z(n17164) );
  BUF_X1 U589 ( .A(n17184), .Z(n17186) );
  BUF_X1 U590 ( .A(n16889), .Z(n16891) );
  BUF_X1 U591 ( .A(n16947), .Z(n16949) );
  BUF_X1 U592 ( .A(n16958), .Z(n16960) );
  BUF_X1 U593 ( .A(n16978), .Z(n16980) );
  BUF_X1 U594 ( .A(n17139), .Z(n17141) );
  BUF_X1 U595 ( .A(n17173), .Z(n17175) );
  BUF_X1 U596 ( .A(n16930), .Z(n16923) );
  BUF_X1 U597 ( .A(n16886), .Z(n16880) );
  BUF_X1 U598 ( .A(n16919), .Z(n16913) );
  BUF_X1 U599 ( .A(n16975), .Z(n16969) );
  BUF_X1 U600 ( .A(n17169), .Z(n17163) );
  BUF_X1 U601 ( .A(n17191), .Z(n17185) );
  BUF_X1 U602 ( .A(n16896), .Z(n16890) );
  BUF_X1 U603 ( .A(n16955), .Z(n16948) );
  BUF_X1 U604 ( .A(n16965), .Z(n16959) );
  BUF_X1 U605 ( .A(n16985), .Z(n16979) );
  BUF_X1 U606 ( .A(n17146), .Z(n17140) );
  BUF_X1 U607 ( .A(n17181), .Z(n17174) );
  BUF_X1 U608 ( .A(n16930), .Z(n16922) );
  BUF_X1 U609 ( .A(n16919), .Z(n16912) );
  BUF_X1 U610 ( .A(n17191), .Z(n17184) );
  BUF_X1 U611 ( .A(n16896), .Z(n16889) );
  BUF_X1 U612 ( .A(n16955), .Z(n16947) );
  BUF_X1 U613 ( .A(n16965), .Z(n16958) );
  BUF_X1 U614 ( .A(n16985), .Z(n16978) );
  BUF_X1 U615 ( .A(n17146), .Z(n17139) );
  BUF_X1 U616 ( .A(n17181), .Z(n17173) );
  BUF_X1 U617 ( .A(n16886), .Z(n16879) );
  BUF_X1 U618 ( .A(n16975), .Z(n16968) );
  BUF_X1 U619 ( .A(n17169), .Z(n17162) );
  BUF_X1 U620 ( .A(n16930), .Z(n16921) );
  BUF_X1 U621 ( .A(n16880), .Z(n16882) );
  BUF_X1 U622 ( .A(n16890), .Z(n16892) );
  BUF_X1 U623 ( .A(n16913), .Z(n16915) );
  BUF_X1 U624 ( .A(n16930), .Z(n16925) );
  BUF_X1 U625 ( .A(n16948), .Z(n16950) );
  BUF_X1 U626 ( .A(n16959), .Z(n16961) );
  BUF_X1 U627 ( .A(n16969), .Z(n16971) );
  BUF_X1 U628 ( .A(n16979), .Z(n16981) );
  BUF_X1 U629 ( .A(n17140), .Z(n17142) );
  BUF_X1 U630 ( .A(n17163), .Z(n17165) );
  BUF_X1 U631 ( .A(n17174), .Z(n17176) );
  BUF_X1 U632 ( .A(n17185), .Z(n17187) );
  BUF_X1 U633 ( .A(n16865), .Z(n16874) );
  BUF_X1 U634 ( .A(n17021), .Z(n17030) );
  BUF_X1 U635 ( .A(n17034), .Z(n17043) );
  BUF_X1 U636 ( .A(n17047), .Z(n17056) );
  BUF_X1 U637 ( .A(n17060), .Z(n17069) );
  BUF_X1 U638 ( .A(n17073), .Z(n17082) );
  BUF_X1 U639 ( .A(n17086), .Z(n17095) );
  BUF_X1 U640 ( .A(n17099), .Z(n17108) );
  BUF_X1 U641 ( .A(n17112), .Z(n17121) );
  BUF_X1 U642 ( .A(n17214), .Z(n17223) );
  BUF_X1 U643 ( .A(n17227), .Z(n17236) );
  BUF_X1 U644 ( .A(n17240), .Z(n17249) );
  BUF_X1 U645 ( .A(n17253), .Z(n17262) );
  BUF_X1 U646 ( .A(n17266), .Z(n17275) );
  BUF_X1 U647 ( .A(n17279), .Z(n17288) );
  BUF_X1 U648 ( .A(n17292), .Z(n17301) );
  BUF_X1 U649 ( .A(n17305), .Z(n17314) );
  BUF_X1 U650 ( .A(n16864), .Z(n16873) );
  BUF_X1 U651 ( .A(n16898), .Z(n16907) );
  BUF_X1 U652 ( .A(n16932), .Z(n16941) );
  BUF_X1 U653 ( .A(n17125), .Z(n17134) );
  BUF_X1 U654 ( .A(n17148), .Z(n17157) );
  BUF_X1 U655 ( .A(n18001), .Z(n18010) );
  BUF_X1 U656 ( .A(n18014), .Z(n18023) );
  BUF_X1 U657 ( .A(n16864), .Z(n16871) );
  BUF_X1 U658 ( .A(n18001), .Z(n18009) );
  BUF_X1 U659 ( .A(n18014), .Z(n18022) );
  BUF_X1 U660 ( .A(n16863), .Z(n16870) );
  BUF_X1 U661 ( .A(n16863), .Z(n16869) );
  BUF_X1 U662 ( .A(n16864), .Z(n16872) );
  BUF_X1 U663 ( .A(n16898), .Z(n16906) );
  BUF_X1 U664 ( .A(n16932), .Z(n16940) );
  BUF_X1 U665 ( .A(n17021), .Z(n17029) );
  BUF_X1 U666 ( .A(n17034), .Z(n17042) );
  BUF_X1 U667 ( .A(n17047), .Z(n17055) );
  BUF_X1 U668 ( .A(n17060), .Z(n17068) );
  BUF_X1 U669 ( .A(n17073), .Z(n17081) );
  BUF_X1 U670 ( .A(n17086), .Z(n17094) );
  BUF_X1 U671 ( .A(n17099), .Z(n17107) );
  BUF_X1 U672 ( .A(n17112), .Z(n17120) );
  BUF_X1 U673 ( .A(n17125), .Z(n17133) );
  BUF_X1 U674 ( .A(n17148), .Z(n17156) );
  BUF_X1 U675 ( .A(n17214), .Z(n17222) );
  BUF_X1 U676 ( .A(n17227), .Z(n17235) );
  BUF_X1 U677 ( .A(n17240), .Z(n17248) );
  BUF_X1 U678 ( .A(n17253), .Z(n17261) );
  BUF_X1 U679 ( .A(n17266), .Z(n17274) );
  BUF_X1 U680 ( .A(n17279), .Z(n17287) );
  BUF_X1 U681 ( .A(n17292), .Z(n17300) );
  BUF_X1 U682 ( .A(n17305), .Z(n17313) );
  BUF_X1 U683 ( .A(n16865), .Z(n16875) );
  BUF_X1 U684 ( .A(n17370), .Z(n17379) );
  BUF_X1 U685 ( .A(n17383), .Z(n17392) );
  BUF_X1 U686 ( .A(n16987), .Z(n16996) );
  BUF_X1 U687 ( .A(n16987), .Z(n16995) );
  BUF_X1 U688 ( .A(n17370), .Z(n17378) );
  BUF_X1 U689 ( .A(n17383), .Z(n17391) );
  BUF_X1 U690 ( .A(n18002), .Z(n18012) );
  BUF_X1 U691 ( .A(n18015), .Z(n18025) );
  BUF_X1 U692 ( .A(n17022), .Z(n17031) );
  BUF_X1 U693 ( .A(n17035), .Z(n17044) );
  BUF_X1 U694 ( .A(n17048), .Z(n17057) );
  BUF_X1 U695 ( .A(n17061), .Z(n17070) );
  BUF_X1 U696 ( .A(n17074), .Z(n17083) );
  BUF_X1 U697 ( .A(n17087), .Z(n17096) );
  BUF_X1 U698 ( .A(n17100), .Z(n17109) );
  BUF_X1 U699 ( .A(n17113), .Z(n17122) );
  BUF_X1 U700 ( .A(n17215), .Z(n17224) );
  BUF_X1 U701 ( .A(n17228), .Z(n17237) );
  BUF_X1 U702 ( .A(n17241), .Z(n17250) );
  BUF_X1 U703 ( .A(n17254), .Z(n17263) );
  BUF_X1 U704 ( .A(n17267), .Z(n17276) );
  BUF_X1 U705 ( .A(n17280), .Z(n17289) );
  BUF_X1 U706 ( .A(n17293), .Z(n17302) );
  BUF_X1 U707 ( .A(n17306), .Z(n17315) );
  BUF_X1 U708 ( .A(n16899), .Z(n16908) );
  BUF_X1 U709 ( .A(n16933), .Z(n16942) );
  BUF_X1 U710 ( .A(n17126), .Z(n17135) );
  BUF_X1 U711 ( .A(n17149), .Z(n17158) );
  BUF_X1 U712 ( .A(n18002), .Z(n18011) );
  BUF_X1 U713 ( .A(n16899), .Z(n16909) );
  BUF_X1 U714 ( .A(n18015), .Z(n18024) );
  BUF_X1 U715 ( .A(n16933), .Z(n16943) );
  BUF_X1 U716 ( .A(n17022), .Z(n17032) );
  BUF_X1 U717 ( .A(n17035), .Z(n17045) );
  BUF_X1 U718 ( .A(n17048), .Z(n17058) );
  BUF_X1 U719 ( .A(n17061), .Z(n17071) );
  BUF_X1 U720 ( .A(n17074), .Z(n17084) );
  BUF_X1 U721 ( .A(n17087), .Z(n17097) );
  BUF_X1 U722 ( .A(n17100), .Z(n17110) );
  BUF_X1 U723 ( .A(n17113), .Z(n17123) );
  BUF_X1 U724 ( .A(n17126), .Z(n17136) );
  BUF_X1 U725 ( .A(n17149), .Z(n17159) );
  BUF_X1 U726 ( .A(n17215), .Z(n17225) );
  BUF_X1 U727 ( .A(n17228), .Z(n17238) );
  BUF_X1 U728 ( .A(n17241), .Z(n17251) );
  BUF_X1 U729 ( .A(n17254), .Z(n17264) );
  BUF_X1 U730 ( .A(n17267), .Z(n17277) );
  BUF_X1 U731 ( .A(n17280), .Z(n17290) );
  BUF_X1 U732 ( .A(n17293), .Z(n17303) );
  BUF_X1 U733 ( .A(n17306), .Z(n17316) );
  BUF_X1 U734 ( .A(n17371), .Z(n17380) );
  BUF_X1 U735 ( .A(n17384), .Z(n17393) );
  BUF_X1 U736 ( .A(n16988), .Z(n16997) );
  BUF_X1 U737 ( .A(n16988), .Z(n16998) );
  BUF_X1 U738 ( .A(n17371), .Z(n17381) );
  BUF_X1 U739 ( .A(n17384), .Z(n17394) );
  BUF_X1 U740 ( .A(n16923), .Z(n16928) );
  BUF_X1 U741 ( .A(n16865), .Z(n16876) );
  BUF_X1 U742 ( .A(n16955), .Z(n16954) );
  BUF_X1 U743 ( .A(n17181), .Z(n17180) );
  BUF_X1 U744 ( .A(n4329), .Z(n17317) );
  BUF_X1 U745 ( .A(n4326), .Z(n17330) );
  BUF_X1 U746 ( .A(n4323), .Z(n17343) );
  BUF_X1 U747 ( .A(n4320), .Z(n17356) );
  BUF_X1 U748 ( .A(n4301), .Z(n17421) );
  BUF_X1 U749 ( .A(n4298), .Z(n17434) );
  BUF_X1 U750 ( .A(n4291), .Z(n17447) );
  BUF_X1 U751 ( .A(n4288), .Z(n17460) );
  BUF_X1 U752 ( .A(n4285), .Z(n17473) );
  BUF_X1 U753 ( .A(n4282), .Z(n17486) );
  BUF_X1 U754 ( .A(n4279), .Z(n17499) );
  BUF_X1 U755 ( .A(n4275), .Z(n17518) );
  BUF_X1 U756 ( .A(n4329), .Z(n17318) );
  BUF_X1 U757 ( .A(n4326), .Z(n17331) );
  BUF_X1 U758 ( .A(n4323), .Z(n17344) );
  BUF_X1 U759 ( .A(n4320), .Z(n17357) );
  BUF_X1 U760 ( .A(n4301), .Z(n17422) );
  BUF_X1 U761 ( .A(n4298), .Z(n17435) );
  BUF_X1 U762 ( .A(n4291), .Z(n17448) );
  BUF_X1 U763 ( .A(n4288), .Z(n17461) );
  BUF_X1 U764 ( .A(n4285), .Z(n17474) );
  BUF_X1 U765 ( .A(n4282), .Z(n17487) );
  BUF_X1 U766 ( .A(n4279), .Z(n17500) );
  BUF_X1 U767 ( .A(n4275), .Z(n17519) );
  BUF_X1 U768 ( .A(n4067), .Z(n17988) );
  BUF_X1 U769 ( .A(n4067), .Z(n17987) );
  BUF_X1 U770 ( .A(n4067), .Z(n17986) );
  BUF_X1 U771 ( .A(n4309), .Z(n17395) );
  BUF_X1 U772 ( .A(n4306), .Z(n17408) );
  BUF_X1 U773 ( .A(n4309), .Z(n17396) );
  BUF_X1 U774 ( .A(n4306), .Z(n17409) );
  BUF_X1 U775 ( .A(n4329), .Z(n17319) );
  BUF_X1 U776 ( .A(n4326), .Z(n17332) );
  BUF_X1 U777 ( .A(n4323), .Z(n17345) );
  BUF_X1 U778 ( .A(n4320), .Z(n17358) );
  BUF_X1 U779 ( .A(n4301), .Z(n17423) );
  BUF_X1 U780 ( .A(n4298), .Z(n17436) );
  BUF_X1 U781 ( .A(n4291), .Z(n17449) );
  BUF_X1 U782 ( .A(n4288), .Z(n17462) );
  BUF_X1 U783 ( .A(n4285), .Z(n17475) );
  BUF_X1 U784 ( .A(n4282), .Z(n17488) );
  BUF_X1 U785 ( .A(n4279), .Z(n17501) );
  BUF_X1 U786 ( .A(n4275), .Z(n17520) );
  BUF_X1 U787 ( .A(n4309), .Z(n17397) );
  BUF_X1 U788 ( .A(n4306), .Z(n17410) );
  INV_X1 U789 ( .A(n16999), .ZN(n17008) );
  INV_X1 U790 ( .A(n4420), .ZN(n17019) );
  INV_X1 U791 ( .A(n17192), .ZN(n17201) );
  INV_X1 U792 ( .A(n4362), .ZN(n17212) );
  INV_X1 U793 ( .A(n18051), .ZN(n18034) );
  INV_X1 U794 ( .A(n18051), .ZN(n18037) );
  INV_X1 U795 ( .A(n17834), .ZN(n17823) );
  OAI21_X1 U796 ( .B1(n14061), .B2(n14063), .A(n18039), .ZN(n4070) );
  BUF_X1 U797 ( .A(n4182), .Z(n17719) );
  BUF_X1 U798 ( .A(n4226), .Z(n17659) );
  BUF_X1 U799 ( .A(n4182), .Z(n17718) );
  BUF_X1 U800 ( .A(n4226), .Z(n17658) );
  BUF_X1 U801 ( .A(n4117), .Z(n17803) );
  BUF_X1 U802 ( .A(n4117), .Z(n17802) );
  BUF_X1 U803 ( .A(n4108), .Z(n17815) );
  BUF_X1 U804 ( .A(n4108), .Z(n17814) );
  BUF_X1 U805 ( .A(n12562), .Z(n16361) );
  BUF_X1 U806 ( .A(n12573), .Z(n16334) );
  BUF_X1 U807 ( .A(n12568), .Z(n16346) );
  BUF_X1 U808 ( .A(n12538), .Z(n16406) );
  BUF_X1 U809 ( .A(n12548), .Z(n16382) );
  BUF_X1 U810 ( .A(n12604), .Z(n16274) );
  BUF_X1 U811 ( .A(n12587), .Z(n16310) );
  BUF_X1 U812 ( .A(n12592), .Z(n16298) );
  BUF_X1 U813 ( .A(n12597), .Z(n16286) );
  BUF_X1 U814 ( .A(n12613), .Z(n16262) );
  BUF_X1 U815 ( .A(n12629), .Z(n16223) );
  BUF_X1 U816 ( .A(n12562), .Z(n16362) );
  BUF_X1 U817 ( .A(n12573), .Z(n16335) );
  BUF_X1 U818 ( .A(n12568), .Z(n16347) );
  BUF_X1 U819 ( .A(n12538), .Z(n16407) );
  BUF_X1 U820 ( .A(n12548), .Z(n16383) );
  BUF_X1 U821 ( .A(n12604), .Z(n16275) );
  BUF_X1 U822 ( .A(n12587), .Z(n16311) );
  BUF_X1 U823 ( .A(n12592), .Z(n16299) );
  BUF_X1 U824 ( .A(n12597), .Z(n16287) );
  BUF_X1 U825 ( .A(n12613), .Z(n16263) );
  BUF_X1 U826 ( .A(n12629), .Z(n16224) );
  BUF_X1 U827 ( .A(n10567), .Z(n16613) );
  BUF_X1 U828 ( .A(n10583), .Z(n16586) );
  BUF_X1 U829 ( .A(n10576), .Z(n16598) );
  BUF_X1 U830 ( .A(n10550), .Z(n16634) );
  BUF_X1 U831 ( .A(n10543), .Z(n16646) );
  BUF_X1 U832 ( .A(n10615), .Z(n16538) );
  BUF_X1 U833 ( .A(n10622), .Z(n16526) );
  BUF_X1 U834 ( .A(n10601), .Z(n16562) );
  BUF_X1 U835 ( .A(n10608), .Z(n16550) );
  BUF_X1 U836 ( .A(n10633), .Z(n16514) );
  BUF_X1 U837 ( .A(n10656), .Z(n16475) );
  BUF_X1 U838 ( .A(n10567), .Z(n16614) );
  BUF_X1 U839 ( .A(n10583), .Z(n16587) );
  BUF_X1 U840 ( .A(n10576), .Z(n16599) );
  BUF_X1 U841 ( .A(n10550), .Z(n16635) );
  BUF_X1 U842 ( .A(n10543), .Z(n16647) );
  BUF_X1 U843 ( .A(n10615), .Z(n16539) );
  BUF_X1 U844 ( .A(n10622), .Z(n16527) );
  BUF_X1 U845 ( .A(n10601), .Z(n16563) );
  BUF_X1 U846 ( .A(n10608), .Z(n16551) );
  BUF_X1 U847 ( .A(n10633), .Z(n16515) );
  BUF_X1 U848 ( .A(n10656), .Z(n16476) );
  BUF_X1 U849 ( .A(n4162), .Z(n17743) );
  BUF_X1 U850 ( .A(n4162), .Z(n17742) );
  BUF_X1 U851 ( .A(n12617), .Z(n16253) );
  BUF_X1 U852 ( .A(n12617), .Z(n16254) );
  BUF_X1 U853 ( .A(n10639), .Z(n16505) );
  BUF_X1 U854 ( .A(n10639), .Z(n16506) );
  OAI21_X1 U855 ( .B1(n14074), .B2(n14236), .A(n18041), .ZN(n4329) );
  OAI21_X1 U856 ( .B1(n14073), .B2(n14236), .A(n18041), .ZN(n4326) );
  OAI21_X1 U857 ( .B1(n14072), .B2(n14236), .A(n18040), .ZN(n4323) );
  OAI21_X1 U858 ( .B1(n14070), .B2(n14236), .A(n18041), .ZN(n4320) );
  OAI21_X1 U859 ( .B1(n12414), .B2(n14236), .A(n18040), .ZN(n4301) );
  OAI21_X1 U860 ( .B1(n14058), .B2(n14236), .A(n18040), .ZN(n4298) );
  OAI21_X1 U861 ( .B1(n14228), .B2(n14236), .A(n18040), .ZN(n4291) );
  OAI21_X1 U862 ( .B1(n14226), .B2(n14236), .A(n18040), .ZN(n4288) );
  OAI21_X1 U863 ( .B1(n14222), .B2(n14236), .A(n18040), .ZN(n4285) );
  OAI21_X1 U864 ( .B1(n14221), .B2(n14236), .A(n18040), .ZN(n4282) );
  OAI21_X1 U865 ( .B1(n14218), .B2(n14236), .A(n18040), .ZN(n4279) );
  OAI21_X1 U866 ( .B1(n14215), .B2(n14236), .A(n18040), .ZN(n4275) );
  BUF_X1 U867 ( .A(n16454), .Z(n16456) );
  BUF_X1 U868 ( .A(n16454), .Z(n16457) );
  BUF_X1 U869 ( .A(n16455), .Z(n16458) );
  BUF_X1 U870 ( .A(n16707), .Z(n16709) );
  BUF_X1 U871 ( .A(n16707), .Z(n16710) );
  BUF_X1 U872 ( .A(n16708), .Z(n16711) );
  BUF_X1 U873 ( .A(n16716), .Z(n16718) );
  BUF_X1 U874 ( .A(n16716), .Z(n16719) );
  BUF_X1 U875 ( .A(n16717), .Z(n16720) );
  BUF_X1 U876 ( .A(n12565), .Z(n16355) );
  BUF_X1 U877 ( .A(n12565), .Z(n16356) );
  BUF_X1 U878 ( .A(n10571), .Z(n16607) );
  BUF_X1 U879 ( .A(n10571), .Z(n16608) );
  BUF_X1 U880 ( .A(n12615), .Z(n16259) );
  BUF_X1 U881 ( .A(n12615), .Z(n16260) );
  BUF_X1 U882 ( .A(n10635), .Z(n16511) );
  BUF_X1 U883 ( .A(n10635), .Z(n16512) );
  BUF_X1 U884 ( .A(n12564), .Z(n16358) );
  BUF_X1 U885 ( .A(n12564), .Z(n16359) );
  BUF_X1 U886 ( .A(n10569), .Z(n16610) );
  BUF_X1 U887 ( .A(n10569), .Z(n16611) );
  BUF_X1 U888 ( .A(n4182), .Z(n17720) );
  BUF_X1 U889 ( .A(n4226), .Z(n17660) );
  BUF_X1 U890 ( .A(n4117), .Z(n17804) );
  BUF_X1 U891 ( .A(n12622), .Z(n16241) );
  BUF_X1 U892 ( .A(n12622), .Z(n16242) );
  BUF_X1 U893 ( .A(n10646), .Z(n16493) );
  BUF_X1 U894 ( .A(n10646), .Z(n16494) );
  BUF_X1 U895 ( .A(n4152), .Z(n17758) );
  BUF_X1 U896 ( .A(n4152), .Z(n17757) );
  BUF_X1 U897 ( .A(n12581), .Z(n16316) );
  BUF_X1 U898 ( .A(n12571), .Z(n16340) );
  BUF_X1 U899 ( .A(n12552), .Z(n16376) );
  BUF_X1 U900 ( .A(n12556), .Z(n16367) );
  BUF_X1 U901 ( .A(n12607), .Z(n16268) );
  BUF_X1 U902 ( .A(n12590), .Z(n16304) );
  BUF_X1 U903 ( .A(n12601), .Z(n16280) );
  BUF_X1 U904 ( .A(n12632), .Z(n16217) );
  BUF_X1 U905 ( .A(n12627), .Z(n16229) );
  BUF_X1 U906 ( .A(n12581), .Z(n16317) );
  BUF_X1 U907 ( .A(n12571), .Z(n16341) );
  BUF_X1 U908 ( .A(n12552), .Z(n16377) );
  BUF_X1 U909 ( .A(n12556), .Z(n16368) );
  BUF_X1 U910 ( .A(n12607), .Z(n16269) );
  BUF_X1 U911 ( .A(n12590), .Z(n16305) );
  BUF_X1 U912 ( .A(n12601), .Z(n16281) );
  BUF_X1 U913 ( .A(n12632), .Z(n16218) );
  BUF_X1 U914 ( .A(n12627), .Z(n16230) );
  BUF_X1 U915 ( .A(n10587), .Z(n16580) );
  BUF_X1 U916 ( .A(n10580), .Z(n16592) );
  BUF_X1 U917 ( .A(n10554), .Z(n16628) );
  BUF_X1 U918 ( .A(n10560), .Z(n16619) );
  BUF_X1 U919 ( .A(n10619), .Z(n16532) );
  BUF_X1 U920 ( .A(n10626), .Z(n16520) );
  BUF_X1 U921 ( .A(n10605), .Z(n16556) );
  BUF_X1 U922 ( .A(n10660), .Z(n16469) );
  BUF_X1 U923 ( .A(n10653), .Z(n16481) );
  BUF_X1 U924 ( .A(n10587), .Z(n16581) );
  BUF_X1 U925 ( .A(n10580), .Z(n16593) );
  BUF_X1 U926 ( .A(n10554), .Z(n16629) );
  BUF_X1 U927 ( .A(n10560), .Z(n16620) );
  BUF_X1 U928 ( .A(n10619), .Z(n16533) );
  BUF_X1 U929 ( .A(n10626), .Z(n16521) );
  BUF_X1 U930 ( .A(n10605), .Z(n16557) );
  BUF_X1 U931 ( .A(n10660), .Z(n16470) );
  BUF_X1 U932 ( .A(n10653), .Z(n16482) );
  BUF_X1 U933 ( .A(n4192), .Z(n17701) );
  BUF_X1 U934 ( .A(n4192), .Z(n17700) );
  BUF_X1 U935 ( .A(n4108), .Z(n17816) );
  BUF_X1 U936 ( .A(n12562), .Z(n16363) );
  BUF_X1 U937 ( .A(n12573), .Z(n16336) );
  BUF_X1 U938 ( .A(n12568), .Z(n16348) );
  BUF_X1 U939 ( .A(n12538), .Z(n16408) );
  BUF_X1 U940 ( .A(n12548), .Z(n16384) );
  BUF_X1 U941 ( .A(n12604), .Z(n16276) );
  BUF_X1 U942 ( .A(n12587), .Z(n16312) );
  BUF_X1 U943 ( .A(n12592), .Z(n16300) );
  BUF_X1 U944 ( .A(n12597), .Z(n16288) );
  BUF_X1 U945 ( .A(n12613), .Z(n16264) );
  BUF_X1 U946 ( .A(n12629), .Z(n16225) );
  BUF_X1 U947 ( .A(n10567), .Z(n16615) );
  BUF_X1 U948 ( .A(n10583), .Z(n16588) );
  BUF_X1 U949 ( .A(n10576), .Z(n16600) );
  BUF_X1 U950 ( .A(n10550), .Z(n16636) );
  BUF_X1 U951 ( .A(n10543), .Z(n16648) );
  BUF_X1 U952 ( .A(n10615), .Z(n16540) );
  BUF_X1 U953 ( .A(n10622), .Z(n16528) );
  BUF_X1 U954 ( .A(n10601), .Z(n16564) );
  BUF_X1 U955 ( .A(n10608), .Z(n16552) );
  BUF_X1 U956 ( .A(n10633), .Z(n16516) );
  BUF_X1 U957 ( .A(n10656), .Z(n16477) );
  BUF_X1 U958 ( .A(n4162), .Z(n17744) );
  BUF_X1 U959 ( .A(n12572), .Z(n16337) );
  BUF_X1 U960 ( .A(n12577), .Z(n16325) );
  BUF_X1 U961 ( .A(n12567), .Z(n16349) );
  BUF_X1 U962 ( .A(n12542), .Z(n16397) );
  BUF_X1 U963 ( .A(n12603), .Z(n16277) );
  BUF_X1 U964 ( .A(n12591), .Z(n16301) );
  BUF_X1 U965 ( .A(n12596), .Z(n16289) );
  BUF_X1 U966 ( .A(n12612), .Z(n16265) );
  BUF_X1 U967 ( .A(n12618), .Z(n16250) );
  BUF_X1 U968 ( .A(n12623), .Z(n16238) );
  BUF_X1 U969 ( .A(n12572), .Z(n16338) );
  BUF_X1 U970 ( .A(n12577), .Z(n16326) );
  BUF_X1 U971 ( .A(n12567), .Z(n16350) );
  BUF_X1 U972 ( .A(n12542), .Z(n16398) );
  BUF_X1 U973 ( .A(n12603), .Z(n16278) );
  BUF_X1 U974 ( .A(n12591), .Z(n16302) );
  BUF_X1 U975 ( .A(n12596), .Z(n16290) );
  BUF_X1 U976 ( .A(n12612), .Z(n16266) );
  BUF_X1 U977 ( .A(n12618), .Z(n16251) );
  BUF_X1 U978 ( .A(n12623), .Z(n16239) );
  BUF_X1 U979 ( .A(n10582), .Z(n16589) );
  BUF_X1 U980 ( .A(n10589), .Z(n16577) );
  BUF_X1 U981 ( .A(n10575), .Z(n16601) );
  BUF_X1 U982 ( .A(n10542), .Z(n16649) );
  BUF_X1 U983 ( .A(n10614), .Z(n16541) );
  BUF_X1 U984 ( .A(n10621), .Z(n16529) );
  BUF_X1 U985 ( .A(n10607), .Z(n16553) );
  BUF_X1 U986 ( .A(n10632), .Z(n16517) );
  BUF_X1 U987 ( .A(n10641), .Z(n16502) );
  BUF_X1 U988 ( .A(n10648), .Z(n16490) );
  BUF_X1 U989 ( .A(n10582), .Z(n16590) );
  BUF_X1 U990 ( .A(n10589), .Z(n16578) );
  BUF_X1 U991 ( .A(n10575), .Z(n16602) );
  BUF_X1 U992 ( .A(n10542), .Z(n16650) );
  BUF_X1 U993 ( .A(n10614), .Z(n16542) );
  BUF_X1 U994 ( .A(n10621), .Z(n16530) );
  BUF_X1 U995 ( .A(n10607), .Z(n16554) );
  BUF_X1 U996 ( .A(n10632), .Z(n16518) );
  BUF_X1 U997 ( .A(n10641), .Z(n16503) );
  BUF_X1 U998 ( .A(n10648), .Z(n16491) );
  BUF_X1 U999 ( .A(n12575), .Z(n16331) );
  BUF_X1 U1000 ( .A(n12550), .Z(n16379) );
  BUF_X1 U1001 ( .A(n12606), .Z(n16271) );
  BUF_X1 U1002 ( .A(n12621), .Z(n16244) );
  BUF_X1 U1003 ( .A(n12575), .Z(n16332) );
  BUF_X1 U1004 ( .A(n12550), .Z(n16380) );
  BUF_X1 U1005 ( .A(n12606), .Z(n16272) );
  BUF_X1 U1006 ( .A(n12621), .Z(n16245) );
  BUF_X1 U1007 ( .A(n10592), .Z(n16571) );
  BUF_X1 U1008 ( .A(n10624), .Z(n16523) );
  BUF_X1 U1009 ( .A(n10644), .Z(n16496) );
  BUF_X1 U1010 ( .A(n10592), .Z(n16572) );
  BUF_X1 U1011 ( .A(n10624), .Z(n16524) );
  BUF_X1 U1012 ( .A(n10644), .Z(n16497) );
  BUF_X1 U1013 ( .A(n12580), .Z(n16319) );
  BUF_X1 U1014 ( .A(n12545), .Z(n16391) );
  BUF_X1 U1015 ( .A(n12555), .Z(n16370) );
  BUF_X1 U1016 ( .A(n12589), .Z(n16307) );
  BUF_X1 U1017 ( .A(n12631), .Z(n16220) );
  BUF_X1 U1018 ( .A(n12580), .Z(n16320) );
  BUF_X1 U1019 ( .A(n12545), .Z(n16392) );
  BUF_X1 U1020 ( .A(n12555), .Z(n16371) );
  BUF_X1 U1021 ( .A(n12589), .Z(n16308) );
  BUF_X1 U1022 ( .A(n12631), .Z(n16221) );
  BUF_X1 U1023 ( .A(n10585), .Z(n16583) );
  BUF_X1 U1024 ( .A(n10552), .Z(n16631) );
  BUF_X1 U1025 ( .A(n10558), .Z(n16622) );
  BUF_X1 U1026 ( .A(n10617), .Z(n16535) );
  BUF_X1 U1027 ( .A(n10603), .Z(n16559) );
  BUF_X1 U1028 ( .A(n10658), .Z(n16472) );
  BUF_X1 U1029 ( .A(n10585), .Z(n16584) );
  BUF_X1 U1030 ( .A(n10552), .Z(n16632) );
  BUF_X1 U1031 ( .A(n10558), .Z(n16623) );
  BUF_X1 U1032 ( .A(n10617), .Z(n16536) );
  BUF_X1 U1033 ( .A(n10603), .Z(n16560) );
  BUF_X1 U1034 ( .A(n10658), .Z(n16473) );
  BUF_X1 U1035 ( .A(n12570), .Z(n16343) );
  BUF_X1 U1036 ( .A(n12594), .Z(n16295) );
  BUF_X1 U1037 ( .A(n12599), .Z(n16283) );
  BUF_X1 U1038 ( .A(n12626), .Z(n16232) );
  BUF_X1 U1039 ( .A(n12570), .Z(n16344) );
  BUF_X1 U1040 ( .A(n12594), .Z(n16296) );
  BUF_X1 U1041 ( .A(n12599), .Z(n16284) );
  BUF_X1 U1042 ( .A(n12626), .Z(n16233) );
  BUF_X1 U1043 ( .A(n10578), .Z(n16595) );
  BUF_X1 U1044 ( .A(n10545), .Z(n16643) );
  BUF_X1 U1045 ( .A(n10610), .Z(n16547) );
  BUF_X1 U1046 ( .A(n10651), .Z(n16484) );
  BUF_X1 U1047 ( .A(n10578), .Z(n16596) );
  BUF_X1 U1048 ( .A(n10545), .Z(n16644) );
  BUF_X1 U1049 ( .A(n10610), .Z(n16548) );
  BUF_X1 U1050 ( .A(n10651), .Z(n16485) );
  BUF_X1 U1051 ( .A(n4164), .Z(n17740) );
  BUF_X1 U1052 ( .A(n4164), .Z(n17739) );
  BUF_X1 U1053 ( .A(n12617), .Z(n16255) );
  BUF_X1 U1054 ( .A(n10639), .Z(n16507) );
  BUF_X1 U1055 ( .A(n12565), .Z(n16357) );
  BUF_X1 U1056 ( .A(n10571), .Z(n16609) );
  BUF_X1 U1057 ( .A(n12615), .Z(n16261) );
  BUF_X1 U1058 ( .A(n10635), .Z(n16513) );
  BUF_X1 U1059 ( .A(n12564), .Z(n16360) );
  BUF_X1 U1060 ( .A(n10569), .Z(n16612) );
  BUF_X1 U1061 ( .A(n4152), .Z(n17759) );
  BUF_X1 U1062 ( .A(n12622), .Z(n16243) );
  BUF_X1 U1063 ( .A(n10646), .Z(n16495) );
  BUF_X1 U1064 ( .A(n12607), .Z(n16270) );
  BUF_X1 U1065 ( .A(n12581), .Z(n16318) );
  BUF_X1 U1066 ( .A(n12571), .Z(n16342) );
  BUF_X1 U1067 ( .A(n12552), .Z(n16378) );
  BUF_X1 U1068 ( .A(n12556), .Z(n16369) );
  BUF_X1 U1069 ( .A(n12590), .Z(n16306) );
  BUF_X1 U1070 ( .A(n12601), .Z(n16282) );
  BUF_X1 U1071 ( .A(n12632), .Z(n16219) );
  BUF_X1 U1072 ( .A(n12627), .Z(n16231) );
  BUF_X1 U1073 ( .A(n10587), .Z(n16582) );
  BUF_X1 U1074 ( .A(n10626), .Z(n16522) );
  BUF_X1 U1075 ( .A(n10580), .Z(n16594) );
  BUF_X1 U1076 ( .A(n10554), .Z(n16630) );
  BUF_X1 U1077 ( .A(n10560), .Z(n16621) );
  BUF_X1 U1078 ( .A(n10619), .Z(n16534) );
  BUF_X1 U1079 ( .A(n10605), .Z(n16558) );
  BUF_X1 U1080 ( .A(n10660), .Z(n16471) );
  BUF_X1 U1081 ( .A(n10653), .Z(n16483) );
  BUF_X1 U1082 ( .A(n4192), .Z(n17702) );
  BUF_X1 U1083 ( .A(n12575), .Z(n16333) );
  BUF_X1 U1084 ( .A(n12550), .Z(n16381) );
  BUF_X1 U1085 ( .A(n12606), .Z(n16273) );
  BUF_X1 U1086 ( .A(n12621), .Z(n16246) );
  BUF_X1 U1087 ( .A(n10592), .Z(n16573) );
  BUF_X1 U1088 ( .A(n10624), .Z(n16525) );
  BUF_X1 U1089 ( .A(n10644), .Z(n16498) );
  BUF_X1 U1090 ( .A(n12572), .Z(n16339) );
  BUF_X1 U1091 ( .A(n12577), .Z(n16327) );
  BUF_X1 U1092 ( .A(n12567), .Z(n16351) );
  BUF_X1 U1093 ( .A(n12542), .Z(n16399) );
  BUF_X1 U1094 ( .A(n12603), .Z(n16279) );
  BUF_X1 U1095 ( .A(n12591), .Z(n16303) );
  BUF_X1 U1096 ( .A(n12596), .Z(n16291) );
  BUF_X1 U1097 ( .A(n12612), .Z(n16267) );
  BUF_X1 U1098 ( .A(n12618), .Z(n16252) );
  BUF_X1 U1099 ( .A(n12623), .Z(n16240) );
  BUF_X1 U1100 ( .A(n10582), .Z(n16591) );
  BUF_X1 U1101 ( .A(n10589), .Z(n16579) );
  BUF_X1 U1102 ( .A(n10575), .Z(n16603) );
  BUF_X1 U1103 ( .A(n10542), .Z(n16651) );
  BUF_X1 U1104 ( .A(n10614), .Z(n16543) );
  BUF_X1 U1105 ( .A(n10621), .Z(n16531) );
  BUF_X1 U1106 ( .A(n10607), .Z(n16555) );
  BUF_X1 U1107 ( .A(n10632), .Z(n16519) );
  BUF_X1 U1108 ( .A(n10641), .Z(n16504) );
  BUF_X1 U1109 ( .A(n10648), .Z(n16492) );
  BUF_X1 U1110 ( .A(n10585), .Z(n16585) );
  BUF_X1 U1111 ( .A(n10552), .Z(n16633) );
  BUF_X1 U1112 ( .A(n10558), .Z(n16624) );
  BUF_X1 U1113 ( .A(n10617), .Z(n16537) );
  BUF_X1 U1114 ( .A(n10603), .Z(n16561) );
  BUF_X1 U1115 ( .A(n10658), .Z(n16474) );
  BUF_X1 U1116 ( .A(n12580), .Z(n16321) );
  BUF_X1 U1117 ( .A(n12545), .Z(n16393) );
  BUF_X1 U1118 ( .A(n12555), .Z(n16372) );
  BUF_X1 U1119 ( .A(n12589), .Z(n16309) );
  BUF_X1 U1120 ( .A(n12631), .Z(n16222) );
  BUF_X1 U1121 ( .A(n12570), .Z(n16345) );
  BUF_X1 U1122 ( .A(n12594), .Z(n16297) );
  BUF_X1 U1123 ( .A(n12599), .Z(n16285) );
  BUF_X1 U1124 ( .A(n12626), .Z(n16234) );
  BUF_X1 U1125 ( .A(n10578), .Z(n16597) );
  BUF_X1 U1126 ( .A(n10545), .Z(n16645) );
  BUF_X1 U1127 ( .A(n10610), .Z(n16549) );
  BUF_X1 U1128 ( .A(n10651), .Z(n16486) );
  BUF_X1 U1129 ( .A(n4164), .Z(n17741) );
  OAI21_X1 U1130 ( .B1(n14061), .B2(n14062), .A(n18039), .ZN(n4067) );
  OAI21_X1 U1131 ( .B1(n14063), .B2(n14237), .A(n18041), .ZN(n4309) );
  OAI21_X1 U1132 ( .B1(n14062), .B2(n14237), .A(n18041), .ZN(n4306) );
  BUF_X1 U1133 ( .A(n18054), .Z(n18052) );
  BUF_X1 U1134 ( .A(n18054), .Z(n18051) );
  NAND2_X1 U1135 ( .A1(n14258), .A2(n14249), .ZN(n14073) );
  NAND2_X1 U1136 ( .A1(n14258), .A2(n14251), .ZN(n14074) );
  BUF_X1 U1137 ( .A(n17822), .Z(n17834) );
  AND2_X1 U1138 ( .A1(n12489), .A2(n12437), .ZN(n12440) );
  BUF_X1 U1139 ( .A(n16688), .Z(n16695) );
  BUF_X1 U1140 ( .A(n16688), .Z(n16694) );
  BUF_X1 U1141 ( .A(n17573), .Z(n17580) );
  BUF_X1 U1142 ( .A(n17573), .Z(n17579) );
  BUF_X1 U1143 ( .A(n18055), .Z(n18050) );
  BUF_X1 U1144 ( .A(n18054), .Z(n18053) );
  NAND2_X1 U1145 ( .A1(n14085), .A2(n14086), .ZN(n4112) );
  NAND2_X1 U1146 ( .A1(n14085), .A2(n14088), .ZN(n4121) );
  NAND2_X1 U1147 ( .A1(n14085), .A2(n14103), .ZN(n4128) );
  BUF_X1 U1148 ( .A(n16689), .Z(n16696) );
  BUF_X1 U1149 ( .A(n17574), .Z(n17581) );
  NAND2_X1 U1150 ( .A1(n13919), .A2(n13920), .ZN(n12540) );
  NAND2_X1 U1151 ( .A1(n13925), .A2(n13920), .ZN(n12546) );
  NAND2_X1 U1152 ( .A1(n12438), .A2(n12439), .ZN(n10538) );
  NAND2_X1 U1153 ( .A1(n12443), .A2(n12439), .ZN(n10547) );
  NAND2_X1 U1154 ( .A1(n14107), .A2(n14085), .ZN(n4248) );
  NAND2_X1 U1155 ( .A1(n13936), .A2(n13918), .ZN(n12566) );
  NAND2_X1 U1156 ( .A1(n13946), .A2(n13918), .ZN(n12576) );
  NAND2_X1 U1157 ( .A1(n13917), .A2(n13918), .ZN(n12541) );
  NAND2_X1 U1158 ( .A1(n13953), .A2(n13918), .ZN(n12595) );
  NAND2_X1 U1159 ( .A1(n13960), .A2(n13918), .ZN(n12616) );
  NAND2_X1 U1160 ( .A1(n12455), .A2(n12437), .ZN(n10573) );
  NAND2_X1 U1161 ( .A1(n12465), .A2(n12437), .ZN(n10594) );
  NAND2_X1 U1162 ( .A1(n12436), .A2(n12437), .ZN(n10540) );
  NAND2_X1 U1163 ( .A1(n12472), .A2(n12437), .ZN(n10612) );
  NAND2_X1 U1164 ( .A1(n12479), .A2(n12437), .ZN(n10637) );
  NAND2_X1 U1165 ( .A1(n14087), .A2(n14088), .ZN(n4110) );
  INV_X1 U1166 ( .A(n14201), .ZN(n14088) );
  AND2_X1 U1167 ( .A1(n13970), .A2(n13918), .ZN(n13928) );
  INV_X1 U1168 ( .A(n14097), .ZN(n14103) );
  BUF_X1 U1169 ( .A(n16455), .Z(n16459) );
  BUF_X1 U1170 ( .A(n16708), .Z(n16712) );
  BUF_X1 U1171 ( .A(n16717), .Z(n16721) );
  AND2_X1 U1172 ( .A1(n13926), .A2(n13918), .ZN(n12553) );
  AND2_X1 U1173 ( .A1(n13969), .A2(n13918), .ZN(n12619) );
  AND2_X1 U1174 ( .A1(n13955), .A2(n13918), .ZN(n12628) );
  AND2_X1 U1175 ( .A1(n12450), .A2(n12437), .ZN(n10556) );
  AND2_X1 U1176 ( .A1(n12488), .A2(n12437), .ZN(n10642) );
  AND2_X1 U1177 ( .A1(n12477), .A2(n12437), .ZN(n10655) );
  AND2_X1 U1178 ( .A1(n13920), .A2(n13923), .ZN(n12537) );
  AND2_X1 U1179 ( .A1(n12439), .A2(n12441), .ZN(n10535) );
  BUF_X1 U1180 ( .A(n16688), .Z(n16693) );
  BUF_X1 U1181 ( .A(n17573), .Z(n17578) );
  AND2_X1 U1182 ( .A1(n13931), .A2(n13920), .ZN(n12561) );
  AND2_X1 U1183 ( .A1(n13929), .A2(n13920), .ZN(n12578) );
  AND2_X1 U1184 ( .A1(n13928), .A2(n13920), .ZN(n12543) );
  AND2_X1 U1185 ( .A1(n13922), .A2(n13920), .ZN(n12547) );
  AND2_X1 U1186 ( .A1(n13933), .A2(n13920), .ZN(n12586) );
  AND2_X1 U1187 ( .A1(n12449), .A2(n12439), .ZN(n10566) );
  AND2_X1 U1188 ( .A1(n12447), .A2(n12439), .ZN(n10590) );
  AND2_X1 U1189 ( .A1(n12440), .A2(n12439), .ZN(n10536) );
  AND2_X1 U1190 ( .A1(n12445), .A2(n12439), .ZN(n10549) );
  AND2_X1 U1191 ( .A1(n12446), .A2(n12439), .ZN(n10600) );
  BUF_X1 U1192 ( .A(n17545), .Z(n17550) );
  BUF_X1 U1193 ( .A(n17559), .Z(n17564) );
  BUF_X1 U1194 ( .A(n17586), .Z(n17591) );
  BUF_X1 U1195 ( .A(n17600), .Z(n17605) );
  BUF_X1 U1196 ( .A(n17614), .Z(n17619) );
  BUF_X1 U1197 ( .A(n17531), .Z(n17536) );
  BUF_X1 U1198 ( .A(n17547), .Z(n17557) );
  BUF_X1 U1199 ( .A(n17561), .Z(n17571) );
  BUF_X1 U1200 ( .A(n17588), .Z(n17598) );
  BUF_X1 U1201 ( .A(n17602), .Z(n17612) );
  BUF_X1 U1202 ( .A(n17616), .Z(n17626) );
  BUF_X1 U1203 ( .A(n16689), .Z(n16698) );
  BUF_X1 U1204 ( .A(n16689), .Z(n16697) );
  BUF_X1 U1205 ( .A(n17533), .Z(n17542) );
  BUF_X1 U1206 ( .A(n17547), .Z(n17556) );
  BUF_X1 U1207 ( .A(n17561), .Z(n17570) );
  BUF_X1 U1208 ( .A(n17588), .Z(n17597) );
  BUF_X1 U1209 ( .A(n17602), .Z(n17611) );
  BUF_X1 U1210 ( .A(n17616), .Z(n17625) );
  BUF_X1 U1211 ( .A(n17532), .Z(n17541) );
  BUF_X1 U1212 ( .A(n17546), .Z(n17555) );
  BUF_X1 U1213 ( .A(n17560), .Z(n17569) );
  BUF_X1 U1214 ( .A(n17574), .Z(n17583) );
  BUF_X1 U1215 ( .A(n17587), .Z(n17596) );
  BUF_X1 U1216 ( .A(n17601), .Z(n17610) );
  BUF_X1 U1217 ( .A(n17615), .Z(n17624) );
  BUF_X1 U1218 ( .A(n17532), .Z(n17539) );
  BUF_X1 U1219 ( .A(n17546), .Z(n17553) );
  BUF_X1 U1220 ( .A(n17560), .Z(n17567) );
  BUF_X1 U1221 ( .A(n17587), .Z(n17594) );
  BUF_X1 U1222 ( .A(n17601), .Z(n17608) );
  BUF_X1 U1223 ( .A(n17615), .Z(n17622) );
  BUF_X1 U1224 ( .A(n17532), .Z(n17540) );
  BUF_X1 U1225 ( .A(n17546), .Z(n17554) );
  BUF_X1 U1226 ( .A(n17560), .Z(n17568) );
  BUF_X1 U1227 ( .A(n17574), .Z(n17582) );
  BUF_X1 U1228 ( .A(n17587), .Z(n17595) );
  BUF_X1 U1229 ( .A(n17601), .Z(n17609) );
  BUF_X1 U1230 ( .A(n17615), .Z(n17623) );
  BUF_X1 U1231 ( .A(n17531), .Z(n17538) );
  BUF_X1 U1232 ( .A(n17545), .Z(n17552) );
  BUF_X1 U1233 ( .A(n17559), .Z(n17566) );
  BUF_X1 U1234 ( .A(n17586), .Z(n17593) );
  BUF_X1 U1235 ( .A(n17600), .Z(n17607) );
  BUF_X1 U1236 ( .A(n17614), .Z(n17621) );
  BUF_X1 U1237 ( .A(n17531), .Z(n17537) );
  BUF_X1 U1238 ( .A(n17545), .Z(n17551) );
  BUF_X1 U1239 ( .A(n17559), .Z(n17565) );
  BUF_X1 U1240 ( .A(n17586), .Z(n17592) );
  BUF_X1 U1241 ( .A(n17600), .Z(n17606) );
  BUF_X1 U1242 ( .A(n17614), .Z(n17620) );
  BUF_X1 U1243 ( .A(n17533), .Z(n17543) );
  BUF_X1 U1244 ( .A(n16690), .Z(n16700) );
  BUF_X1 U1245 ( .A(n17575), .Z(n17585) );
  BUF_X1 U1246 ( .A(n16690), .Z(n16699) );
  BUF_X1 U1247 ( .A(n17575), .Z(n17584) );
  BUF_X1 U1248 ( .A(n4367), .Z(n17192) );
  OAI21_X1 U1249 ( .B1(n14063), .B2(n14244), .A(n18042), .ZN(n4367) );
  BUF_X1 U1250 ( .A(n4423), .Z(n16999) );
  OAI21_X1 U1251 ( .B1(n14063), .B2(n14252), .A(n18042), .ZN(n4423) );
  OAI21_X1 U1252 ( .B1(n14062), .B2(n14252), .A(n18043), .ZN(n4420) );
  OAI21_X1 U1253 ( .B1(n14062), .B2(n14244), .A(n18042), .ZN(n4362) );
  BUF_X1 U1254 ( .A(n17533), .Z(n17544) );
  BUF_X1 U1255 ( .A(n17547), .Z(n17558) );
  BUF_X1 U1256 ( .A(n17561), .Z(n17572) );
  BUF_X1 U1257 ( .A(n17588), .Z(n17599) );
  BUF_X1 U1258 ( .A(n17602), .Z(n17613) );
  INV_X1 U1259 ( .A(n14089), .ZN(n14086) );
  INV_X1 U1260 ( .A(n14098), .ZN(n14158) );
  BUF_X1 U1261 ( .A(n17616), .Z(n17627) );
  BUF_X1 U1262 ( .A(n4062), .Z(n18000) );
  BUF_X1 U1263 ( .A(n4456), .Z(n16897) );
  BUF_X1 U1264 ( .A(n4467), .Z(n16865) );
  BUF_X1 U1265 ( .A(n4062), .Z(n18001) );
  BUF_X1 U1266 ( .A(n4467), .Z(n16864) );
  BUF_X1 U1267 ( .A(n4456), .Z(n16898) );
  BUF_X1 U1268 ( .A(n4467), .Z(n16863) );
  BUF_X1 U1269 ( .A(n4385), .Z(n17124) );
  BUF_X1 U1270 ( .A(n4379), .Z(n17147) );
  BUF_X1 U1271 ( .A(n4359), .Z(n17213) );
  BUF_X1 U1272 ( .A(n4356), .Z(n17226) );
  BUF_X1 U1273 ( .A(n4351), .Z(n17239) );
  BUF_X1 U1274 ( .A(n4348), .Z(n17252) );
  BUF_X1 U1275 ( .A(n4341), .Z(n17265) );
  BUF_X1 U1276 ( .A(n4338), .Z(n17278) );
  BUF_X1 U1277 ( .A(n4335), .Z(n17291) );
  BUF_X1 U1278 ( .A(n4332), .Z(n17304) );
  BUF_X1 U1279 ( .A(n4385), .Z(n17125) );
  BUF_X1 U1280 ( .A(n4379), .Z(n17148) );
  BUF_X1 U1281 ( .A(n4359), .Z(n17214) );
  BUF_X1 U1282 ( .A(n4356), .Z(n17227) );
  BUF_X1 U1283 ( .A(n4351), .Z(n17240) );
  BUF_X1 U1284 ( .A(n4348), .Z(n17253) );
  BUF_X1 U1285 ( .A(n4341), .Z(n17266) );
  BUF_X1 U1286 ( .A(n4338), .Z(n17279) );
  BUF_X1 U1287 ( .A(n4335), .Z(n17292) );
  BUF_X1 U1288 ( .A(n4332), .Z(n17305) );
  BUF_X1 U1289 ( .A(n4441), .Z(n16931) );
  BUF_X1 U1290 ( .A(n4417), .Z(n17020) );
  BUF_X1 U1291 ( .A(n4412), .Z(n17033) );
  BUF_X1 U1292 ( .A(n4409), .Z(n17046) );
  BUF_X1 U1293 ( .A(n4406), .Z(n17059) );
  BUF_X1 U1294 ( .A(n4401), .Z(n17072) );
  BUF_X1 U1295 ( .A(n4398), .Z(n17085) );
  BUF_X1 U1296 ( .A(n4391), .Z(n17098) );
  BUF_X1 U1297 ( .A(n4388), .Z(n17111) );
  BUF_X1 U1298 ( .A(n4441), .Z(n16932) );
  BUF_X1 U1299 ( .A(n4417), .Z(n17021) );
  BUF_X1 U1300 ( .A(n4412), .Z(n17034) );
  BUF_X1 U1301 ( .A(n4409), .Z(n17047) );
  BUF_X1 U1302 ( .A(n4406), .Z(n17060) );
  BUF_X1 U1303 ( .A(n4401), .Z(n17073) );
  BUF_X1 U1304 ( .A(n4398), .Z(n17086) );
  BUF_X1 U1305 ( .A(n4391), .Z(n17099) );
  BUF_X1 U1306 ( .A(n4388), .Z(n17112) );
  BUF_X1 U1307 ( .A(n4059), .Z(n18013) );
  BUF_X1 U1308 ( .A(n4059), .Z(n18014) );
  BUF_X1 U1309 ( .A(n4317), .Z(n17369) );
  BUF_X1 U1310 ( .A(n4317), .Z(n17370) );
  BUF_X1 U1311 ( .A(n4426), .Z(n16986) );
  BUF_X1 U1312 ( .A(n4312), .Z(n17382) );
  BUF_X1 U1313 ( .A(n4426), .Z(n16987) );
  BUF_X1 U1314 ( .A(n4312), .Z(n17383) );
  BUF_X1 U1315 ( .A(n4062), .Z(n18002) );
  BUF_X1 U1316 ( .A(n4456), .Z(n16899) );
  BUF_X1 U1317 ( .A(n4385), .Z(n17126) );
  BUF_X1 U1318 ( .A(n4379), .Z(n17149) );
  BUF_X1 U1319 ( .A(n4359), .Z(n17215) );
  BUF_X1 U1320 ( .A(n4356), .Z(n17228) );
  BUF_X1 U1321 ( .A(n4351), .Z(n17241) );
  BUF_X1 U1322 ( .A(n4348), .Z(n17254) );
  BUF_X1 U1323 ( .A(n4341), .Z(n17267) );
  BUF_X1 U1324 ( .A(n4338), .Z(n17280) );
  BUF_X1 U1325 ( .A(n4335), .Z(n17293) );
  BUF_X1 U1326 ( .A(n4332), .Z(n17306) );
  BUF_X1 U1327 ( .A(n4441), .Z(n16933) );
  BUF_X1 U1328 ( .A(n4417), .Z(n17022) );
  BUF_X1 U1329 ( .A(n4412), .Z(n17035) );
  BUF_X1 U1330 ( .A(n4409), .Z(n17048) );
  BUF_X1 U1331 ( .A(n4406), .Z(n17061) );
  BUF_X1 U1332 ( .A(n4401), .Z(n17074) );
  BUF_X1 U1333 ( .A(n4398), .Z(n17087) );
  BUF_X1 U1334 ( .A(n4391), .Z(n17100) );
  BUF_X1 U1335 ( .A(n4388), .Z(n17113) );
  BUF_X1 U1336 ( .A(n4059), .Z(n18015) );
  BUF_X1 U1337 ( .A(n4317), .Z(n17371) );
  BUF_X1 U1338 ( .A(n4426), .Z(n16988) );
  BUF_X1 U1339 ( .A(n4312), .Z(n17384) );
  INV_X1 U1340 ( .A(n16944), .ZN(n16955) );
  INV_X1 U1341 ( .A(n16956), .ZN(n16965) );
  INV_X1 U1342 ( .A(n16966), .ZN(n16975) );
  INV_X1 U1343 ( .A(n17137), .ZN(n17146) );
  INV_X1 U1344 ( .A(n17160), .ZN(n17169) );
  INV_X1 U1345 ( .A(n16877), .ZN(n16886) );
  INV_X1 U1346 ( .A(n16887), .ZN(n16896) );
  INV_X1 U1347 ( .A(n16910), .ZN(n16919) );
  INV_X1 U1348 ( .A(n4448), .ZN(n16930) );
  INV_X1 U1349 ( .A(n16976), .ZN(n16985) );
  INV_X1 U1350 ( .A(n17170), .ZN(n17181) );
  INV_X1 U1351 ( .A(n17182), .ZN(n17191) );
  BUF_X1 U1352 ( .A(n18055), .Z(n18048) );
  BUF_X1 U1353 ( .A(n18048), .Z(n18047) );
  BUF_X1 U1354 ( .A(n18049), .Z(n18046) );
  BUF_X1 U1355 ( .A(n18049), .Z(n18045) );
  BUF_X1 U1356 ( .A(n18055), .Z(n18049) );
  BUF_X1 U1357 ( .A(n17822), .Z(n17832) );
  BUF_X1 U1358 ( .A(n17821), .Z(n17831) );
  BUF_X1 U1359 ( .A(n17821), .Z(n17830) );
  BUF_X1 U1360 ( .A(n17821), .Z(n17829) );
  BUF_X1 U1361 ( .A(n17820), .Z(n17828) );
  BUF_X1 U1362 ( .A(n17820), .Z(n17827) );
  BUF_X1 U1363 ( .A(n17820), .Z(n17826) );
  BUF_X1 U1364 ( .A(n17822), .Z(n17833) );
  NAND3_X1 U1365 ( .A1(n14239), .A2(n14234), .A3(n14240), .ZN(n14236) );
  OAI22_X1 U1366 ( .A1(n14022), .A2(n14136), .B1(n14096), .B2(n14134), .ZN(
        n4152) );
  OAI22_X1 U1367 ( .A1(n14166), .A2(n14124), .B1(n14167), .B2(n14125), .ZN(
        n4226) );
  OAI22_X1 U1368 ( .A1(n14120), .A2(n14124), .B1(n14121), .B2(n14125), .ZN(
        n4182) );
  OAI21_X1 U1369 ( .B1(n14066), .B2(n14061), .A(n18040), .ZN(n4076) );
  OAI21_X1 U1370 ( .B1(n14064), .B2(n14061), .A(n18039), .ZN(n4073) );
  NOR2_X1 U1371 ( .A1(n14257), .A2(n14259), .ZN(n14258) );
  NOR2_X1 U1372 ( .A1(n14096), .A2(n14097), .ZN(n4117) );
  BUF_X1 U1373 ( .A(n12624), .Z(n16235) );
  BUF_X1 U1374 ( .A(n12624), .Z(n16236) );
  INV_X1 U1375 ( .A(n14099), .ZN(n14085) );
  AND3_X1 U1376 ( .A1(n13980), .A2(n13963), .A3(n13962), .ZN(n13920) );
  AND3_X1 U1377 ( .A1(n12499), .A2(n12482), .A3(n12481), .ZN(n12439) );
  INV_X1 U1378 ( .A(n14162), .ZN(n4192) );
  OAI22_X1 U1379 ( .A1(n14163), .A2(n14124), .B1(n14164), .B2(n14125), .ZN(
        n14162) );
  OAI21_X1 U1380 ( .B1(n14059), .B2(n14228), .A(n18041), .ZN(n4467) );
  OAI21_X1 U1381 ( .B1(n14059), .B2(n12414), .A(n18039), .ZN(n4062) );
  OAI21_X1 U1382 ( .B1(n14059), .B2(n14221), .A(n18044), .ZN(n4456) );
  BUF_X1 U1383 ( .A(n10523), .Z(n16670) );
  BUF_X1 U1384 ( .A(n10517), .Z(n16682) );
  BUF_X1 U1385 ( .A(n10662), .Z(n16466) );
  BUF_X1 U1386 ( .A(n10649), .Z(n16487) );
  BUF_X1 U1387 ( .A(n4153), .Z(n17755) );
  BUF_X1 U1388 ( .A(n4153), .Z(n17754) );
  BUF_X1 U1389 ( .A(n4198), .Z(n17695) );
  BUF_X1 U1390 ( .A(n4198), .Z(n17694) );
  BUF_X1 U1391 ( .A(n4233), .Z(n17647) );
  BUF_X1 U1392 ( .A(n4233), .Z(n17646) );
  BUF_X1 U1393 ( .A(n4207), .Z(n17683) );
  BUF_X1 U1394 ( .A(n4207), .Z(n17682) );
  BUF_X1 U1395 ( .A(n4220), .Z(n17671) );
  BUF_X1 U1396 ( .A(n4220), .Z(n17670) );
  BUF_X1 U1397 ( .A(n4142), .Z(n17767) );
  BUF_X1 U1398 ( .A(n4189), .Z(n17707) );
  BUF_X1 U1399 ( .A(n4142), .Z(n17766) );
  BUF_X1 U1400 ( .A(n4189), .Z(n17706) );
  BUF_X1 U1401 ( .A(n4171), .Z(n17731) );
  BUF_X1 U1402 ( .A(n4124), .Z(n17791) );
  BUF_X1 U1403 ( .A(n4131), .Z(n17779) );
  BUF_X1 U1404 ( .A(n4171), .Z(n17730) );
  BUF_X1 U1405 ( .A(n4124), .Z(n17790) );
  BUF_X1 U1406 ( .A(n4131), .Z(n17778) );
  BUF_X1 U1407 ( .A(n10663), .Z(n16463) );
  BUF_X1 U1408 ( .A(n10649), .Z(n16488) );
  BUF_X1 U1409 ( .A(n10519), .Z(n16679) );
  BUF_X1 U1410 ( .A(n10662), .Z(n16467) );
  BUF_X1 U1411 ( .A(n10523), .Z(n16671) );
  BUF_X1 U1412 ( .A(n10517), .Z(n16683) );
  NOR2_X1 U1413 ( .A1(n14089), .A2(n14090), .ZN(n4108) );
  BUF_X1 U1414 ( .A(n10519), .Z(n16680) );
  BUF_X1 U1415 ( .A(n4058), .Z(n18026) );
  BUF_X1 U1416 ( .A(n4058), .Z(n18030) );
  BUF_X1 U1417 ( .A(n4058), .Z(n18029) );
  BUF_X1 U1418 ( .A(n4058), .Z(n18028) );
  BUF_X1 U1419 ( .A(n4058), .Z(n18027) );
  BUF_X1 U1420 ( .A(n10510), .Z(n16701) );
  INV_X1 U1421 ( .A(n14034), .ZN(n14033) );
  BUF_X1 U1422 ( .A(n4058), .Z(n18031) );
  BUF_X1 U1423 ( .A(n12522), .Z(n16427) );
  BUF_X1 U1424 ( .A(n12522), .Z(n16428) );
  BUF_X1 U1425 ( .A(n10510), .Z(n16702) );
  OAI21_X1 U1426 ( .B1(n14074), .B2(n14241), .A(n18042), .ZN(n4385) );
  OAI21_X1 U1427 ( .B1(n14072), .B2(n14241), .A(n18042), .ZN(n4379) );
  OAI21_X1 U1428 ( .B1(n12414), .B2(n14241), .A(n18042), .ZN(n4359) );
  OAI21_X1 U1429 ( .B1(n14058), .B2(n14241), .A(n18041), .ZN(n4356) );
  OAI21_X1 U1430 ( .B1(n14228), .B2(n14241), .A(n18042), .ZN(n4351) );
  OAI21_X1 U1431 ( .B1(n14226), .B2(n14241), .A(n18041), .ZN(n4348) );
  OAI21_X1 U1432 ( .B1(n14222), .B2(n14241), .A(n18039), .ZN(n4341) );
  OAI21_X1 U1433 ( .B1(n14221), .B2(n14241), .A(n18041), .ZN(n4338) );
  OAI21_X1 U1434 ( .B1(n14218), .B2(n14241), .A(n18041), .ZN(n4335) );
  OAI21_X1 U1435 ( .B1(n14215), .B2(n14241), .A(n18041), .ZN(n4332) );
  BUF_X1 U1436 ( .A(n7537), .Z(n16731) );
  BUF_X1 U1437 ( .A(n7537), .Z(n16732) );
  BUF_X1 U1438 ( .A(n7537), .Z(n16733) );
  BUF_X1 U1439 ( .A(n7537), .Z(n16734) );
  BUF_X1 U1440 ( .A(n7537), .Z(n16735) );
  BUF_X1 U1441 ( .A(n7537), .Z(n16736) );
  BUF_X1 U1442 ( .A(n7428), .Z(n16737) );
  BUF_X1 U1443 ( .A(n7428), .Z(n16738) );
  BUF_X1 U1444 ( .A(n7428), .Z(n16739) );
  BUF_X1 U1445 ( .A(n7428), .Z(n16740) );
  BUF_X1 U1446 ( .A(n7428), .Z(n16741) );
  BUF_X1 U1447 ( .A(n7428), .Z(n16742) );
  BUF_X1 U1448 ( .A(n7319), .Z(n16743) );
  BUF_X1 U1449 ( .A(n7319), .Z(n16744) );
  BUF_X1 U1450 ( .A(n7319), .Z(n16745) );
  BUF_X1 U1451 ( .A(n7319), .Z(n16746) );
  BUF_X1 U1452 ( .A(n7319), .Z(n16747) );
  BUF_X1 U1453 ( .A(n7319), .Z(n16748) );
  BUF_X1 U1454 ( .A(n7205), .Z(n16749) );
  BUF_X1 U1455 ( .A(n7205), .Z(n16750) );
  BUF_X1 U1456 ( .A(n7205), .Z(n16751) );
  BUF_X1 U1457 ( .A(n7205), .Z(n16752) );
  BUF_X1 U1458 ( .A(n7205), .Z(n16753) );
  BUF_X1 U1459 ( .A(n7205), .Z(n16754) );
  BUF_X1 U1460 ( .A(n7096), .Z(n16755) );
  BUF_X1 U1461 ( .A(n7096), .Z(n16756) );
  BUF_X1 U1462 ( .A(n7096), .Z(n16757) );
  BUF_X1 U1463 ( .A(n7096), .Z(n16758) );
  BUF_X1 U1464 ( .A(n7096), .Z(n16759) );
  BUF_X1 U1465 ( .A(n7096), .Z(n16760) );
  BUF_X1 U1466 ( .A(n6987), .Z(n16761) );
  BUF_X1 U1467 ( .A(n6987), .Z(n16762) );
  BUF_X1 U1468 ( .A(n6987), .Z(n16763) );
  BUF_X1 U1469 ( .A(n6987), .Z(n16764) );
  BUF_X1 U1470 ( .A(n6987), .Z(n16765) );
  BUF_X1 U1471 ( .A(n6987), .Z(n16766) );
  BUF_X1 U1472 ( .A(n6878), .Z(n16767) );
  BUF_X1 U1473 ( .A(n6878), .Z(n16768) );
  BUF_X1 U1474 ( .A(n6878), .Z(n16769) );
  BUF_X1 U1475 ( .A(n6878), .Z(n16770) );
  BUF_X1 U1476 ( .A(n6878), .Z(n16771) );
  BUF_X1 U1477 ( .A(n6878), .Z(n16772) );
  BUF_X1 U1478 ( .A(n6769), .Z(n16773) );
  BUF_X1 U1479 ( .A(n6769), .Z(n16774) );
  BUF_X1 U1480 ( .A(n6769), .Z(n16775) );
  BUF_X1 U1481 ( .A(n6769), .Z(n16776) );
  BUF_X1 U1482 ( .A(n6769), .Z(n16777) );
  BUF_X1 U1483 ( .A(n6769), .Z(n16778) );
  BUF_X1 U1484 ( .A(n6635), .Z(n16779) );
  BUF_X1 U1485 ( .A(n6635), .Z(n16780) );
  BUF_X1 U1486 ( .A(n6635), .Z(n16781) );
  BUF_X1 U1487 ( .A(n6635), .Z(n16782) );
  BUF_X1 U1488 ( .A(n6635), .Z(n16783) );
  BUF_X1 U1489 ( .A(n6635), .Z(n16784) );
  BUF_X1 U1490 ( .A(n6448), .Z(n16785) );
  BUF_X1 U1491 ( .A(n6448), .Z(n16786) );
  BUF_X1 U1492 ( .A(n6448), .Z(n16787) );
  BUF_X1 U1493 ( .A(n6448), .Z(n16788) );
  BUF_X1 U1494 ( .A(n6448), .Z(n16789) );
  BUF_X1 U1495 ( .A(n6448), .Z(n16790) );
  BUF_X1 U1496 ( .A(n6261), .Z(n16791) );
  BUF_X1 U1497 ( .A(n6261), .Z(n16792) );
  BUF_X1 U1498 ( .A(n6261), .Z(n16793) );
  BUF_X1 U1499 ( .A(n6261), .Z(n16794) );
  BUF_X1 U1500 ( .A(n6261), .Z(n16795) );
  BUF_X1 U1501 ( .A(n6261), .Z(n16796) );
  BUF_X1 U1502 ( .A(n6076), .Z(n16797) );
  BUF_X1 U1503 ( .A(n6076), .Z(n16798) );
  BUF_X1 U1504 ( .A(n6076), .Z(n16799) );
  BUF_X1 U1505 ( .A(n6076), .Z(n16800) );
  BUF_X1 U1506 ( .A(n6076), .Z(n16801) );
  BUF_X1 U1507 ( .A(n6076), .Z(n16802) );
  BUF_X1 U1508 ( .A(n5889), .Z(n16803) );
  BUF_X1 U1509 ( .A(n5889), .Z(n16804) );
  BUF_X1 U1510 ( .A(n5889), .Z(n16805) );
  BUF_X1 U1511 ( .A(n5889), .Z(n16806) );
  BUF_X1 U1512 ( .A(n5889), .Z(n16807) );
  BUF_X1 U1513 ( .A(n5889), .Z(n16808) );
  BUF_X1 U1514 ( .A(n5717), .Z(n16809) );
  BUF_X1 U1515 ( .A(n5717), .Z(n16810) );
  BUF_X1 U1516 ( .A(n5717), .Z(n16811) );
  BUF_X1 U1517 ( .A(n5717), .Z(n16812) );
  BUF_X1 U1518 ( .A(n5717), .Z(n16813) );
  BUF_X1 U1519 ( .A(n5717), .Z(n16814) );
  BUF_X1 U1520 ( .A(n5530), .Z(n16815) );
  BUF_X1 U1521 ( .A(n5530), .Z(n16816) );
  BUF_X1 U1522 ( .A(n5530), .Z(n16817) );
  BUF_X1 U1523 ( .A(n5530), .Z(n16818) );
  BUF_X1 U1524 ( .A(n5530), .Z(n16819) );
  BUF_X1 U1525 ( .A(n5530), .Z(n16820) );
  BUF_X1 U1526 ( .A(n5343), .Z(n16821) );
  BUF_X1 U1527 ( .A(n5343), .Z(n16822) );
  BUF_X1 U1528 ( .A(n5343), .Z(n16823) );
  BUF_X1 U1529 ( .A(n5343), .Z(n16824) );
  BUF_X1 U1530 ( .A(n5343), .Z(n16825) );
  BUF_X1 U1531 ( .A(n5343), .Z(n16826) );
  BUF_X1 U1532 ( .A(n5157), .Z(n16827) );
  BUF_X1 U1533 ( .A(n5157), .Z(n16828) );
  BUF_X1 U1534 ( .A(n5157), .Z(n16829) );
  BUF_X1 U1535 ( .A(n5157), .Z(n16830) );
  BUF_X1 U1536 ( .A(n5157), .Z(n16831) );
  BUF_X1 U1537 ( .A(n5157), .Z(n16832) );
  BUF_X1 U1538 ( .A(n5040), .Z(n16833) );
  BUF_X1 U1539 ( .A(n5040), .Z(n16834) );
  BUF_X1 U1540 ( .A(n5040), .Z(n16835) );
  BUF_X1 U1541 ( .A(n5040), .Z(n16836) );
  BUF_X1 U1542 ( .A(n5040), .Z(n16837) );
  BUF_X1 U1543 ( .A(n5040), .Z(n16838) );
  BUF_X1 U1544 ( .A(n4924), .Z(n16839) );
  BUF_X1 U1545 ( .A(n4924), .Z(n16840) );
  BUF_X1 U1546 ( .A(n4924), .Z(n16841) );
  BUF_X1 U1547 ( .A(n4924), .Z(n16842) );
  BUF_X1 U1548 ( .A(n4924), .Z(n16843) );
  BUF_X1 U1549 ( .A(n4924), .Z(n16844) );
  BUF_X1 U1550 ( .A(n4791), .Z(n16845) );
  BUF_X1 U1551 ( .A(n4791), .Z(n16846) );
  BUF_X1 U1552 ( .A(n4791), .Z(n16847) );
  BUF_X1 U1553 ( .A(n4791), .Z(n16848) );
  BUF_X1 U1554 ( .A(n4791), .Z(n16849) );
  BUF_X1 U1555 ( .A(n4791), .Z(n16850) );
  BUF_X1 U1556 ( .A(n4664), .Z(n16851) );
  BUF_X1 U1557 ( .A(n4664), .Z(n16852) );
  BUF_X1 U1558 ( .A(n4664), .Z(n16853) );
  BUF_X1 U1559 ( .A(n4664), .Z(n16854) );
  BUF_X1 U1560 ( .A(n4664), .Z(n16855) );
  BUF_X1 U1561 ( .A(n4664), .Z(n16856) );
  BUF_X1 U1562 ( .A(n4533), .Z(n16857) );
  BUF_X1 U1563 ( .A(n4533), .Z(n16858) );
  BUF_X1 U1564 ( .A(n4533), .Z(n16859) );
  BUF_X1 U1565 ( .A(n4533), .Z(n16860) );
  BUF_X1 U1566 ( .A(n4533), .Z(n16861) );
  BUF_X1 U1567 ( .A(n4533), .Z(n16862) );
  BUF_X1 U1568 ( .A(n4278), .Z(n17512) );
  BUF_X1 U1569 ( .A(n4278), .Z(n17513) );
  BUF_X1 U1570 ( .A(n4278), .Z(n17514) );
  BUF_X1 U1571 ( .A(n4278), .Z(n17515) );
  BUF_X1 U1572 ( .A(n4278), .Z(n17516) );
  BUF_X1 U1573 ( .A(n4278), .Z(n17517) );
  BUF_X1 U1574 ( .A(n10510), .Z(n16706) );
  BUF_X1 U1575 ( .A(n10510), .Z(n16705) );
  BUF_X1 U1576 ( .A(n10510), .Z(n16704) );
  BUF_X1 U1577 ( .A(n10510), .Z(n16703) );
  BUF_X1 U1578 ( .A(n7652), .Z(n16725) );
  BUF_X1 U1579 ( .A(n7652), .Z(n16726) );
  BUF_X1 U1580 ( .A(n7652), .Z(n16727) );
  BUF_X1 U1581 ( .A(n7652), .Z(n16728) );
  BUF_X1 U1582 ( .A(n7652), .Z(n16729) );
  BUF_X1 U1583 ( .A(n12338), .Z(n16436) );
  BUF_X1 U1584 ( .A(n12338), .Z(n16437) );
  BUF_X1 U1585 ( .A(n12338), .Z(n16438) );
  BUF_X1 U1586 ( .A(n12184), .Z(n16442) );
  BUF_X1 U1587 ( .A(n12184), .Z(n16443) );
  BUF_X1 U1588 ( .A(n12184), .Z(n16444) );
  BUF_X1 U1589 ( .A(n12029), .Z(n16448) );
  BUF_X1 U1590 ( .A(n12029), .Z(n16449) );
  BUF_X1 U1591 ( .A(n12029), .Z(n16450) );
  OAI21_X1 U1592 ( .B1(n14074), .B2(n14248), .A(n18044), .ZN(n4441) );
  OAI21_X1 U1593 ( .B1(n12414), .B2(n14248), .A(n18043), .ZN(n4417) );
  OAI21_X1 U1594 ( .B1(n14058), .B2(n14248), .A(n18043), .ZN(n4412) );
  OAI21_X1 U1595 ( .B1(n14228), .B2(n14248), .A(n18043), .ZN(n4409) );
  OAI21_X1 U1596 ( .B1(n14226), .B2(n14248), .A(n18043), .ZN(n4406) );
  OAI21_X1 U1597 ( .B1(n14222), .B2(n14248), .A(n18043), .ZN(n4401) );
  OAI21_X1 U1598 ( .B1(n14221), .B2(n14248), .A(n18042), .ZN(n4398) );
  OAI21_X1 U1599 ( .B1(n14218), .B2(n14248), .A(n18043), .ZN(n4391) );
  OAI21_X1 U1600 ( .B1(n14215), .B2(n14248), .A(n18042), .ZN(n4388) );
  BUF_X1 U1601 ( .A(n12523), .Z(n16424) );
  BUF_X1 U1602 ( .A(n12523), .Z(n16425) );
  BUF_X1 U1603 ( .A(n10520), .Z(n16677) );
  BUF_X1 U1604 ( .A(n10520), .Z(n16676) );
  BUF_X1 U1605 ( .A(n10663), .Z(n16464) );
  OAI21_X1 U1606 ( .B1(n14058), .B2(n14059), .A(n18039), .ZN(n4059) );
  BUF_X1 U1607 ( .A(n12524), .Z(n16421) );
  BUF_X1 U1608 ( .A(n12519), .Z(n16433) );
  BUF_X1 U1609 ( .A(n12524), .Z(n16422) );
  BUF_X1 U1610 ( .A(n12519), .Z(n16434) );
  BUF_X1 U1611 ( .A(n10522), .Z(n16674) );
  BUF_X1 U1612 ( .A(n10516), .Z(n16686) );
  BUF_X1 U1613 ( .A(n10522), .Z(n16673) );
  BUF_X1 U1614 ( .A(n10516), .Z(n16685) );
  BUF_X1 U1615 ( .A(n4153), .Z(n17756) );
  BUF_X1 U1616 ( .A(n4198), .Z(n17696) );
  BUF_X1 U1617 ( .A(n4233), .Z(n17648) );
  BUF_X1 U1618 ( .A(n4207), .Z(n17684) );
  BUF_X1 U1619 ( .A(n4220), .Z(n17672) );
  BUF_X1 U1620 ( .A(n4142), .Z(n17768) );
  BUF_X1 U1621 ( .A(n4189), .Z(n17708) );
  BUF_X1 U1622 ( .A(n4168), .Z(n17737) );
  BUF_X1 U1623 ( .A(n4237), .Z(n17641) );
  BUF_X1 U1624 ( .A(n4168), .Z(n17736) );
  BUF_X1 U1625 ( .A(n4237), .Z(n17640) );
  BUF_X1 U1626 ( .A(n4230), .Z(n17653) );
  BUF_X1 U1627 ( .A(n4230), .Z(n17652) );
  BUF_X1 U1628 ( .A(n4159), .Z(n17749) );
  BUF_X1 U1629 ( .A(n4211), .Z(n17677) );
  BUF_X1 U1630 ( .A(n4159), .Z(n17748) );
  BUF_X1 U1631 ( .A(n4211), .Z(n17676) );
  BUF_X1 U1632 ( .A(n4135), .Z(n17773) );
  BUF_X1 U1633 ( .A(n4135), .Z(n17772) );
  BUF_X1 U1634 ( .A(n4175), .Z(n17725) );
  BUF_X1 U1635 ( .A(n4186), .Z(n17713) );
  BUF_X1 U1636 ( .A(n4175), .Z(n17724) );
  BUF_X1 U1637 ( .A(n4186), .Z(n17712) );
  BUF_X1 U1638 ( .A(n4150), .Z(n17761) );
  BUF_X1 U1639 ( .A(n4150), .Z(n17760) );
  BUF_X1 U1640 ( .A(n4161), .Z(n17746) );
  BUF_X1 U1641 ( .A(n4195), .Z(n17698) );
  BUF_X1 U1642 ( .A(n4161), .Z(n17745) );
  BUF_X1 U1643 ( .A(n4195), .Z(n17697) );
  BUF_X1 U1644 ( .A(n4232), .Z(n17650) );
  BUF_X1 U1645 ( .A(n4232), .Z(n17649) );
  BUF_X1 U1646 ( .A(n4206), .Z(n17686) );
  BUF_X1 U1647 ( .A(n4206), .Z(n17685) );
  BUF_X1 U1648 ( .A(n4188), .Z(n17710) );
  BUF_X1 U1649 ( .A(n4219), .Z(n17674) );
  BUF_X1 U1650 ( .A(n4188), .Z(n17709) );
  BUF_X1 U1651 ( .A(n4219), .Z(n17673) );
  BUF_X1 U1652 ( .A(n4141), .Z(n17770) );
  BUF_X1 U1653 ( .A(n4181), .Z(n17722) );
  BUF_X1 U1654 ( .A(n4225), .Z(n17662) );
  BUF_X1 U1655 ( .A(n4239), .Z(n17638) );
  BUF_X1 U1656 ( .A(n4114), .Z(n17806) );
  BUF_X1 U1657 ( .A(n4141), .Z(n17769) );
  BUF_X1 U1658 ( .A(n4181), .Z(n17721) );
  BUF_X1 U1659 ( .A(n4225), .Z(n17661) );
  BUF_X1 U1660 ( .A(n4239), .Z(n17637) );
  BUF_X1 U1661 ( .A(n4114), .Z(n17805) );
  BUF_X1 U1662 ( .A(n4200), .Z(n17692) );
  BUF_X1 U1663 ( .A(n4209), .Z(n17680) );
  BUF_X1 U1664 ( .A(n4200), .Z(n17691) );
  BUF_X1 U1665 ( .A(n4209), .Z(n17679) );
  BUF_X1 U1666 ( .A(n4157), .Z(n17752) );
  BUF_X1 U1667 ( .A(n4235), .Z(n17644) );
  BUF_X1 U1668 ( .A(n4228), .Z(n17656) );
  BUF_X1 U1669 ( .A(n4157), .Z(n17751) );
  BUF_X1 U1670 ( .A(n4235), .Z(n17643) );
  BUF_X1 U1671 ( .A(n4228), .Z(n17655) );
  BUF_X1 U1672 ( .A(n12633), .Z(n16214) );
  BUF_X1 U1673 ( .A(n12633), .Z(n16215) );
  BUF_X1 U1674 ( .A(n12525), .Z(n16418) );
  BUF_X1 U1675 ( .A(n12520), .Z(n16430) );
  BUF_X1 U1676 ( .A(n12525), .Z(n16419) );
  BUF_X1 U1677 ( .A(n12520), .Z(n16431) );
  BUF_X1 U1678 ( .A(n4124), .Z(n17792) );
  BUF_X1 U1679 ( .A(n4131), .Z(n17780) );
  BUF_X1 U1680 ( .A(n4171), .Z(n17732) );
  BUF_X1 U1681 ( .A(n4184), .Z(n17716) );
  BUF_X1 U1682 ( .A(n4119), .Z(n17800) );
  BUF_X1 U1683 ( .A(n4126), .Z(n17788) );
  BUF_X1 U1684 ( .A(n4133), .Z(n17776) );
  BUF_X1 U1685 ( .A(n4184), .Z(n17715) );
  BUF_X1 U1686 ( .A(n4119), .Z(n17799) );
  BUF_X1 U1687 ( .A(n4126), .Z(n17787) );
  BUF_X1 U1688 ( .A(n4133), .Z(n17775) );
  BUF_X1 U1689 ( .A(n4173), .Z(n17728) );
  BUF_X1 U1690 ( .A(n4242), .Z(n17632) );
  BUF_X1 U1691 ( .A(n4173), .Z(n17727) );
  BUF_X1 U1692 ( .A(n4242), .Z(n17631) );
  BUF_X1 U1693 ( .A(n4170), .Z(n17734) );
  BUF_X1 U1694 ( .A(n4107), .Z(n17818) );
  BUF_X1 U1695 ( .A(n4123), .Z(n17794) );
  BUF_X1 U1696 ( .A(n4130), .Z(n17782) );
  BUF_X1 U1697 ( .A(n4170), .Z(n17733) );
  BUF_X1 U1698 ( .A(n4107), .Z(n17817) );
  BUF_X1 U1699 ( .A(n4123), .Z(n17793) );
  BUF_X1 U1700 ( .A(n4130), .Z(n17781) );
  BUF_X1 U1701 ( .A(n4148), .Z(n17764) );
  BUF_X1 U1702 ( .A(n4191), .Z(n17704) );
  BUF_X1 U1703 ( .A(n4222), .Z(n17668) );
  BUF_X1 U1704 ( .A(n4148), .Z(n17763) );
  BUF_X1 U1705 ( .A(n4191), .Z(n17703) );
  BUF_X1 U1706 ( .A(n4222), .Z(n17667) );
  BUF_X1 U1707 ( .A(n12522), .Z(n16429) );
  NOR2_X1 U1708 ( .A1(n13975), .A2(n13976), .ZN(n13970) );
  NOR2_X1 U1709 ( .A1(n12494), .A2(n12495), .ZN(n12489) );
  BUF_X1 U1710 ( .A(n12523), .Z(n16426) );
  BUF_X1 U1711 ( .A(n12634), .Z(n16212) );
  BUF_X1 U1712 ( .A(n12634), .Z(n16211) );
  NAND2_X1 U1713 ( .A1(n14260), .A2(n14253), .ZN(n14215) );
  NAND2_X1 U1714 ( .A1(n13932), .A2(n13960), .ZN(n12615) );
  BUF_X1 U1715 ( .A(n12524), .Z(n16423) );
  BUF_X1 U1716 ( .A(n12519), .Z(n16435) );
  BUF_X1 U1717 ( .A(n10520), .Z(n16678) );
  NAND2_X1 U1718 ( .A1(n14260), .A2(n14251), .ZN(n14222) );
  NAND2_X1 U1719 ( .A1(n14260), .A2(n14249), .ZN(n14221) );
  NAND2_X1 U1720 ( .A1(n14253), .A2(n14250), .ZN(n14226) );
  NAND2_X1 U1721 ( .A1(n14260), .A2(n14254), .ZN(n14218) );
  NAND2_X1 U1722 ( .A1(n14254), .A2(n14250), .ZN(n14228) );
  BUF_X1 U1723 ( .A(n4161), .Z(n17747) );
  BUF_X1 U1724 ( .A(n4195), .Z(n17699) );
  BUF_X1 U1725 ( .A(n4232), .Z(n17651) );
  BUF_X1 U1726 ( .A(n4168), .Z(n17738) );
  BUF_X1 U1727 ( .A(n4237), .Z(n17642) );
  BUF_X1 U1728 ( .A(n4230), .Z(n17654) );
  BUF_X1 U1729 ( .A(n4206), .Z(n17687) );
  BUF_X1 U1730 ( .A(n4188), .Z(n17711) );
  BUF_X1 U1731 ( .A(n4219), .Z(n17675) );
  BUF_X1 U1732 ( .A(n4159), .Z(n17750) );
  BUF_X1 U1733 ( .A(n4211), .Z(n17678) );
  BUF_X1 U1734 ( .A(n4141), .Z(n17771) );
  BUF_X1 U1735 ( .A(n4181), .Z(n17723) );
  BUF_X1 U1736 ( .A(n4225), .Z(n17663) );
  BUF_X1 U1737 ( .A(n4239), .Z(n17639) );
  BUF_X1 U1738 ( .A(n4114), .Z(n17807) );
  BUF_X1 U1739 ( .A(n10522), .Z(n16675) );
  BUF_X1 U1740 ( .A(n10516), .Z(n16687) );
  BUF_X1 U1741 ( .A(n4135), .Z(n17774) );
  BUF_X1 U1742 ( .A(n4200), .Z(n17693) );
  BUF_X1 U1743 ( .A(n4209), .Z(n17681) );
  BUF_X1 U1744 ( .A(n4175), .Z(n17726) );
  BUF_X1 U1745 ( .A(n4186), .Z(n17714) );
  BUF_X1 U1746 ( .A(n4157), .Z(n17753) );
  BUF_X1 U1747 ( .A(n4235), .Z(n17645) );
  BUF_X1 U1748 ( .A(n4228), .Z(n17657) );
  BUF_X1 U1749 ( .A(n4150), .Z(n17762) );
  NAND2_X1 U1750 ( .A1(n14251), .A2(n14250), .ZN(n12414) );
  BUF_X1 U1751 ( .A(n12624), .Z(n16237) );
  BUF_X1 U1752 ( .A(n12633), .Z(n16216) );
  BUF_X1 U1753 ( .A(n12525), .Z(n16420) );
  BUF_X1 U1754 ( .A(n12520), .Z(n16432) );
  BUF_X1 U1755 ( .A(n4184), .Z(n17717) );
  BUF_X1 U1756 ( .A(n4119), .Z(n17801) );
  BUF_X1 U1757 ( .A(n4126), .Z(n17789) );
  BUF_X1 U1758 ( .A(n4133), .Z(n17777) );
  BUF_X1 U1759 ( .A(n4173), .Z(n17729) );
  BUF_X1 U1760 ( .A(n4242), .Z(n17633) );
  BUF_X1 U1761 ( .A(n4123), .Z(n17795) );
  BUF_X1 U1762 ( .A(n4130), .Z(n17783) );
  BUF_X1 U1763 ( .A(n4170), .Z(n17735) );
  BUF_X1 U1764 ( .A(n4107), .Z(n17819) );
  BUF_X1 U1765 ( .A(n4148), .Z(n17765) );
  BUF_X1 U1766 ( .A(n4191), .Z(n17705) );
  BUF_X1 U1767 ( .A(n4222), .Z(n17669) );
  NAND2_X1 U1768 ( .A1(n12452), .A2(n12479), .ZN(n10635) );
  NAND2_X1 U1769 ( .A1(n14249), .A2(n14250), .ZN(n14058) );
  NAND2_X1 U1770 ( .A1(n14138), .A2(n14205), .ZN(n14089) );
  NAND2_X1 U1771 ( .A1(n14137), .A2(n14205), .ZN(n14098) );
  OAI21_X1 U1772 ( .B1(n14066), .B2(n14237), .A(n18041), .ZN(n4317) );
  BUF_X1 U1773 ( .A(n12634), .Z(n16213) );
  BUF_X1 U1774 ( .A(n4088), .Z(n17835) );
  OAI21_X1 U1775 ( .B1(n14059), .B2(n14074), .A(n18040), .ZN(n4088) );
  BUF_X1 U1776 ( .A(n4085), .Z(n17857) );
  OAI21_X1 U1777 ( .B1(n14059), .B2(n14073), .A(n18040), .ZN(n4085) );
  BUF_X1 U1778 ( .A(n4082), .Z(n17879) );
  OAI21_X1 U1779 ( .B1(n14059), .B2(n14072), .A(n18040), .ZN(n4082) );
  BUF_X1 U1780 ( .A(n4079), .Z(n17901) );
  OAI21_X1 U1781 ( .B1(n14059), .B2(n14070), .A(n18039), .ZN(n4079) );
  OAI21_X1 U1782 ( .B1(n14064), .B2(n14252), .A(n18043), .ZN(n4426) );
  OAI21_X1 U1783 ( .B1(n14064), .B2(n14237), .A(n18041), .ZN(n4312) );
  INV_X1 U1784 ( .A(n14207), .ZN(n14197) );
  NAND2_X1 U1785 ( .A1(n14245), .A2(n14067), .ZN(n14244) );
  INV_X1 U1786 ( .A(n14241), .ZN(n14245) );
  NAND2_X1 U1787 ( .A1(n14256), .A2(n14067), .ZN(n14252) );
  INV_X1 U1788 ( .A(n14248), .ZN(n14256) );
  NAND2_X1 U1789 ( .A1(n14238), .A2(n14067), .ZN(n14237) );
  INV_X1 U1790 ( .A(n14236), .ZN(n14238) );
  NAND2_X1 U1791 ( .A1(n14258), .A2(n14253), .ZN(n14070) );
  NAND2_X1 U1792 ( .A1(n14143), .A2(n14205), .ZN(n14097) );
  NAND2_X1 U1793 ( .A1(n14202), .A2(n14205), .ZN(n14201) );
  NAND2_X1 U1794 ( .A1(n14067), .A2(n14068), .ZN(n14061) );
  INV_X1 U1795 ( .A(n14059), .ZN(n14068) );
  NAND2_X1 U1796 ( .A1(n14258), .A2(n14254), .ZN(n14072) );
  INV_X1 U1797 ( .A(n14183), .ZN(n14176) );
  AND2_X1 U1798 ( .A1(n14000), .A2(n14001), .ZN(n14004) );
  INV_X1 U1799 ( .A(n14096), .ZN(n14087) );
  NAND2_X1 U1800 ( .A1(n13946), .A2(n13932), .ZN(n12575) );
  NAND2_X1 U1801 ( .A1(n13926), .A2(n13932), .ZN(n12550) );
  NAND2_X1 U1802 ( .A1(n13936), .A2(n13932), .ZN(n12606) );
  NAND2_X1 U1803 ( .A1(n13955), .A2(n13932), .ZN(n12621) );
  NAND2_X1 U1804 ( .A1(n13969), .A2(n13932), .ZN(n12622) );
  BUF_X1 U1805 ( .A(n10649), .Z(n16489) );
  NAND2_X1 U1806 ( .A1(n12465), .A2(n12452), .ZN(n10592) );
  NAND2_X1 U1807 ( .A1(n12455), .A2(n12452), .ZN(n10624) );
  NAND2_X1 U1808 ( .A1(n12477), .A2(n12452), .ZN(n10644) );
  NAND2_X1 U1809 ( .A1(n12488), .A2(n12452), .ZN(n10646) );
  BUF_X1 U1810 ( .A(n10662), .Z(n16468) );
  BUF_X1 U1811 ( .A(n10523), .Z(n16672) );
  BUF_X1 U1812 ( .A(n10517), .Z(n16684) );
  AND2_X1 U1813 ( .A1(n12463), .A2(n12456), .ZN(n12465) );
  AND2_X1 U1814 ( .A1(n13944), .A2(n13937), .ZN(n13946) );
  BUF_X1 U1815 ( .A(n10519), .Z(n16681) );
  AND2_X1 U1816 ( .A1(n12444), .A2(n12480), .ZN(n12455) );
  AND2_X1 U1817 ( .A1(n13921), .A2(n13961), .ZN(n13936) );
  INV_X1 U1818 ( .A(n14253), .ZN(n14062) );
  AND2_X1 U1819 ( .A1(n13970), .A2(n13932), .ZN(n13925) );
  AND2_X1 U1820 ( .A1(n13957), .A2(n13937), .ZN(n13960) );
  AND2_X1 U1821 ( .A1(n12489), .A2(n12452), .ZN(n12443) );
  AND2_X1 U1822 ( .A1(n12474), .A2(n12456), .ZN(n12479) );
  BUF_X1 U1823 ( .A(n10663), .Z(n16465) );
  NAND2_X1 U1824 ( .A1(n12451), .A2(n12479), .ZN(n10626) );
  NAND2_X1 U1825 ( .A1(n18044), .A2(n14000), .ZN(n14001) );
  INV_X1 U1826 ( .A(n14254), .ZN(n14063) );
  NAND2_X1 U1827 ( .A1(n13927), .A2(n13960), .ZN(n12607) );
  NAND2_X1 U1828 ( .A1(n13935), .A2(n13969), .ZN(n12617) );
  NAND2_X1 U1829 ( .A1(n12454), .A2(n12488), .ZN(n10639) );
  INV_X1 U1830 ( .A(n14134), .ZN(n14094) );
  AND2_X1 U1831 ( .A1(n12463), .A2(n12480), .ZN(n12472) );
  AND2_X1 U1832 ( .A1(n13944), .A2(n13961), .ZN(n13953) );
  AND2_X1 U1833 ( .A1(n13920), .A2(n13961), .ZN(n13917) );
  AND2_X1 U1834 ( .A1(n12439), .A2(n12480), .ZN(n12436) );
  AND2_X1 U1835 ( .A1(n13921), .A2(n13937), .ZN(n13926) );
  INV_X1 U1836 ( .A(n14066), .ZN(n14251) );
  NAND2_X1 U1837 ( .A1(n12465), .A2(n12451), .ZN(n10585) );
  NAND2_X1 U1838 ( .A1(n12450), .A2(n12451), .ZN(n10552) );
  NAND2_X1 U1839 ( .A1(n12455), .A2(n12451), .ZN(n10558) );
  NAND2_X1 U1840 ( .A1(n12477), .A2(n12451), .ZN(n10617) );
  NAND2_X1 U1841 ( .A1(n12472), .A2(n12451), .ZN(n10603) );
  NAND2_X1 U1842 ( .A1(n12436), .A2(n12451), .ZN(n10658) );
  NAND2_X1 U1843 ( .A1(n13946), .A2(n13927), .ZN(n12580) );
  NAND2_X1 U1844 ( .A1(n13926), .A2(n13927), .ZN(n12545) );
  NAND2_X1 U1845 ( .A1(n13936), .A2(n13927), .ZN(n12555) );
  NAND2_X1 U1846 ( .A1(n13953), .A2(n13927), .ZN(n12589) );
  NAND2_X1 U1847 ( .A1(n13917), .A2(n13927), .ZN(n12631) );
  AND2_X1 U1848 ( .A1(n12475), .A2(n12454), .ZN(n12445) );
  AND2_X1 U1849 ( .A1(n13961), .A2(n13957), .ZN(n13969) );
  AND2_X1 U1850 ( .A1(n12480), .A2(n12474), .ZN(n12488) );
  INV_X1 U1851 ( .A(n14064), .ZN(n14249) );
  AND2_X1 U1852 ( .A1(n13958), .A2(n13927), .ZN(n13929) );
  AND2_X1 U1853 ( .A1(n13958), .A2(n13935), .ZN(n13922) );
  NAND2_X1 U1854 ( .A1(n12463), .A2(n12440), .ZN(n10619) );
  NAND2_X1 U1855 ( .A1(n12463), .A2(n12443), .ZN(n10610) );
  AND2_X1 U1856 ( .A1(n12444), .A2(n12456), .ZN(n12450) );
  AND2_X1 U1857 ( .A1(n12439), .A2(n12456), .ZN(n12477) );
  INV_X1 U1858 ( .A(n14131), .ZN(n14104) );
  NAND2_X1 U1859 ( .A1(n13944), .A2(n13925), .ZN(n12594) );
  NAND2_X1 U1860 ( .A1(n13922), .A2(n13957), .ZN(n12601) );
  NAND2_X1 U1861 ( .A1(n13929), .A2(n13957), .ZN(n12599) );
  NAND2_X1 U1862 ( .A1(n13928), .A2(n13957), .ZN(n12627) );
  NAND2_X1 U1863 ( .A1(n13925), .A2(n13957), .ZN(n12626) );
  NAND2_X1 U1864 ( .A1(n13936), .A2(n13935), .ZN(n12565) );
  NAND2_X1 U1865 ( .A1(n13946), .A2(n13935), .ZN(n12581) );
  NAND2_X1 U1866 ( .A1(n13926), .A2(n13935), .ZN(n12556) );
  NAND2_X1 U1867 ( .A1(n13953), .A2(n13935), .ZN(n12590) );
  NAND2_X1 U1868 ( .A1(n13917), .A2(n13935), .ZN(n12632) );
  NAND2_X1 U1869 ( .A1(n12455), .A2(n12454), .ZN(n10571) );
  NAND2_X1 U1870 ( .A1(n12465), .A2(n12454), .ZN(n10587) );
  NAND2_X1 U1871 ( .A1(n12450), .A2(n12454), .ZN(n10560) );
  NAND2_X1 U1872 ( .A1(n12472), .A2(n12454), .ZN(n10605) );
  NAND2_X1 U1873 ( .A1(n12436), .A2(n12454), .ZN(n10660) );
  NAND2_X1 U1874 ( .A1(n12445), .A2(n12463), .ZN(n10580) );
  NAND2_X1 U1875 ( .A1(n12447), .A2(n12463), .ZN(n10578) );
  AND2_X1 U1876 ( .A1(n13958), .A2(n13932), .ZN(n13931) );
  AND2_X1 U1877 ( .A1(n12475), .A2(n12452), .ZN(n12449) );
  NAND2_X1 U1878 ( .A1(n12444), .A2(n12441), .ZN(n10569) );
  NAND2_X1 U1879 ( .A1(n12444), .A2(n12449), .ZN(n10554) );
  NAND2_X1 U1880 ( .A1(n12444), .A2(n12445), .ZN(n10545) );
  NAND2_X1 U1881 ( .A1(n13922), .A2(n13944), .ZN(n12571) );
  NAND2_X1 U1882 ( .A1(n13929), .A2(n13944), .ZN(n12570) );
  INV_X1 U1883 ( .A(n14145), .ZN(n14107) );
  NAND2_X1 U1884 ( .A1(n12440), .A2(n12474), .ZN(n10653) );
  NAND2_X1 U1885 ( .A1(n12443), .A2(n12474), .ZN(n10651) );
  NAND2_X1 U1886 ( .A1(n14108), .A2(n14085), .ZN(n4164) );
  NAND2_X1 U1887 ( .A1(n13921), .A2(n13931), .ZN(n12552) );
  NAND2_X1 U1888 ( .A1(n13921), .A2(n13923), .ZN(n12564) );
  AND2_X1 U1889 ( .A1(n12489), .A2(n12451), .ZN(n12441) );
  AND2_X1 U1890 ( .A1(n13970), .A2(n13927), .ZN(n13923) );
  AND2_X1 U1891 ( .A1(n13917), .A2(n13932), .ZN(n12577) );
  AND2_X1 U1892 ( .A1(n13953), .A2(n13932), .ZN(n12629) );
  AND2_X1 U1893 ( .A1(n12436), .A2(n12452), .ZN(n10589) );
  AND2_X1 U1894 ( .A1(n12450), .A2(n12452), .ZN(n10550) );
  AND2_X1 U1895 ( .A1(n12472), .A2(n12452), .ZN(n10656) );
  AND2_X1 U1896 ( .A1(n13970), .A2(n13935), .ZN(n13919) );
  AND2_X1 U1897 ( .A1(n12489), .A2(n12454), .ZN(n12438) );
  AND2_X1 U1898 ( .A1(n12475), .A2(n12451), .ZN(n12447) );
  AND2_X1 U1899 ( .A1(n13920), .A2(n13937), .ZN(n13955) );
  AND2_X1 U1900 ( .A1(n12451), .A2(n12488), .ZN(n10632) );
  AND2_X1 U1901 ( .A1(n13927), .A2(n13969), .ZN(n12612) );
  AND2_X1 U1902 ( .A1(n13935), .A2(n13960), .ZN(n12604) );
  AND2_X1 U1903 ( .A1(n12454), .A2(n12479), .ZN(n10622) );
  AND2_X1 U1904 ( .A1(n12463), .A2(n12441), .ZN(n10601) );
  AND2_X1 U1905 ( .A1(n12463), .A2(n12438), .ZN(n10607) );
  AND2_X1 U1906 ( .A1(n13955), .A2(n13927), .ZN(n12592) );
  AND2_X1 U1907 ( .A1(n13955), .A2(n13935), .ZN(n12618) );
  AND2_X1 U1908 ( .A1(n12477), .A2(n12454), .ZN(n10641) );
  AND2_X1 U1909 ( .A1(n13944), .A2(n13923), .ZN(n12587) );
  AND2_X1 U1910 ( .A1(n13944), .A2(n13919), .ZN(n12591) );
  AND2_X1 U1911 ( .A1(n13944), .A2(n13928), .ZN(n12596) );
  AND2_X1 U1912 ( .A1(n12444), .A2(n12438), .ZN(n10567) );
  AND2_X1 U1913 ( .A1(n12444), .A2(n12440), .ZN(n10575) );
  AND2_X1 U1914 ( .A1(n12444), .A2(n12443), .ZN(n10576) );
  AND2_X1 U1915 ( .A1(n12444), .A2(n12447), .ZN(n10542) );
  AND2_X1 U1916 ( .A1(n12444), .A2(n12446), .ZN(n10543) );
  AND2_X1 U1917 ( .A1(n13921), .A2(n13919), .ZN(n12562) );
  AND2_X1 U1918 ( .A1(n13921), .A2(n13928), .ZN(n12567) );
  AND2_X1 U1919 ( .A1(n13921), .A2(n13925), .ZN(n12568) );
  AND2_X1 U1920 ( .A1(n13921), .A2(n13922), .ZN(n12538) );
  AND2_X1 U1921 ( .A1(n13921), .A2(n13929), .ZN(n12542) );
  AND2_X1 U1922 ( .A1(n13921), .A2(n13933), .ZN(n12548) );
  AND2_X1 U1923 ( .A1(n13931), .A2(n13957), .ZN(n12603) );
  AND2_X1 U1924 ( .A1(n13933), .A2(n13957), .ZN(n12597) );
  AND2_X1 U1925 ( .A1(n13923), .A2(n13957), .ZN(n12613) );
  AND2_X1 U1926 ( .A1(n13919), .A2(n13957), .ZN(n12623) );
  AND2_X1 U1927 ( .A1(n12446), .A2(n12463), .ZN(n10582) );
  AND2_X1 U1928 ( .A1(n12449), .A2(n12463), .ZN(n10583) );
  AND2_X1 U1929 ( .A1(n13933), .A2(n13944), .ZN(n12572) );
  AND2_X1 U1930 ( .A1(n13931), .A2(n13944), .ZN(n12573) );
  AND2_X1 U1931 ( .A1(n12445), .A2(n12474), .ZN(n10614) );
  AND2_X1 U1932 ( .A1(n12446), .A2(n12474), .ZN(n10615) );
  AND2_X1 U1933 ( .A1(n12449), .A2(n12474), .ZN(n10621) );
  AND2_X1 U1934 ( .A1(n12447), .A2(n12474), .ZN(n10608) );
  AND2_X1 U1935 ( .A1(n12441), .A2(n12474), .ZN(n10633) );
  AND2_X1 U1936 ( .A1(n12438), .A2(n12474), .ZN(n10648) );
  AND2_X1 U1937 ( .A1(n14108), .A2(n14087), .ZN(n4162) );
  BUF_X1 U1938 ( .A(n4462), .Z(n16877) );
  OAI21_X1 U1939 ( .B1(n14059), .B2(n14226), .A(n18044), .ZN(n4462) );
  BUF_X1 U1940 ( .A(n4459), .Z(n16887) );
  OAI21_X1 U1941 ( .B1(n14059), .B2(n14222), .A(n18044), .ZN(n4459) );
  BUF_X1 U1942 ( .A(n4451), .Z(n16910) );
  OAI21_X1 U1943 ( .B1(n14059), .B2(n14218), .A(n18044), .ZN(n4451) );
  OAI21_X1 U1944 ( .B1(n14059), .B2(n14215), .A(n18043), .ZN(n4448) );
  BUF_X1 U1945 ( .A(n4382), .Z(n17137) );
  OAI21_X1 U1946 ( .B1(n14073), .B2(n14241), .A(n18042), .ZN(n4382) );
  BUF_X1 U1947 ( .A(n4376), .Z(n17160) );
  OAI21_X1 U1948 ( .B1(n14070), .B2(n14241), .A(n18042), .ZN(n4376) );
  BUF_X1 U1949 ( .A(n4438), .Z(n16944) );
  OAI21_X1 U1950 ( .B1(n14073), .B2(n14248), .A(n18043), .ZN(n4438) );
  BUF_X1 U1951 ( .A(n4435), .Z(n16956) );
  OAI21_X1 U1952 ( .B1(n14072), .B2(n14248), .A(n18043), .ZN(n4435) );
  BUF_X1 U1953 ( .A(n4432), .Z(n16966) );
  OAI21_X1 U1954 ( .B1(n14070), .B2(n14248), .A(n18043), .ZN(n4432) );
  BUF_X1 U1955 ( .A(n4373), .Z(n17170) );
  OAI21_X1 U1956 ( .B1(n14066), .B2(n14244), .A(n18042), .ZN(n4373) );
  BUF_X1 U1957 ( .A(n4429), .Z(n16976) );
  OAI21_X1 U1958 ( .B1(n14066), .B2(n14252), .A(n18043), .ZN(n4429) );
  BUF_X1 U1959 ( .A(n4370), .Z(n17182) );
  OAI21_X1 U1960 ( .B1(n14064), .B2(n14244), .A(n18042), .ZN(n4370) );
  AND2_X1 U1961 ( .A1(n13958), .A2(n13918), .ZN(n13933) );
  AND2_X1 U1962 ( .A1(n12475), .A2(n12437), .ZN(n12446) );
  INV_X1 U1963 ( .A(n14133), .ZN(n14022) );
  BUF_X1 U1964 ( .A(n10425), .Z(n16707) );
  BUF_X1 U1965 ( .A(n10315), .Z(n16716) );
  BUF_X1 U1966 ( .A(n11868), .Z(n16454) );
  INV_X1 U1967 ( .A(n14180), .ZN(n14182) );
  INV_X1 U1968 ( .A(n14204), .ZN(n14208) );
  BUF_X1 U1969 ( .A(n10425), .Z(n16708) );
  BUF_X1 U1970 ( .A(n10315), .Z(n16717) );
  BUF_X1 U1971 ( .A(n11868), .Z(n16455) );
  BUF_X1 U1972 ( .A(n10511), .Z(n16688) );
  BUF_X1 U1973 ( .A(n4273), .Z(n17533) );
  BUF_X1 U1974 ( .A(n4270), .Z(n17547) );
  BUF_X1 U1975 ( .A(n4267), .Z(n17561) );
  BUF_X1 U1976 ( .A(n10511), .Z(n16689) );
  BUF_X1 U1977 ( .A(n4273), .Z(n17532) );
  BUF_X1 U1978 ( .A(n4270), .Z(n17546) );
  BUF_X1 U1979 ( .A(n4267), .Z(n17560) );
  BUF_X1 U1980 ( .A(n4273), .Z(n17531) );
  BUF_X1 U1981 ( .A(n4270), .Z(n17545) );
  BUF_X1 U1982 ( .A(n4267), .Z(n17559) );
  BUF_X1 U1983 ( .A(n4262), .Z(n17573) );
  BUF_X1 U1984 ( .A(n4259), .Z(n17588) );
  BUF_X1 U1985 ( .A(n4262), .Z(n17574) );
  BUF_X1 U1986 ( .A(n4259), .Z(n17587) );
  BUF_X1 U1987 ( .A(n4259), .Z(n17586) );
  BUF_X1 U1988 ( .A(n4256), .Z(n17602) );
  BUF_X1 U1989 ( .A(n4251), .Z(n17616) );
  BUF_X1 U1990 ( .A(n4256), .Z(n17601) );
  BUF_X1 U1991 ( .A(n4251), .Z(n17615) );
  BUF_X1 U1992 ( .A(n4256), .Z(n17600) );
  BUF_X1 U1993 ( .A(n4251), .Z(n17614) );
  BUF_X1 U1994 ( .A(n4090), .Z(n17822) );
  BUF_X1 U1995 ( .A(n10511), .Z(n16690) );
  BUF_X1 U1996 ( .A(n4262), .Z(n17575) );
  INV_X1 U1997 ( .A(n18032), .ZN(n18054) );
  INV_X1 U1998 ( .A(n18032), .ZN(n18055) );
  BUF_X1 U1999 ( .A(n12302), .Z(n16439) );
  BUF_X1 U2000 ( .A(n12302), .Z(n16440) );
  BUF_X1 U2001 ( .A(n12302), .Z(n16441) );
  BUF_X1 U2002 ( .A(n12149), .Z(n16445) );
  BUF_X1 U2003 ( .A(n12149), .Z(n16446) );
  BUF_X1 U2004 ( .A(n12149), .Z(n16447) );
  BUF_X1 U2005 ( .A(n11996), .Z(n16451) );
  BUF_X1 U2006 ( .A(n11996), .Z(n16452) );
  BUF_X1 U2007 ( .A(n11996), .Z(n16453) );
  BUF_X1 U2008 ( .A(n10400), .Z(n16714) );
  BUF_X1 U2009 ( .A(n10400), .Z(n16713) );
  BUF_X1 U2010 ( .A(n11843), .Z(n16461) );
  BUF_X1 U2011 ( .A(n11843), .Z(n16460) );
  BUF_X1 U2012 ( .A(n10290), .Z(n16723) );
  BUF_X1 U2013 ( .A(n10290), .Z(n16722) );
  BUF_X1 U2014 ( .A(n11843), .Z(n16462) );
  BUF_X1 U2015 ( .A(n10290), .Z(n16724) );
  BUF_X1 U2016 ( .A(n10400), .Z(n16715) );
  BUF_X1 U2017 ( .A(n4090), .Z(n17821) );
  BUF_X1 U2018 ( .A(n4090), .Z(n17820) );
  NOR3_X1 U2019 ( .A1(n14174), .A2(N9924), .A3(n14173), .ZN(n14151) );
  NAND4_X1 U2020 ( .A1(N9924), .A2(n14173), .A3(n14174), .A4(n14020), .ZN(
        n14096) );
  NAND3_X1 U2021 ( .A1(n14247), .A2(n14234), .A3(n14240), .ZN(n14248) );
  NOR2_X1 U2022 ( .A1(n17825), .A2(n14005), .ZN(n14034) );
  NAND3_X1 U2023 ( .A1(n14240), .A2(n14247), .A3(N276), .ZN(n14059) );
  NOR3_X1 U2024 ( .A1(n14006), .A2(n14231), .A3(n14266), .ZN(n14240) );
  INV_X1 U2025 ( .A(n14232), .ZN(n14266) );
  NOR3_X1 U2026 ( .A1(N9922), .A2(N9924), .A3(n14174), .ZN(n14091) );
  NAND4_X1 U2027 ( .A1(n14231), .A2(n14232), .A3(n14233), .A4(n14234), .ZN(
        n12415) );
  BUF_X1 U2028 ( .A(n12527), .Z(n16413) );
  BUF_X1 U2029 ( .A(n12527), .Z(n16412) );
  BUF_X1 U2030 ( .A(n10525), .Z(n16665) );
  BUF_X1 U2031 ( .A(n10525), .Z(n16664) );
  BUF_X1 U2032 ( .A(n12527), .Z(n16414) );
  BUF_X1 U2033 ( .A(n10525), .Z(n16666) );
  OAI22_X1 U2034 ( .A1(n14135), .A2(n14136), .B1(n14096), .B2(n14131), .ZN(
        n4153) );
  INV_X1 U2035 ( .A(n14129), .ZN(n14135) );
  OAI22_X1 U2036 ( .A1(n14144), .A2(n14136), .B1(n14145), .B2(n14096), .ZN(
        n4161) );
  OAI22_X1 U2037 ( .A1(n14172), .A2(n14142), .B1(n14089), .B2(n14096), .ZN(
        n4195) );
  OAI22_X1 U2038 ( .A1(n14172), .A2(n14101), .B1(n14098), .B2(n14096), .ZN(
        n4198) );
  OAI22_X1 U2039 ( .A1(n14181), .A2(n14208), .B1(n14207), .B2(n14184), .ZN(
        n4232) );
  OAI22_X1 U2040 ( .A1(n14208), .A2(n14185), .B1(n14207), .B2(n14186), .ZN(
        n4233) );
  OAI22_X1 U2041 ( .A1(n14185), .A2(n14182), .B1(n14183), .B2(n14186), .ZN(
        n4206) );
  OAI22_X1 U2042 ( .A1(n14181), .A2(n14182), .B1(n14183), .B2(n14184), .ZN(
        n4207) );
  OAI22_X1 U2043 ( .A1(n14163), .A2(n14115), .B1(n14164), .B2(n14117), .ZN(
        n4188) );
  OAI22_X1 U2044 ( .A1(n14163), .A2(n14122), .B1(n14164), .B2(n14123), .ZN(
        n4219) );
  NAND2_X1 U2045 ( .A1(N9925), .A2(n14197), .ZN(n14164) );
  OAI22_X1 U2046 ( .A1(n14120), .A2(n14159), .B1(n14121), .B2(n14160), .ZN(
        n4220) );
  OAI22_X1 U2047 ( .A1(n14124), .A2(n14116), .B1(n14125), .B2(n14118), .ZN(
        n4141) );
  OAI22_X1 U2048 ( .A1(n14159), .A2(n14116), .B1(n14160), .B2(n14118), .ZN(
        n4181) );
  OAI22_X1 U2049 ( .A1(n14122), .A2(n14116), .B1(n14123), .B2(n14118), .ZN(
        n4239) );
  OAI22_X1 U2050 ( .A1(n14122), .A2(n14166), .B1(n14123), .B2(n14167), .ZN(
        n4189) );
  OAI22_X1 U2051 ( .A1(n14159), .A2(n14166), .B1(n14160), .B2(n14167), .ZN(
        n4225) );
  OAI22_X1 U2052 ( .A1(n14122), .A2(n14120), .B1(n14123), .B2(n14121), .ZN(
        n4142) );
  OAI22_X1 U2053 ( .A1(n14098), .A2(n14099), .B1(n14100), .B2(n14101), .ZN(
        n4114) );
  NOR2_X1 U2054 ( .A1(n14259), .A2(N275), .ZN(n14250) );
  AOI22_X1 U2055 ( .A1(n14140), .A2(n14141), .B1(n14105), .B2(n14086), .ZN(
        n4168) );
  INV_X1 U2056 ( .A(n14142), .ZN(n14141) );
  AOI22_X1 U2057 ( .A1(n14140), .A2(n14171), .B1(n14105), .B2(n14158), .ZN(
        n4200) );
  INV_X1 U2058 ( .A(n14101), .ZN(n14171) );
  NOR2_X1 U2059 ( .A1(n14257), .A2(N274), .ZN(n14067) );
  NOR2_X1 U2060 ( .A1(n14263), .A2(N273), .ZN(n14253) );
  NOR2_X1 U2061 ( .A1(n14262), .A2(N273), .ZN(n14254) );
  OAI21_X1 U2062 ( .B1(n14005), .B2(n14006), .A(n18039), .ZN(n14000) );
  OAI221_X1 U2063 ( .B1(n14220), .B2(n12413), .C1(n14058), .C2(n12415), .A(
        n18036), .ZN(n4273) );
  OAI221_X1 U2064 ( .B1(n14217), .B2(n12413), .C1(n12415), .C2(n14228), .A(
        n18035), .ZN(n4270) );
  OAI221_X1 U2065 ( .B1(n14213), .B2(n12413), .C1(n12415), .C2(n14226), .A(
        n18035), .ZN(n4267) );
  OAI221_X1 U2066 ( .B1(n12412), .B2(n12413), .C1(n12414), .C2(n12415), .A(
        n18035), .ZN(n10511) );
  OAI221_X1 U2067 ( .B1(n14214), .B2(n14220), .C1(n12415), .C2(n14221), .A(
        n18035), .ZN(n4259) );
  OAI221_X1 U2068 ( .B1(n14214), .B2(n12412), .C1(n12415), .C2(n14222), .A(
        n18035), .ZN(n4262) );
  OAI221_X1 U2069 ( .B1(n14214), .B2(n14217), .C1(n12415), .C2(n14218), .A(
        n18035), .ZN(n4256) );
  OAI221_X1 U2070 ( .B1(n14213), .B2(n14214), .C1(n12415), .C2(n14215), .A(
        n18035), .ZN(n4251) );
  NOR2_X1 U2071 ( .A1(N275), .A2(N274), .ZN(n14260) );
  NAND4_X1 U2072 ( .A1(N9922), .A2(N9924), .A3(n14174), .A4(n14020), .ZN(
        n14099) );
  NOR2_X1 U2073 ( .A1(N9641), .A2(N9909), .ZN(n14133) );
  INV_X1 U2074 ( .A(N9925), .ZN(n14205) );
  AOI22_X1 U2075 ( .A1(n14170), .A2(n14180), .B1(n14176), .B2(n14092), .ZN(
        n4209) );
  AOI22_X1 U2076 ( .A1(n14204), .A2(n14170), .B1(n14197), .B2(n14092), .ZN(
        n4237) );
  NAND2_X1 U2077 ( .A1(N9925), .A2(n14138), .ZN(n14134) );
  AOI21_X1 U2078 ( .B1(n14105), .B2(n14088), .A(n14200), .ZN(n4228) );
  AND3_X1 U2079 ( .A1(n14147), .A2(n14140), .A3(n14179), .ZN(n14200) );
  AND3_X1 U2080 ( .A1(N46302), .A2(n13962), .A3(N46303), .ZN(n13957) );
  AOI21_X1 U2081 ( .B1(n14103), .B2(n14105), .A(n14199), .ZN(n4230) );
  AND3_X1 U2082 ( .A1(n14194), .A2(n14140), .A3(n14147), .ZN(n14199) );
  AND3_X1 U2083 ( .A1(n12481), .A2(n12499), .A3(N45789), .ZN(n12463) );
  NAND2_X1 U2084 ( .A1(n13998), .A2(n13997), .ZN(n14007) );
  NAND2_X1 U2085 ( .A1(n14091), .A2(N9925), .ZN(n14118) );
  NAND2_X1 U2086 ( .A1(n14176), .A2(N9925), .ZN(n14167) );
  NAND2_X1 U2087 ( .A1(n14151), .A2(N9925), .ZN(n14121) );
  NOR3_X1 U2088 ( .A1(n16414), .A2(n13981), .A3(n13983), .ZN(n13987) );
  NOR3_X1 U2089 ( .A1(n16666), .A2(n12500), .A3(n12502), .ZN(n12506) );
  AOI21_X1 U2090 ( .B1(n14085), .B2(n14104), .A(n14127), .ZN(n4159) );
  AND3_X1 U2091 ( .A1(n14128), .A2(n14129), .A3(n14130), .ZN(n14127) );
  AOI21_X1 U2092 ( .B1(n14085), .B2(n14094), .A(n14132), .ZN(n4157) );
  AND3_X1 U2093 ( .A1(n14128), .A2(n14133), .A3(n14130), .ZN(n14132) );
  AOI21_X1 U2094 ( .B1(n14176), .B2(n14152), .A(n14177), .ZN(n4211) );
  AND3_X1 U2095 ( .A1(n14178), .A2(n14179), .A3(n14180), .ZN(n14177) );
  AOI21_X1 U2096 ( .B1(n14197), .B2(n14152), .A(n14206), .ZN(n4235) );
  AND3_X1 U2097 ( .A1(n14178), .A2(n14179), .A3(n14204), .ZN(n14206) );
  AND3_X1 U2098 ( .A1(n13962), .A2(n13980), .A3(N46303), .ZN(n13944) );
  AND3_X1 U2099 ( .A1(n12481), .A2(n12482), .A3(N45788), .ZN(n12444) );
  AND3_X1 U2100 ( .A1(N45788), .A2(n12481), .A3(N45789), .ZN(n12474) );
  INV_X1 U2101 ( .A(n14165), .ZN(n4191) );
  OAI22_X1 U2102 ( .A1(n14163), .A2(n14159), .B1(n14164), .B2(n14160), .ZN(
        n14165) );
  NOR2_X1 U2103 ( .A1(n14020), .A2(n14178), .ZN(n14147) );
  NOR2_X1 U2104 ( .A1(N9921), .A2(N9923), .ZN(n14138) );
  NAND2_X1 U2105 ( .A1(datain[30]), .A2(n18039), .ZN(n4058) );
  NAND2_X1 U2106 ( .A1(datain[31]), .A2(n18039), .ZN(n10510) );
  NAND2_X1 U2107 ( .A1(datain[24]), .A2(n18038), .ZN(n5040) );
  NAND2_X1 U2108 ( .A1(datain[26]), .A2(n18038), .ZN(n4791) );
  NAND2_X1 U2109 ( .A1(datain[28]), .A2(n18038), .ZN(n4533) );
  NAND2_X1 U2110 ( .A1(datain[7]), .A2(n18033), .ZN(n7537) );
  NAND2_X1 U2111 ( .A1(datain[8]), .A2(n18037), .ZN(n7428) );
  NAND2_X1 U2112 ( .A1(datain[9]), .A2(n18034), .ZN(n7319) );
  NAND2_X1 U2113 ( .A1(datain[10]), .A2(n18033), .ZN(n7205) );
  NAND2_X1 U2114 ( .A1(datain[11]), .A2(n18034), .ZN(n7096) );
  NAND2_X1 U2115 ( .A1(datain[12]), .A2(n18033), .ZN(n6987) );
  NAND2_X1 U2116 ( .A1(datain[13]), .A2(n18037), .ZN(n6878) );
  NAND2_X1 U2117 ( .A1(datain[14]), .A2(n18034), .ZN(n6769) );
  NAND2_X1 U2118 ( .A1(datain[15]), .A2(n18033), .ZN(n6635) );
  NAND2_X1 U2119 ( .A1(datain[16]), .A2(n18037), .ZN(n6448) );
  NAND2_X1 U2120 ( .A1(datain[17]), .A2(n18037), .ZN(n6261) );
  NAND2_X1 U2121 ( .A1(datain[18]), .A2(n18038), .ZN(n6076) );
  NAND2_X1 U2122 ( .A1(datain[19]), .A2(n18037), .ZN(n5889) );
  NAND2_X1 U2123 ( .A1(datain[20]), .A2(n18034), .ZN(n5717) );
  NAND2_X1 U2124 ( .A1(datain[21]), .A2(n18033), .ZN(n5530) );
  NAND2_X1 U2125 ( .A1(datain[22]), .A2(n18034), .ZN(n5343) );
  NAND2_X1 U2126 ( .A1(datain[23]), .A2(n18038), .ZN(n5157) );
  NAND2_X1 U2127 ( .A1(datain[25]), .A2(n18037), .ZN(n4924) );
  NAND2_X1 U2128 ( .A1(datain[27]), .A2(n18034), .ZN(n4664) );
  NAND2_X1 U2129 ( .A1(datain[29]), .A2(n18038), .ZN(n4278) );
  AND3_X1 U2130 ( .A1(n13962), .A2(n13963), .A3(N46302), .ZN(n13921) );
  OAI221_X1 U2131 ( .B1(n17836), .B2(n14296), .C1(n17854), .C2(n16461), .A(
        n18034), .ZN(n8030) );
  OAI221_X1 U2132 ( .B1(n17858), .B2(n14997), .C1(n17876), .C2(n16461), .A(
        n18034), .ZN(n8031) );
  OAI221_X1 U2133 ( .B1(n17880), .B2(n15361), .C1(n17898), .C2(n16461), .A(
        n18034), .ZN(n8032) );
  OAI221_X1 U2134 ( .B1(n17902), .B2(n14635), .C1(n17920), .C2(n16461), .A(
        n18034), .ZN(n8033) );
  OAI221_X1 U2135 ( .B1(n17923), .B2(n15353), .C1(n17941), .C2(n16461), .A(
        n18034), .ZN(n8034) );
  OAI221_X1 U2136 ( .B1(n17944), .B2(n14863), .C1(n17962), .C2(n16461), .A(
        n18034), .ZN(n8035) );
  OAI221_X1 U2137 ( .B1(n17965), .B2(n15240), .C1(n17983), .C2(n16461), .A(
        n18034), .ZN(n8036) );
  OAI221_X1 U2138 ( .B1(n17836), .B2(n14297), .C1(n17854), .C2(n16714), .A(
        n18036), .ZN(n8158) );
  OAI221_X1 U2139 ( .B1(n17858), .B2(n14998), .C1(n17875), .C2(n16714), .A(
        n18036), .ZN(n8159) );
  OAI221_X1 U2140 ( .B1(n17880), .B2(n15362), .C1(n17897), .C2(n16714), .A(
        n18036), .ZN(n8160) );
  OAI221_X1 U2141 ( .B1(n17902), .B2(n14636), .C1(n17920), .C2(n16714), .A(
        n18036), .ZN(n8161) );
  OAI221_X1 U2142 ( .B1(n17923), .B2(n15354), .C1(n17940), .C2(n16714), .A(
        n18037), .ZN(n8162) );
  OAI221_X1 U2143 ( .B1(n17944), .B2(n14864), .C1(n17962), .C2(n16714), .A(
        n18033), .ZN(n8163) );
  OAI221_X1 U2144 ( .B1(n17965), .B2(n15241), .C1(n17983), .C2(n16714), .A(
        n18034), .ZN(n8164) );
  OAI221_X1 U2145 ( .B1(n17836), .B2(n14298), .C1(n17853), .C2(n16723), .A(
        n18037), .ZN(n8230) );
  OAI221_X1 U2146 ( .B1(n17858), .B2(n14999), .C1(n17876), .C2(n16723), .A(
        n18034), .ZN(n8231) );
  OAI221_X1 U2147 ( .B1(n17880), .B2(n15364), .C1(n17898), .C2(n16723), .A(
        n18037), .ZN(n8232) );
  OAI221_X1 U2148 ( .B1(n17902), .B2(n14637), .C1(n17919), .C2(n16723), .A(
        n18038), .ZN(n8233) );
  OAI221_X1 U2149 ( .B1(n17923), .B2(n15355), .C1(n17941), .C2(n16723), .A(
        n18037), .ZN(n8234) );
  OAI221_X1 U2150 ( .B1(n17944), .B2(n14865), .C1(n17961), .C2(n16723), .A(
        n18038), .ZN(n8235) );
  OAI221_X1 U2151 ( .B1(n17965), .B2(n15242), .C1(n17982), .C2(n16723), .A(
        n18034), .ZN(n8236) );
  OAI221_X1 U2152 ( .B1(n17170), .B2(n12016), .C1(n17179), .C2(n16460), .A(
        n18033), .ZN(n8050) );
  OAI221_X1 U2153 ( .B1(n17182), .B2(n12340), .C1(n17190), .C2(n16460), .A(
        n18033), .ZN(n8051) );
  OAI221_X1 U2154 ( .B1(n17192), .B2(n14282), .C1(n17200), .C2(n16460), .A(
        n18033), .ZN(n8052) );
  OAI221_X1 U2155 ( .B1(n16944), .B2(n11905), .C1(n16953), .C2(n16461), .A(
        n18034), .ZN(n8039) );
  OAI221_X1 U2156 ( .B1(n16956), .B2(n14641), .C1(n16964), .C2(n16460), .A(
        n18033), .ZN(n8040) );
  OAI221_X1 U2157 ( .B1(n16966), .B2(n15356), .C1(n16974), .C2(n16460), .A(
        n18033), .ZN(n8041) );
  OAI221_X1 U2158 ( .B1(n16976), .B2(n14861), .C1(n16984), .C2(n16460), .A(
        n18033), .ZN(n8042) );
  OAI221_X1 U2159 ( .B1(n16999), .B2(n14292), .C1(n17007), .C2(n16460), .A(
        n18033), .ZN(n8044) );
  OAI221_X1 U2160 ( .B1(n17137), .B2(n14638), .C1(n17145), .C2(n16460), .A(
        n18033), .ZN(n8047) );
  OAI221_X1 U2161 ( .B1(n17160), .B2(n14989), .C1(n17168), .C2(n16460), .A(
        n18033), .ZN(n8049) );
  OAI221_X1 U2162 ( .B1(n16877), .B2(n14866), .C1(n16885), .C2(n16713), .A(
        n18037), .ZN(n8169) );
  OAI221_X1 U2163 ( .B1(n16887), .B2(n15351), .C1(n16895), .C2(n16713), .A(
        n18038), .ZN(n8170) );
  OAI221_X1 U2164 ( .B1(n16910), .B2(n14294), .C1(n16918), .C2(n16713), .A(
        n18034), .ZN(n8172) );
  OAI221_X1 U2165 ( .B1(n4382), .B2(n14639), .C1(n17145), .C2(n16713), .A(
        n18038), .ZN(n8175) );
  OAI221_X1 U2166 ( .B1(n4376), .B2(n14990), .C1(n17168), .C2(n16713), .A(
        n18033), .ZN(n8177) );
  OAI221_X1 U2167 ( .B1(n4373), .B2(n12017), .C1(n17179), .C2(n16713), .A(
        n18037), .ZN(n8178) );
  OAI221_X1 U2168 ( .B1(n4370), .B2(n12341), .C1(n17190), .C2(n16713), .A(
        n18037), .ZN(n8179) );
  OAI221_X1 U2169 ( .B1(n4367), .B2(n14283), .C1(n17200), .C2(n16713), .A(
        n18037), .ZN(n8180) );
  OAI221_X1 U2170 ( .B1(n16877), .B2(n14867), .C1(n16885), .C2(n16722), .A(
        n18038), .ZN(n8241) );
  OAI221_X1 U2171 ( .B1(n16887), .B2(n15352), .C1(n16895), .C2(n16722), .A(
        n18037), .ZN(n8242) );
  OAI221_X1 U2172 ( .B1(n16910), .B2(n14295), .C1(n16918), .C2(n16722), .A(
        n18038), .ZN(n8244) );
  OAI221_X1 U2173 ( .B1(n16944), .B2(n11906), .C1(n16953), .C2(n16722), .A(
        n18033), .ZN(n8247) );
  OAI221_X1 U2174 ( .B1(n16956), .B2(n14642), .C1(n16964), .C2(n16722), .A(
        n18038), .ZN(n8248) );
  OAI221_X1 U2175 ( .B1(n16966), .B2(n15357), .C1(n16974), .C2(n16722), .A(
        n18037), .ZN(n8249) );
  OAI221_X1 U2176 ( .B1(n4429), .B2(n14862), .C1(n16984), .C2(n16722), .A(
        n18038), .ZN(n8250) );
  OAI221_X1 U2177 ( .B1(n16999), .B2(n14293), .C1(n17007), .C2(n16722), .A(
        n18034), .ZN(n8252) );
  OAI22_X1 U2178 ( .A1(n16681), .A2(n14960), .B1(n16678), .B2(n14284), .ZN(
        n12419) );
  OAI22_X1 U2179 ( .A1(n16681), .A2(n14961), .B1(n16678), .B2(n14285), .ZN(
        n12262) );
  OAI22_X1 U2180 ( .A1(n16681), .A2(n14962), .B1(n16678), .B2(n14286), .ZN(
        n12109) );
  OAI22_X1 U2181 ( .A1(n16681), .A2(n14980), .B1(n16678), .B2(n14287), .ZN(
        n11956) );
  OAI22_X1 U2182 ( .A1(n14051), .A2(n16679), .B1(n16678), .B2(n14856), .ZN(
        n10518) );
  OAI22_X1 U2183 ( .A1(n17729), .A2(n15620), .B1(n17726), .B2(n12332), .ZN(
        n5295) );
  OAI22_X1 U2184 ( .A1(n17717), .A2(n15631), .B1(n17714), .B2(n11867), .ZN(
        n5303) );
  OAI22_X1 U2185 ( .A1(n17729), .A2(n15621), .B1(n17726), .B2(n12333), .ZN(
        n5129) );
  OAI22_X1 U2186 ( .A1(n17717), .A2(n15632), .B1(n17714), .B2(n11869), .ZN(
        n5134) );
  OAI22_X1 U2187 ( .A1(n17729), .A2(n15622), .B1(n17726), .B2(n12334), .ZN(
        n5013) );
  OAI22_X1 U2188 ( .A1(n17717), .A2(n15633), .B1(n17714), .B2(n11870), .ZN(
        n5020) );
  OAI22_X1 U2189 ( .A1(n17729), .A2(n15623), .B1(n17726), .B2(n12335), .ZN(
        n4891) );
  OAI22_X1 U2190 ( .A1(n17717), .A2(n15634), .B1(n17714), .B2(n11871), .ZN(
        n4900) );
  OAI22_X1 U2191 ( .A1(n17729), .A2(n15624), .B1(n17726), .B2(n12336), .ZN(
        n4764) );
  OAI22_X1 U2192 ( .A1(n17717), .A2(n15635), .B1(n17714), .B2(n11872), .ZN(
        n4771) );
  OAI22_X1 U2193 ( .A1(n17729), .A2(n15625), .B1(n17726), .B2(n12337), .ZN(
        n4633) );
  OAI22_X1 U2194 ( .A1(n17717), .A2(n15636), .B1(n17714), .B2(n11873), .ZN(
        n4638) );
  OAI22_X1 U2195 ( .A1(n17729), .A2(n15614), .B1(n17726), .B2(n12339), .ZN(
        n4506) );
  OAI22_X1 U2196 ( .A1(n17717), .A2(n15615), .B1(n17714), .B2(n11861), .ZN(
        n4511) );
  OAI22_X1 U2197 ( .A1(n17729), .A2(n15278), .B1(n17726), .B2(n12163), .ZN(
        n4172) );
  OAI22_X1 U2198 ( .A1(n17717), .A2(n15279), .B1(n17714), .B2(n11498), .ZN(
        n4183) );
  OAI22_X1 U2199 ( .A1(n16333), .A2(n15060), .B1(n16330), .B2(n12165), .ZN(
        n12913) );
  OAI22_X1 U2200 ( .A1(n16321), .A2(n15176), .B1(n16318), .B2(n14403), .ZN(
        n12914) );
  OAI22_X1 U2201 ( .A1(n16345), .A2(n12333), .B1(n16342), .B2(n11869), .ZN(
        n12912) );
  OAI22_X1 U2202 ( .A1(n16393), .A2(n14825), .B1(n16390), .B2(n11875), .ZN(
        n12904) );
  OAI22_X1 U2203 ( .A1(n16381), .A2(n15396), .B1(n16378), .B2(n14414), .ZN(
        n12905) );
  OAI22_X1 U2204 ( .A1(n16333), .A2(n15061), .B1(n16330), .B2(n12166), .ZN(
        n12871) );
  OAI22_X1 U2205 ( .A1(n16321), .A2(n15177), .B1(n16318), .B2(n14404), .ZN(
        n12872) );
  OAI22_X1 U2206 ( .A1(n16345), .A2(n12334), .B1(n16342), .B2(n11870), .ZN(
        n12870) );
  OAI22_X1 U2207 ( .A1(n16393), .A2(n14826), .B1(n16390), .B2(n11876), .ZN(
        n12862) );
  OAI22_X1 U2208 ( .A1(n16381), .A2(n15397), .B1(n16378), .B2(n14415), .ZN(
        n12863) );
  OAI22_X1 U2209 ( .A1(n16333), .A2(n15062), .B1(n16330), .B2(n12167), .ZN(
        n12829) );
  OAI22_X1 U2210 ( .A1(n16321), .A2(n15178), .B1(n16318), .B2(n14405), .ZN(
        n12830) );
  OAI22_X1 U2211 ( .A1(n16345), .A2(n12335), .B1(n16342), .B2(n11871), .ZN(
        n12828) );
  OAI22_X1 U2212 ( .A1(n16393), .A2(n14827), .B1(n16390), .B2(n11877), .ZN(
        n12820) );
  OAI22_X1 U2213 ( .A1(n16381), .A2(n15398), .B1(n16378), .B2(n14416), .ZN(
        n12821) );
  OAI22_X1 U2214 ( .A1(n16333), .A2(n15063), .B1(n16330), .B2(n12168), .ZN(
        n12787) );
  OAI22_X1 U2215 ( .A1(n16321), .A2(n15179), .B1(n16318), .B2(n14406), .ZN(
        n12788) );
  OAI22_X1 U2216 ( .A1(n16345), .A2(n12336), .B1(n16342), .B2(n11872), .ZN(
        n12786) );
  OAI22_X1 U2217 ( .A1(n16393), .A2(n14828), .B1(n16390), .B2(n11878), .ZN(
        n12778) );
  OAI22_X1 U2218 ( .A1(n16381), .A2(n15399), .B1(n16378), .B2(n14417), .ZN(
        n12779) );
  OAI22_X1 U2219 ( .A1(n16333), .A2(n15064), .B1(n16330), .B2(n12169), .ZN(
        n12745) );
  OAI22_X1 U2220 ( .A1(n16321), .A2(n15180), .B1(n16318), .B2(n14407), .ZN(
        n12746) );
  OAI22_X1 U2221 ( .A1(n16345), .A2(n12337), .B1(n16342), .B2(n11873), .ZN(
        n12744) );
  OAI22_X1 U2222 ( .A1(n16393), .A2(n14829), .B1(n16390), .B2(n11879), .ZN(
        n12736) );
  OAI22_X1 U2223 ( .A1(n16381), .A2(n15400), .B1(n16378), .B2(n14418), .ZN(
        n12737) );
  OAI22_X1 U2224 ( .A1(n16333), .A2(n15054), .B1(n16330), .B2(n12170), .ZN(
        n12703) );
  OAI22_X1 U2225 ( .A1(n16321), .A2(n15169), .B1(n16318), .B2(n14396), .ZN(
        n12704) );
  OAI22_X1 U2226 ( .A1(n16345), .A2(n12339), .B1(n16342), .B2(n11861), .ZN(
        n12702) );
  OAI22_X1 U2227 ( .A1(n16393), .A2(n14830), .B1(n16390), .B2(n11880), .ZN(
        n12694) );
  OAI22_X1 U2228 ( .A1(n16381), .A2(n15390), .B1(n16378), .B2(n14397), .ZN(
        n12695) );
  OAI22_X1 U2229 ( .A1(n16333), .A2(n14869), .B1(n16330), .B2(n12160), .ZN(
        n12660) );
  OAI22_X1 U2230 ( .A1(n16321), .A2(n14872), .B1(n16318), .B2(n14056), .ZN(
        n12661) );
  OAI22_X1 U2231 ( .A1(n16345), .A2(n12163), .B1(n16342), .B2(n11498), .ZN(
        n12659) );
  OAI22_X1 U2232 ( .A1(n16393), .A2(n14822), .B1(n16390), .B2(n11541), .ZN(
        n12650) );
  OAI22_X1 U2233 ( .A1(n16381), .A2(n15273), .B1(n16378), .B2(n14057), .ZN(
        n12651) );
  OAI22_X1 U2234 ( .A1(n16333), .A2(n15041), .B1(n16330), .B2(n12194), .ZN(
        n12574) );
  OAI22_X1 U2235 ( .A1(n16321), .A2(n15156), .B1(n16318), .B2(n14370), .ZN(
        n12579) );
  OAI22_X1 U2236 ( .A1(n16345), .A2(n12314), .B1(n16342), .B2(n11845), .ZN(
        n12569) );
  OAI22_X1 U2237 ( .A1(n16393), .A2(n14853), .B1(n16390), .B2(n11903), .ZN(
        n12544) );
  OAI22_X1 U2238 ( .A1(n16381), .A2(n15377), .B1(n16378), .B2(n14371), .ZN(
        n12549) );
  OAI22_X1 U2239 ( .A1(n16585), .A2(n15176), .B1(n16582), .B2(n14403), .ZN(
        n10963) );
  OAI22_X1 U2240 ( .A1(n16573), .A2(n15060), .B1(n16570), .B2(n12165), .ZN(
        n10964) );
  OAI22_X1 U2241 ( .A1(n16597), .A2(n12333), .B1(n16594), .B2(n11869), .ZN(
        n10962) );
  OAI22_X1 U2242 ( .A1(n16633), .A2(n14825), .B1(n16630), .B2(n14414), .ZN(
        n10955) );
  OAI22_X1 U2243 ( .A1(n16645), .A2(n14599), .B1(n16642), .B2(n11875), .ZN(
        n10954) );
  OAI22_X1 U2244 ( .A1(n16585), .A2(n15177), .B1(n16582), .B2(n14404), .ZN(
        n10920) );
  OAI22_X1 U2245 ( .A1(n16573), .A2(n15061), .B1(n16570), .B2(n12166), .ZN(
        n10921) );
  OAI22_X1 U2246 ( .A1(n16597), .A2(n12334), .B1(n16594), .B2(n11870), .ZN(
        n10919) );
  OAI22_X1 U2247 ( .A1(n16633), .A2(n14826), .B1(n16630), .B2(n14415), .ZN(
        n10912) );
  OAI22_X1 U2248 ( .A1(n16645), .A2(n14600), .B1(n16642), .B2(n11876), .ZN(
        n10911) );
  OAI22_X1 U2249 ( .A1(n16585), .A2(n15178), .B1(n16582), .B2(n14405), .ZN(
        n10877) );
  OAI22_X1 U2250 ( .A1(n16573), .A2(n15062), .B1(n16570), .B2(n12167), .ZN(
        n10878) );
  OAI22_X1 U2251 ( .A1(n16597), .A2(n12335), .B1(n16594), .B2(n11871), .ZN(
        n10876) );
  OAI22_X1 U2252 ( .A1(n16633), .A2(n14827), .B1(n16630), .B2(n14416), .ZN(
        n10869) );
  OAI22_X1 U2253 ( .A1(n16645), .A2(n14601), .B1(n16642), .B2(n11877), .ZN(
        n10868) );
  OAI22_X1 U2254 ( .A1(n16585), .A2(n15179), .B1(n16582), .B2(n14406), .ZN(
        n10834) );
  OAI22_X1 U2255 ( .A1(n16573), .A2(n15063), .B1(n16570), .B2(n12168), .ZN(
        n10835) );
  OAI22_X1 U2256 ( .A1(n16597), .A2(n12336), .B1(n16594), .B2(n11872), .ZN(
        n10833) );
  OAI22_X1 U2257 ( .A1(n16633), .A2(n14828), .B1(n16630), .B2(n14417), .ZN(
        n10826) );
  OAI22_X1 U2258 ( .A1(n16645), .A2(n14602), .B1(n16642), .B2(n11878), .ZN(
        n10825) );
  OAI22_X1 U2259 ( .A1(n16585), .A2(n15180), .B1(n16582), .B2(n14407), .ZN(
        n10791) );
  OAI22_X1 U2260 ( .A1(n16573), .A2(n15064), .B1(n16570), .B2(n12169), .ZN(
        n10792) );
  OAI22_X1 U2261 ( .A1(n16597), .A2(n12337), .B1(n16594), .B2(n11873), .ZN(
        n10790) );
  OAI22_X1 U2262 ( .A1(n16633), .A2(n14829), .B1(n16630), .B2(n14418), .ZN(
        n10783) );
  OAI22_X1 U2263 ( .A1(n16645), .A2(n14603), .B1(n16642), .B2(n11879), .ZN(
        n10782) );
  OAI22_X1 U2264 ( .A1(n16585), .A2(n15169), .B1(n16582), .B2(n14396), .ZN(
        n10748) );
  OAI22_X1 U2265 ( .A1(n16573), .A2(n15054), .B1(n16570), .B2(n12170), .ZN(
        n10749) );
  OAI22_X1 U2266 ( .A1(n16597), .A2(n12339), .B1(n16594), .B2(n11861), .ZN(
        n10747) );
  OAI22_X1 U2267 ( .A1(n16633), .A2(n14830), .B1(n16630), .B2(n14397), .ZN(
        n10740) );
  OAI22_X1 U2268 ( .A1(n16645), .A2(n14604), .B1(n16642), .B2(n11880), .ZN(
        n10739) );
  OAI22_X1 U2269 ( .A1(n16585), .A2(n14872), .B1(n16582), .B2(n14056), .ZN(
        n10695) );
  OAI22_X1 U2270 ( .A1(n16573), .A2(n14869), .B1(n16570), .B2(n12160), .ZN(
        n10698) );
  OAI22_X1 U2271 ( .A1(n16597), .A2(n12163), .B1(n16594), .B2(n11498), .ZN(
        n10694) );
  OAI22_X1 U2272 ( .A1(n16633), .A2(n14822), .B1(n16630), .B2(n14057), .ZN(
        n10683) );
  OAI22_X1 U2273 ( .A1(n16645), .A2(n14299), .B1(n16642), .B2(n11541), .ZN(
        n10682) );
  OAI22_X1 U2274 ( .A1(n16585), .A2(n15156), .B1(n16582), .B2(n14370), .ZN(
        n10584) );
  OAI22_X1 U2275 ( .A1(n16573), .A2(n15041), .B1(n16570), .B2(n12194), .ZN(
        n10591) );
  OAI22_X1 U2276 ( .A1(n16597), .A2(n12314), .B1(n16594), .B2(n11845), .ZN(
        n10577) );
  OAI22_X1 U2277 ( .A1(n16633), .A2(n14853), .B1(n16630), .B2(n14371), .ZN(
        n10551) );
  OAI22_X1 U2278 ( .A1(n16645), .A2(n14627), .B1(n16642), .B2(n11903), .ZN(
        n10544) );
  OAI22_X1 U2279 ( .A1(n17765), .A2(n15420), .B1(n17762), .B2(n14505), .ZN(
        n5292) );
  OAI22_X1 U2280 ( .A1(n17753), .A2(n14049), .B1(n17750), .B2(n12040), .ZN(
        n5293) );
  OAI22_X1 U2281 ( .A1(n17681), .A2(n14568), .B1(n17678), .B2(n12015), .ZN(
        n5307) );
  OAI22_X1 U2282 ( .A1(n17705), .A2(n15654), .B1(n17702), .B2(n14663), .ZN(
        n5304) );
  OAI22_X1 U2283 ( .A1(n17765), .A2(n15421), .B1(n17762), .B2(n14471), .ZN(
        n5124) );
  OAI22_X1 U2284 ( .A1(n17753), .A2(n12349), .B1(n17750), .B2(n12041), .ZN(
        n5125) );
  OAI22_X1 U2285 ( .A1(n17681), .A2(n14540), .B1(n17678), .B2(n11907), .ZN(
        n5137) );
  OAI22_X1 U2286 ( .A1(n17705), .A2(n15655), .B1(n17702), .B2(n14664), .ZN(
        n5135) );
  OAI22_X1 U2287 ( .A1(n17765), .A2(n15422), .B1(n17762), .B2(n14472), .ZN(
        n5010) );
  OAI22_X1 U2288 ( .A1(n17753), .A2(n12350), .B1(n17750), .B2(n12042), .ZN(
        n5011) );
  OAI22_X1 U2289 ( .A1(n17681), .A2(n14541), .B1(n17678), .B2(n11945), .ZN(
        n5023) );
  OAI22_X1 U2290 ( .A1(n17705), .A2(n15656), .B1(n17702), .B2(n14665), .ZN(
        n5021) );
  OAI22_X1 U2291 ( .A1(n17765), .A2(n15423), .B1(n17762), .B2(n14473), .ZN(
        n4888) );
  OAI22_X1 U2292 ( .A1(n17753), .A2(n12351), .B1(n17750), .B2(n12043), .ZN(
        n4889) );
  OAI22_X1 U2293 ( .A1(n17681), .A2(n14542), .B1(n17678), .B2(n11946), .ZN(
        n4903) );
  OAI22_X1 U2294 ( .A1(n17705), .A2(n15657), .B1(n17702), .B2(n14666), .ZN(
        n4901) );
  OAI22_X1 U2295 ( .A1(n17765), .A2(n15424), .B1(n17762), .B2(n14474), .ZN(
        n4761) );
  OAI22_X1 U2296 ( .A1(n17753), .A2(n12352), .B1(n17750), .B2(n12044), .ZN(
        n4762) );
  OAI22_X1 U2297 ( .A1(n17681), .A2(n14543), .B1(n17678), .B2(n11947), .ZN(
        n4774) );
  OAI22_X1 U2298 ( .A1(n17705), .A2(n15658), .B1(n17702), .B2(n14667), .ZN(
        n4772) );
  OAI22_X1 U2299 ( .A1(n17765), .A2(n15425), .B1(n17762), .B2(n14475), .ZN(
        n4630) );
  OAI22_X1 U2300 ( .A1(n17753), .A2(n12353), .B1(n17750), .B2(n12045), .ZN(
        n4631) );
  OAI22_X1 U2301 ( .A1(n17681), .A2(n14544), .B1(n17678), .B2(n11948), .ZN(
        n4641) );
  OAI22_X1 U2302 ( .A1(n17705), .A2(n15659), .B1(n17702), .B2(n14668), .ZN(
        n4639) );
  OAI22_X1 U2303 ( .A1(n17765), .A2(n15426), .B1(n17762), .B2(n14476), .ZN(
        n4501) );
  OAI22_X1 U2304 ( .A1(n17753), .A2(n12354), .B1(n17750), .B2(n12046), .ZN(
        n4502) );
  OAI22_X1 U2305 ( .A1(n17681), .A2(n14545), .B1(n17678), .B2(n11949), .ZN(
        n4514) );
  OAI22_X1 U2306 ( .A1(n17705), .A2(n15660), .B1(n17702), .B2(n14644), .ZN(
        n4512) );
  OAI22_X1 U2307 ( .A1(n17765), .A2(n15272), .B1(n17762), .B2(n14065), .ZN(
        n4145) );
  OAI22_X1 U2308 ( .A1(n17753), .A2(n12197), .B1(n17750), .B2(n11904), .ZN(
        n4156) );
  OAI22_X1 U2309 ( .A1(n17681), .A2(n14279), .B1(n17678), .B2(n11670), .ZN(
        n4208) );
  OAI22_X1 U2310 ( .A1(n17705), .A2(n15316), .B1(n17702), .B2(n14633), .ZN(
        n4190) );
  NOR2_X1 U2311 ( .A1(n14209), .A2(N9921), .ZN(n14202) );
  OAI221_X1 U2312 ( .B1(n17322), .B2(n15284), .C1(n17321), .C2(n16462), .A(
        n18035), .ZN(n8014) );
  OAI221_X1 U2313 ( .B1(n17335), .B2(n11627), .C1(n17334), .C2(n16462), .A(
        n18035), .ZN(n8015) );
  OAI221_X1 U2314 ( .B1(n17348), .B2(n14994), .C1(n17347), .C2(n16462), .A(
        n18035), .ZN(n8016) );
  OAI221_X1 U2315 ( .B1(n17361), .B2(n15365), .C1(n17360), .C2(n16462), .A(
        n18035), .ZN(n8017) );
  OAI221_X1 U2316 ( .B1(n17374), .B2(n14291), .C1(n17373), .C2(n16462), .A(
        n18035), .ZN(n8018) );
  OAI221_X1 U2317 ( .B1(n17387), .B2(n14640), .C1(n17386), .C2(n16461), .A(
        n18034), .ZN(n8019) );
  OAI221_X1 U2318 ( .B1(n17400), .B2(n14288), .C1(n17399), .C2(n16461), .A(
        n18034), .ZN(n8020) );
  OAI221_X1 U2319 ( .B1(n17413), .B2(n15003), .C1(n17412), .C2(n16461), .A(
        n18034), .ZN(n8021) );
  OAI221_X1 U2320 ( .B1(n16936), .B2(n14536), .C1(n16935), .C2(n16461), .A(
        n18034), .ZN(n8038) );
  OAI221_X1 U2321 ( .B1(n17009), .B2(n14995), .C1(n17017), .C2(n16460), .A(
        n18033), .ZN(n8045) );
  OAI221_X1 U2322 ( .B1(n16693), .B2(n14868), .C1(n16692), .C2(n10285), .A(
        n18036), .ZN(n8059) );
  OAI221_X1 U2323 ( .B1(n17129), .B2(n15367), .C1(n17128), .C2(n16460), .A(
        n18033), .ZN(n8046) );
  OAI221_X1 U2324 ( .B1(n17202), .B2(n15001), .C1(n17210), .C2(n16460), .A(
        n18033), .ZN(n8053) );
  OAI221_X1 U2325 ( .B1(n17231), .B2(n15350), .C1(n17230), .C2(n16715), .A(
        n18036), .ZN(n8135) );
  OAI221_X1 U2326 ( .B1(n17244), .B2(n12195), .C1(n17243), .C2(n16715), .A(
        n18036), .ZN(n8136) );
  OAI221_X1 U2327 ( .B1(n17257), .B2(n14823), .C1(n17256), .C2(n16714), .A(
        n18036), .ZN(n8137) );
  OAI221_X1 U2328 ( .B1(n17283), .B2(n14289), .C1(n17282), .C2(n16714), .A(
        n18036), .ZN(n8139) );
  OAI221_X1 U2329 ( .B1(n17296), .B2(n14569), .C1(n17295), .C2(n16714), .A(
        n18036), .ZN(n8140) );
  OAI221_X1 U2330 ( .B1(n17309), .B2(n15366), .C1(n17308), .C2(n16714), .A(
        n18036), .ZN(n8141) );
  OAI221_X1 U2331 ( .B1(n18005), .B2(n12050), .C1(n18004), .C2(n16714), .A(
        n18034), .ZN(n8166) );
  OAI221_X1 U2332 ( .B1(n18018), .B2(n14538), .C1(n18017), .C2(n16713), .A(
        n18033), .ZN(n8167) );
  OAI221_X1 U2333 ( .B1(n16920), .B2(n15359), .C1(n16928), .C2(n16713), .A(
        n18037), .ZN(n8173) );
  OAI221_X1 U2334 ( .B1(n17129), .B2(n15368), .C1(n17127), .C2(n16713), .A(
        n18033), .ZN(n8174) );
  OAI221_X1 U2335 ( .B1(n4362), .B2(n15002), .C1(n17210), .C2(n16713), .A(
        n18038), .ZN(n8181) );
  OAI221_X1 U2336 ( .B1(n17025), .B2(n12162), .C1(n17024), .C2(n16724), .A(
        n18037), .ZN(n8190) );
  OAI221_X1 U2337 ( .B1(n17038), .B2(n14993), .C1(n17037), .C2(n16724), .A(
        n18037), .ZN(n8191) );
  OAI221_X1 U2338 ( .B1(n17051), .B2(n14290), .C1(n17050), .C2(n16724), .A(
        n18037), .ZN(n8192) );
  OAI221_X1 U2339 ( .B1(n17064), .B2(n15000), .C1(n17063), .C2(n16724), .A(
        n18038), .ZN(n8193) );
  OAI221_X1 U2340 ( .B1(n17077), .B2(n15363), .C1(n17076), .C2(n16723), .A(
        n18037), .ZN(n8194) );
  OAI221_X1 U2341 ( .B1(n17090), .B2(n15358), .C1(n17089), .C2(n16723), .A(
        n18033), .ZN(n8195) );
  OAI221_X1 U2342 ( .B1(n17103), .B2(n11584), .C1(n17102), .C2(n16723), .A(
        n18037), .ZN(n8196) );
  OAI221_X1 U2343 ( .B1(n17116), .B2(n12308), .C1(n17115), .C2(n16723), .A(
        n18033), .ZN(n8197) );
  OAI221_X1 U2344 ( .B1(n18005), .B2(n12051), .C1(n18003), .C2(n16723), .A(
        n18038), .ZN(n8238) );
  OAI221_X1 U2345 ( .B1(n18018), .B2(n14539), .C1(n18016), .C2(n16722), .A(
        n18037), .ZN(n8239) );
  OAI221_X1 U2346 ( .B1(n16920), .B2(n15360), .C1(n16928), .C2(n16722), .A(
        n18038), .ZN(n8245) );
  OAI221_X1 U2347 ( .B1(n16936), .B2(n14537), .C1(n16934), .C2(n16722), .A(
        n18038), .ZN(n8246) );
  OAI221_X1 U2348 ( .B1(n4420), .B2(n14996), .C1(n17017), .C2(n16722), .A(
        n18038), .ZN(n8253) );
  OAI221_X1 U2349 ( .B1(n17578), .B2(n14053), .C1(n17577), .C2(n10285), .A(
        n18037), .ZN(n8257) );
  OAI22_X1 U2350 ( .A1(n14983), .A2(n16429), .B1(n14273), .B2(n16426), .ZN(
        n12892) );
  OAI22_X1 U2351 ( .A1(n14984), .A2(n16429), .B1(n14274), .B2(n16426), .ZN(
        n12850) );
  OAI22_X1 U2352 ( .A1(n14985), .A2(n16429), .B1(n14275), .B2(n16426), .ZN(
        n12808) );
  OAI22_X1 U2353 ( .A1(n14986), .A2(n16429), .B1(n14276), .B2(n16426), .ZN(
        n12766) );
  OAI22_X1 U2354 ( .A1(n14987), .A2(n16429), .B1(n14277), .B2(n16426), .ZN(
        n12724) );
  OAI22_X1 U2355 ( .A1(n14988), .A2(n16429), .B1(n14278), .B2(n16426), .ZN(
        n12682) );
  OAI22_X1 U2356 ( .A1(n14860), .A2(n16429), .B1(n14052), .B2(n16426), .ZN(
        n12638) );
  OAI22_X1 U2357 ( .A1(n14051), .A2(n16429), .B1(n14856), .B2(n16426), .ZN(
        n12521) );
  OAI22_X1 U2358 ( .A1(n16681), .A2(n14963), .B1(n14071), .B2(n16678), .ZN(
        n11803) );
  OAI22_X1 U2359 ( .A1(n16681), .A2(n14964), .B1(n14212), .B2(n16678), .ZN(
        n11760) );
  OAI22_X1 U2360 ( .A1(n16680), .A2(n14868), .B1(n14053), .B2(n16678), .ZN(
        n11717) );
  OAI22_X1 U2361 ( .A1(n16331), .A2(n15037), .B1(n16328), .B2(n12171), .ZN(
        n13945) );
  OAI22_X1 U2362 ( .A1(n16319), .A2(n15152), .B1(n16316), .B2(n14359), .ZN(
        n13947) );
  OAI22_X1 U2363 ( .A1(n16343), .A2(n12309), .B1(n16340), .B2(n11713), .ZN(
        n13943) );
  OAI22_X1 U2364 ( .A1(n16391), .A2(n14831), .B1(n16388), .B2(n11881), .ZN(
        n13924) );
  OAI22_X1 U2365 ( .A1(n16379), .A2(n15373), .B1(n16376), .B2(n14362), .ZN(
        n13930) );
  OAI22_X1 U2366 ( .A1(n16331), .A2(n15035), .B1(n16328), .B2(n12172), .ZN(
        n13879) );
  OAI22_X1 U2367 ( .A1(n16319), .A2(n15153), .B1(n16316), .B2(n14363), .ZN(
        n13880) );
  OAI22_X1 U2368 ( .A1(n16343), .A2(n12310), .B1(n16340), .B2(n11756), .ZN(
        n13878) );
  OAI22_X1 U2369 ( .A1(n16391), .A2(n14832), .B1(n16388), .B2(n11882), .ZN(
        n13870) );
  OAI22_X1 U2370 ( .A1(n16379), .A2(n15371), .B1(n16376), .B2(n14360), .ZN(
        n13871) );
  OAI22_X1 U2371 ( .A1(n16331), .A2(n15036), .B1(n16328), .B2(n12173), .ZN(
        n13837) );
  OAI22_X1 U2372 ( .A1(n16319), .A2(n15151), .B1(n16316), .B2(n14361), .ZN(
        n13838) );
  OAI22_X1 U2373 ( .A1(n16343), .A2(n12311), .B1(n16340), .B2(n11799), .ZN(
        n13836) );
  OAI22_X1 U2374 ( .A1(n16391), .A2(n14833), .B1(n16388), .B2(n11883), .ZN(
        n13828) );
  OAI22_X1 U2375 ( .A1(n16379), .A2(n15372), .B1(n16376), .B2(n14364), .ZN(
        n13829) );
  OAI22_X1 U2376 ( .A1(n16331), .A2(n15038), .B1(n16328), .B2(n12174), .ZN(
        n13795) );
  OAI22_X1 U2377 ( .A1(n16319), .A2(n15154), .B1(n16316), .B2(n14365), .ZN(
        n13796) );
  OAI22_X1 U2378 ( .A1(n16343), .A2(n12312), .B1(n16340), .B2(n11842), .ZN(
        n13794) );
  OAI22_X1 U2379 ( .A1(n16391), .A2(n14834), .B1(n16388), .B2(n11627), .ZN(
        n13786) );
  OAI22_X1 U2380 ( .A1(n16379), .A2(n15374), .B1(n16376), .B2(n14366), .ZN(
        n13787) );
  OAI22_X1 U2381 ( .A1(n16331), .A2(n15039), .B1(n16328), .B2(n12175), .ZN(
        n13753) );
  OAI22_X1 U2382 ( .A1(n16319), .A2(n15155), .B1(n16316), .B2(n14367), .ZN(
        n13754) );
  OAI22_X1 U2383 ( .A1(n16343), .A2(n12313), .B1(n16340), .B2(n11844), .ZN(
        n13752) );
  OAI22_X1 U2384 ( .A1(n16391), .A2(n14823), .B1(n16388), .B2(n11884), .ZN(
        n13744) );
  OAI22_X1 U2385 ( .A1(n16379), .A2(n15350), .B1(n16376), .B2(n14289), .ZN(
        n13745) );
  OAI22_X1 U2386 ( .A1(n16331), .A2(n14993), .B1(n16328), .B2(n12162), .ZN(
        n13711) );
  OAI22_X1 U2387 ( .A1(n16319), .A2(n15000), .B1(n16316), .B2(n14290), .ZN(
        n13712) );
  OAI22_X1 U2388 ( .A1(n16343), .A2(n12308), .B1(n16340), .B2(n11584), .ZN(
        n13710) );
  OAI22_X1 U2389 ( .A1(n16391), .A2(n14835), .B1(n16388), .B2(n11885), .ZN(
        n13702) );
  OAI22_X1 U2390 ( .A1(n16379), .A2(n15375), .B1(n16376), .B2(n14368), .ZN(
        n13703) );
  OAI22_X1 U2391 ( .A1(n16331), .A2(n15040), .B1(n16328), .B2(n12176), .ZN(
        n13669) );
  OAI22_X1 U2392 ( .A1(n16319), .A2(n15157), .B1(n16316), .B2(n14369), .ZN(
        n13670) );
  OAI22_X1 U2393 ( .A1(n16343), .A2(n12315), .B1(n16340), .B2(n11846), .ZN(
        n13668) );
  OAI22_X1 U2394 ( .A1(n16391), .A2(n14836), .B1(n16388), .B2(n11886), .ZN(
        n13660) );
  OAI22_X1 U2395 ( .A1(n16379), .A2(n15376), .B1(n16376), .B2(n14372), .ZN(
        n13661) );
  OAI22_X1 U2396 ( .A1(n16331), .A2(n15042), .B1(n16328), .B2(n12177), .ZN(
        n13627) );
  OAI22_X1 U2397 ( .A1(n16319), .A2(n15158), .B1(n16316), .B2(n14373), .ZN(
        n13628) );
  OAI22_X1 U2398 ( .A1(n16343), .A2(n12316), .B1(n16340), .B2(n11847), .ZN(
        n13626) );
  OAI22_X1 U2399 ( .A1(n16391), .A2(n14837), .B1(n16388), .B2(n11887), .ZN(
        n13618) );
  OAI22_X1 U2400 ( .A1(n16379), .A2(n15378), .B1(n16376), .B2(n14374), .ZN(
        n13619) );
  OAI22_X1 U2401 ( .A1(n16331), .A2(n15043), .B1(n16328), .B2(n12178), .ZN(
        n13585) );
  OAI22_X1 U2402 ( .A1(n16319), .A2(n15159), .B1(n16316), .B2(n14375), .ZN(
        n13586) );
  OAI22_X1 U2403 ( .A1(n16343), .A2(n12317), .B1(n16340), .B2(n11849), .ZN(
        n13584) );
  OAI22_X1 U2404 ( .A1(n16391), .A2(n14838), .B1(n16388), .B2(n11888), .ZN(
        n13576) );
  OAI22_X1 U2405 ( .A1(n16379), .A2(n15379), .B1(n16376), .B2(n14376), .ZN(
        n13577) );
  OAI22_X1 U2406 ( .A1(n16331), .A2(n15044), .B1(n16328), .B2(n12179), .ZN(
        n13543) );
  OAI22_X1 U2407 ( .A1(n16319), .A2(n15160), .B1(n16316), .B2(n14377), .ZN(
        n13544) );
  OAI22_X1 U2408 ( .A1(n16343), .A2(n12318), .B1(n16340), .B2(n11850), .ZN(
        n13542) );
  OAI22_X1 U2409 ( .A1(n16391), .A2(n14839), .B1(n16388), .B2(n11889), .ZN(
        n13534) );
  OAI22_X1 U2410 ( .A1(n16379), .A2(n15380), .B1(n16376), .B2(n14378), .ZN(
        n13535) );
  OAI22_X1 U2411 ( .A1(n16331), .A2(n15045), .B1(n16328), .B2(n12180), .ZN(
        n13501) );
  OAI22_X1 U2412 ( .A1(n16319), .A2(n15161), .B1(n16316), .B2(n14379), .ZN(
        n13502) );
  OAI22_X1 U2413 ( .A1(n16343), .A2(n12319), .B1(n16340), .B2(n11851), .ZN(
        n13500) );
  OAI22_X1 U2414 ( .A1(n16391), .A2(n14840), .B1(n16388), .B2(n11890), .ZN(
        n13492) );
  OAI22_X1 U2415 ( .A1(n16379), .A2(n15381), .B1(n16376), .B2(n14380), .ZN(
        n13493) );
  OAI22_X1 U2416 ( .A1(n16331), .A2(n15046), .B1(n16328), .B2(n12181), .ZN(
        n13459) );
  OAI22_X1 U2417 ( .A1(n16319), .A2(n15162), .B1(n16316), .B2(n14381), .ZN(
        n13460) );
  OAI22_X1 U2418 ( .A1(n16343), .A2(n12320), .B1(n16340), .B2(n11852), .ZN(
        n13458) );
  OAI22_X1 U2419 ( .A1(n16391), .A2(n14841), .B1(n16388), .B2(n11891), .ZN(
        n13450) );
  OAI22_X1 U2420 ( .A1(n16379), .A2(n15382), .B1(n16376), .B2(n14382), .ZN(
        n13451) );
  OAI22_X1 U2421 ( .A1(n16332), .A2(n15047), .B1(n16329), .B2(n12182), .ZN(
        n13417) );
  OAI22_X1 U2422 ( .A1(n16320), .A2(n15163), .B1(n16317), .B2(n14383), .ZN(
        n13418) );
  OAI22_X1 U2423 ( .A1(n16344), .A2(n12321), .B1(n16341), .B2(n11854), .ZN(
        n13416) );
  OAI22_X1 U2424 ( .A1(n16392), .A2(n14842), .B1(n16389), .B2(n11892), .ZN(
        n13408) );
  OAI22_X1 U2425 ( .A1(n16380), .A2(n15383), .B1(n16377), .B2(n14384), .ZN(
        n13409) );
  OAI22_X1 U2426 ( .A1(n16332), .A2(n15048), .B1(n16329), .B2(n12183), .ZN(
        n13375) );
  OAI22_X1 U2427 ( .A1(n16320), .A2(n15164), .B1(n16317), .B2(n14385), .ZN(
        n13376) );
  OAI22_X1 U2428 ( .A1(n16344), .A2(n12322), .B1(n16341), .B2(n11855), .ZN(
        n13374) );
  OAI22_X1 U2429 ( .A1(n16392), .A2(n14843), .B1(n16389), .B2(n11893), .ZN(
        n13366) );
  OAI22_X1 U2430 ( .A1(n16380), .A2(n15384), .B1(n16377), .B2(n14386), .ZN(
        n13367) );
  OAI22_X1 U2431 ( .A1(n16332), .A2(n15049), .B1(n16329), .B2(n12185), .ZN(
        n13333) );
  OAI22_X1 U2432 ( .A1(n16320), .A2(n15165), .B1(n16317), .B2(n14387), .ZN(
        n13334) );
  OAI22_X1 U2433 ( .A1(n16344), .A2(n12323), .B1(n16341), .B2(n11856), .ZN(
        n13332) );
  OAI22_X1 U2434 ( .A1(n16392), .A2(n14844), .B1(n16389), .B2(n11894), .ZN(
        n13324) );
  OAI22_X1 U2435 ( .A1(n16380), .A2(n15385), .B1(n16377), .B2(n14388), .ZN(
        n13325) );
  OAI22_X1 U2436 ( .A1(n16332), .A2(n15050), .B1(n16329), .B2(n12186), .ZN(
        n13291) );
  OAI22_X1 U2437 ( .A1(n16320), .A2(n15166), .B1(n16317), .B2(n14389), .ZN(
        n13292) );
  OAI22_X1 U2438 ( .A1(n16344), .A2(n12324), .B1(n16341), .B2(n11857), .ZN(
        n13290) );
  OAI22_X1 U2439 ( .A1(n16392), .A2(n14845), .B1(n16389), .B2(n11895), .ZN(
        n13282) );
  OAI22_X1 U2440 ( .A1(n16380), .A2(n15386), .B1(n16377), .B2(n14390), .ZN(
        n13283) );
  OAI22_X1 U2441 ( .A1(n16332), .A2(n15051), .B1(n16329), .B2(n12187), .ZN(
        n13249) );
  OAI22_X1 U2442 ( .A1(n16320), .A2(n15167), .B1(n16317), .B2(n14391), .ZN(
        n13250) );
  OAI22_X1 U2443 ( .A1(n16344), .A2(n12325), .B1(n16341), .B2(n11858), .ZN(
        n13248) );
  OAI22_X1 U2444 ( .A1(n16392), .A2(n14846), .B1(n16389), .B2(n11896), .ZN(
        n13240) );
  OAI22_X1 U2445 ( .A1(n16380), .A2(n15387), .B1(n16377), .B2(n14392), .ZN(
        n13241) );
  OAI22_X1 U2446 ( .A1(n16332), .A2(n15052), .B1(n16329), .B2(n12188), .ZN(
        n13207) );
  OAI22_X1 U2447 ( .A1(n16320), .A2(n15168), .B1(n16317), .B2(n14393), .ZN(
        n13208) );
  OAI22_X1 U2448 ( .A1(n16344), .A2(n12326), .B1(n16341), .B2(n11860), .ZN(
        n13206) );
  OAI22_X1 U2449 ( .A1(n16392), .A2(n14847), .B1(n16389), .B2(n11897), .ZN(
        n13198) );
  OAI22_X1 U2450 ( .A1(n16380), .A2(n15388), .B1(n16377), .B2(n14394), .ZN(
        n13199) );
  OAI22_X1 U2451 ( .A1(n16332), .A2(n15053), .B1(n16329), .B2(n12189), .ZN(
        n13165) );
  OAI22_X1 U2452 ( .A1(n16320), .A2(n15170), .B1(n16317), .B2(n14395), .ZN(
        n13166) );
  OAI22_X1 U2453 ( .A1(n16344), .A2(n12327), .B1(n16341), .B2(n11862), .ZN(
        n13164) );
  OAI22_X1 U2454 ( .A1(n16392), .A2(n14848), .B1(n16389), .B2(n11898), .ZN(
        n13156) );
  OAI22_X1 U2455 ( .A1(n16380), .A2(n15389), .B1(n16377), .B2(n14408), .ZN(
        n13157) );
  OAI22_X1 U2456 ( .A1(n16332), .A2(n15055), .B1(n16329), .B2(n12190), .ZN(
        n13123) );
  OAI22_X1 U2457 ( .A1(n16320), .A2(n15171), .B1(n16317), .B2(n14398), .ZN(
        n13124) );
  OAI22_X1 U2458 ( .A1(n16344), .A2(n12328), .B1(n16341), .B2(n11863), .ZN(
        n13122) );
  OAI22_X1 U2459 ( .A1(n16392), .A2(n14849), .B1(n16389), .B2(n11899), .ZN(
        n13114) );
  OAI22_X1 U2460 ( .A1(n16380), .A2(n15391), .B1(n16377), .B2(n14409), .ZN(
        n13115) );
  OAI22_X1 U2461 ( .A1(n16332), .A2(n15056), .B1(n16329), .B2(n12191), .ZN(
        n13081) );
  OAI22_X1 U2462 ( .A1(n16320), .A2(n15172), .B1(n16317), .B2(n14399), .ZN(
        n13082) );
  OAI22_X1 U2463 ( .A1(n16344), .A2(n12329), .B1(n16341), .B2(n11864), .ZN(
        n13080) );
  OAI22_X1 U2464 ( .A1(n16392), .A2(n14850), .B1(n16389), .B2(n11900), .ZN(
        n13072) );
  OAI22_X1 U2465 ( .A1(n16380), .A2(n15392), .B1(n16377), .B2(n14410), .ZN(
        n13073) );
  OAI22_X1 U2466 ( .A1(n16332), .A2(n15057), .B1(n16329), .B2(n12192), .ZN(
        n13039) );
  OAI22_X1 U2467 ( .A1(n16320), .A2(n15173), .B1(n16317), .B2(n14400), .ZN(
        n13040) );
  OAI22_X1 U2468 ( .A1(n16344), .A2(n12330), .B1(n16341), .B2(n11865), .ZN(
        n13038) );
  OAI22_X1 U2469 ( .A1(n16392), .A2(n14851), .B1(n16389), .B2(n11901), .ZN(
        n13030) );
  OAI22_X1 U2470 ( .A1(n16380), .A2(n15393), .B1(n16377), .B2(n14411), .ZN(
        n13031) );
  OAI22_X1 U2471 ( .A1(n16332), .A2(n15058), .B1(n16329), .B2(n12193), .ZN(
        n12997) );
  OAI22_X1 U2472 ( .A1(n16320), .A2(n15174), .B1(n16317), .B2(n14401), .ZN(
        n12998) );
  OAI22_X1 U2473 ( .A1(n16344), .A2(n12331), .B1(n16341), .B2(n11866), .ZN(
        n12996) );
  OAI22_X1 U2474 ( .A1(n16392), .A2(n14852), .B1(n16389), .B2(n11902), .ZN(
        n12988) );
  OAI22_X1 U2475 ( .A1(n16380), .A2(n15394), .B1(n16377), .B2(n14412), .ZN(
        n12989) );
  OAI22_X1 U2476 ( .A1(n16332), .A2(n15059), .B1(n16329), .B2(n12164), .ZN(
        n12955) );
  OAI22_X1 U2477 ( .A1(n16320), .A2(n15175), .B1(n16317), .B2(n14402), .ZN(
        n12956) );
  OAI22_X1 U2478 ( .A1(n16344), .A2(n12332), .B1(n16341), .B2(n11867), .ZN(
        n12954) );
  OAI22_X1 U2479 ( .A1(n16392), .A2(n14824), .B1(n16389), .B2(n11874), .ZN(
        n12946) );
  OAI22_X1 U2480 ( .A1(n16380), .A2(n15395), .B1(n16377), .B2(n14413), .ZN(
        n12947) );
  OAI22_X1 U2481 ( .A1(n16583), .A2(n15152), .B1(n16580), .B2(n14359), .ZN(
        n12464) );
  OAI22_X1 U2482 ( .A1(n16571), .A2(n15037), .B1(n16568), .B2(n12171), .ZN(
        n12466) );
  OAI22_X1 U2483 ( .A1(n16595), .A2(n12309), .B1(n16592), .B2(n11713), .ZN(
        n12462) );
  OAI22_X1 U2484 ( .A1(n16631), .A2(n14831), .B1(n16628), .B2(n14362), .ZN(
        n12448) );
  OAI22_X1 U2485 ( .A1(n16643), .A2(n14605), .B1(n16640), .B2(n11881), .ZN(
        n12442) );
  OAI22_X1 U2486 ( .A1(n16583), .A2(n15153), .B1(n16580), .B2(n14363), .ZN(
        n12283) );
  OAI22_X1 U2487 ( .A1(n16571), .A2(n15035), .B1(n16568), .B2(n12172), .ZN(
        n12284) );
  OAI22_X1 U2488 ( .A1(n16595), .A2(n12310), .B1(n16592), .B2(n11756), .ZN(
        n12282) );
  OAI22_X1 U2489 ( .A1(n16631), .A2(n14832), .B1(n16628), .B2(n14360), .ZN(
        n12275) );
  OAI22_X1 U2490 ( .A1(n16643), .A2(n14606), .B1(n16640), .B2(n11882), .ZN(
        n12274) );
  OAI22_X1 U2491 ( .A1(n16583), .A2(n15151), .B1(n16580), .B2(n14361), .ZN(
        n12130) );
  OAI22_X1 U2492 ( .A1(n16571), .A2(n15036), .B1(n16568), .B2(n12173), .ZN(
        n12131) );
  OAI22_X1 U2493 ( .A1(n16595), .A2(n12311), .B1(n16592), .B2(n11799), .ZN(
        n12129) );
  OAI22_X1 U2494 ( .A1(n16631), .A2(n14833), .B1(n16628), .B2(n14364), .ZN(
        n12122) );
  OAI22_X1 U2495 ( .A1(n16643), .A2(n14607), .B1(n16640), .B2(n11883), .ZN(
        n12121) );
  OAI22_X1 U2496 ( .A1(n16583), .A2(n15154), .B1(n16580), .B2(n14365), .ZN(
        n11977) );
  OAI22_X1 U2497 ( .A1(n16571), .A2(n15038), .B1(n16568), .B2(n12174), .ZN(
        n11978) );
  OAI22_X1 U2498 ( .A1(n16595), .A2(n12312), .B1(n16592), .B2(n11842), .ZN(
        n11976) );
  OAI22_X1 U2499 ( .A1(n16631), .A2(n14834), .B1(n16628), .B2(n14366), .ZN(
        n11969) );
  OAI22_X1 U2500 ( .A1(n16643), .A2(n14608), .B1(n16640), .B2(n11627), .ZN(
        n11968) );
  OAI22_X1 U2501 ( .A1(n16583), .A2(n15155), .B1(n16580), .B2(n14367), .ZN(
        n11824) );
  OAI22_X1 U2502 ( .A1(n16571), .A2(n15039), .B1(n16568), .B2(n12175), .ZN(
        n11825) );
  OAI22_X1 U2503 ( .A1(n16595), .A2(n12313), .B1(n16592), .B2(n11844), .ZN(
        n11823) );
  OAI22_X1 U2504 ( .A1(n16631), .A2(n14823), .B1(n16628), .B2(n14289), .ZN(
        n11816) );
  OAI22_X1 U2505 ( .A1(n16643), .A2(n14569), .B1(n16640), .B2(n11884), .ZN(
        n11815) );
  OAI22_X1 U2506 ( .A1(n16583), .A2(n15000), .B1(n16580), .B2(n14290), .ZN(
        n11781) );
  OAI22_X1 U2507 ( .A1(n16571), .A2(n14993), .B1(n16568), .B2(n12162), .ZN(
        n11782) );
  OAI22_X1 U2508 ( .A1(n16595), .A2(n12308), .B1(n16592), .B2(n11584), .ZN(
        n11780) );
  OAI22_X1 U2509 ( .A1(n16631), .A2(n14835), .B1(n16628), .B2(n14368), .ZN(
        n11773) );
  OAI22_X1 U2510 ( .A1(n16643), .A2(n14609), .B1(n16640), .B2(n11885), .ZN(
        n11772) );
  OAI22_X1 U2511 ( .A1(n16583), .A2(n15157), .B1(n16580), .B2(n14369), .ZN(
        n11738) );
  OAI22_X1 U2512 ( .A1(n16571), .A2(n15040), .B1(n16568), .B2(n12176), .ZN(
        n11739) );
  OAI22_X1 U2513 ( .A1(n16595), .A2(n12315), .B1(n16592), .B2(n11846), .ZN(
        n11737) );
  OAI22_X1 U2514 ( .A1(n16631), .A2(n14836), .B1(n16628), .B2(n14372), .ZN(
        n11730) );
  OAI22_X1 U2515 ( .A1(n16643), .A2(n14610), .B1(n16640), .B2(n11886), .ZN(
        n11729) );
  OAI22_X1 U2516 ( .A1(n16583), .A2(n15158), .B1(n16580), .B2(n14373), .ZN(
        n11695) );
  OAI22_X1 U2517 ( .A1(n16571), .A2(n15042), .B1(n16568), .B2(n12177), .ZN(
        n11696) );
  OAI22_X1 U2518 ( .A1(n16595), .A2(n12316), .B1(n16592), .B2(n11847), .ZN(
        n11694) );
  OAI22_X1 U2519 ( .A1(n16631), .A2(n14837), .B1(n16628), .B2(n14374), .ZN(
        n11687) );
  OAI22_X1 U2520 ( .A1(n16643), .A2(n14611), .B1(n16640), .B2(n11887), .ZN(
        n11686) );
  OAI22_X1 U2521 ( .A1(n16583), .A2(n15159), .B1(n16580), .B2(n14375), .ZN(
        n11652) );
  OAI22_X1 U2522 ( .A1(n16571), .A2(n15043), .B1(n16568), .B2(n12178), .ZN(
        n11653) );
  OAI22_X1 U2523 ( .A1(n16595), .A2(n12317), .B1(n16592), .B2(n11849), .ZN(
        n11651) );
  OAI22_X1 U2524 ( .A1(n16631), .A2(n14838), .B1(n16628), .B2(n14376), .ZN(
        n11644) );
  OAI22_X1 U2525 ( .A1(n16643), .A2(n14612), .B1(n16640), .B2(n11888), .ZN(
        n11643) );
  OAI22_X1 U2526 ( .A1(n16583), .A2(n15160), .B1(n16580), .B2(n14377), .ZN(
        n11609) );
  OAI22_X1 U2527 ( .A1(n16571), .A2(n15044), .B1(n16568), .B2(n12179), .ZN(
        n11610) );
  OAI22_X1 U2528 ( .A1(n16595), .A2(n12318), .B1(n16592), .B2(n11850), .ZN(
        n11608) );
  OAI22_X1 U2529 ( .A1(n16631), .A2(n14839), .B1(n16628), .B2(n14378), .ZN(
        n11601) );
  OAI22_X1 U2530 ( .A1(n16643), .A2(n14613), .B1(n16640), .B2(n11889), .ZN(
        n11600) );
  OAI22_X1 U2531 ( .A1(n16583), .A2(n15161), .B1(n16580), .B2(n14379), .ZN(
        n11566) );
  OAI22_X1 U2532 ( .A1(n16571), .A2(n15045), .B1(n16568), .B2(n12180), .ZN(
        n11567) );
  OAI22_X1 U2533 ( .A1(n16595), .A2(n12319), .B1(n16592), .B2(n11851), .ZN(
        n11565) );
  OAI22_X1 U2534 ( .A1(n16631), .A2(n14840), .B1(n16628), .B2(n14380), .ZN(
        n11558) );
  OAI22_X1 U2535 ( .A1(n16643), .A2(n14614), .B1(n16640), .B2(n11890), .ZN(
        n11557) );
  OAI22_X1 U2536 ( .A1(n16583), .A2(n15162), .B1(n16580), .B2(n14381), .ZN(
        n11523) );
  OAI22_X1 U2537 ( .A1(n16571), .A2(n15046), .B1(n16568), .B2(n12181), .ZN(
        n11524) );
  OAI22_X1 U2538 ( .A1(n16595), .A2(n12320), .B1(n16592), .B2(n11852), .ZN(
        n11522) );
  OAI22_X1 U2539 ( .A1(n16631), .A2(n14841), .B1(n16628), .B2(n14382), .ZN(
        n11515) );
  OAI22_X1 U2540 ( .A1(n16643), .A2(n14615), .B1(n16640), .B2(n11891), .ZN(
        n11514) );
  OAI22_X1 U2541 ( .A1(n16584), .A2(n15163), .B1(n16581), .B2(n14383), .ZN(
        n11480) );
  OAI22_X1 U2542 ( .A1(n16572), .A2(n15047), .B1(n16569), .B2(n12182), .ZN(
        n11481) );
  OAI22_X1 U2543 ( .A1(n16596), .A2(n12321), .B1(n16593), .B2(n11854), .ZN(
        n11479) );
  OAI22_X1 U2544 ( .A1(n16632), .A2(n14842), .B1(n16629), .B2(n14384), .ZN(
        n11472) );
  OAI22_X1 U2545 ( .A1(n16644), .A2(n14616), .B1(n16641), .B2(n11892), .ZN(
        n11471) );
  OAI22_X1 U2546 ( .A1(n16584), .A2(n15164), .B1(n16581), .B2(n14385), .ZN(
        n11436) );
  OAI22_X1 U2547 ( .A1(n16572), .A2(n15048), .B1(n16569), .B2(n12183), .ZN(
        n11437) );
  OAI22_X1 U2548 ( .A1(n16596), .A2(n12322), .B1(n16593), .B2(n11855), .ZN(
        n11435) );
  OAI22_X1 U2549 ( .A1(n16632), .A2(n14843), .B1(n16629), .B2(n14386), .ZN(
        n11428) );
  OAI22_X1 U2550 ( .A1(n16644), .A2(n14617), .B1(n16641), .B2(n11893), .ZN(
        n11427) );
  OAI22_X1 U2551 ( .A1(n16584), .A2(n15165), .B1(n16581), .B2(n14387), .ZN(
        n11393) );
  OAI22_X1 U2552 ( .A1(n16572), .A2(n15049), .B1(n16569), .B2(n12185), .ZN(
        n11394) );
  OAI22_X1 U2553 ( .A1(n16596), .A2(n12323), .B1(n16593), .B2(n11856), .ZN(
        n11392) );
  OAI22_X1 U2554 ( .A1(n16632), .A2(n14844), .B1(n16629), .B2(n14388), .ZN(
        n11385) );
  OAI22_X1 U2555 ( .A1(n16644), .A2(n14618), .B1(n16641), .B2(n11894), .ZN(
        n11384) );
  OAI22_X1 U2556 ( .A1(n16584), .A2(n15166), .B1(n16581), .B2(n14389), .ZN(
        n11350) );
  OAI22_X1 U2557 ( .A1(n16572), .A2(n15050), .B1(n16569), .B2(n12186), .ZN(
        n11351) );
  OAI22_X1 U2558 ( .A1(n16596), .A2(n12324), .B1(n16593), .B2(n11857), .ZN(
        n11349) );
  OAI22_X1 U2559 ( .A1(n16632), .A2(n14845), .B1(n16629), .B2(n14390), .ZN(
        n11342) );
  OAI22_X1 U2560 ( .A1(n16644), .A2(n14619), .B1(n16641), .B2(n11895), .ZN(
        n11341) );
  OAI22_X1 U2561 ( .A1(n16584), .A2(n15167), .B1(n16581), .B2(n14391), .ZN(
        n11307) );
  OAI22_X1 U2562 ( .A1(n16572), .A2(n15051), .B1(n16569), .B2(n12187), .ZN(
        n11308) );
  OAI22_X1 U2563 ( .A1(n16596), .A2(n12325), .B1(n16593), .B2(n11858), .ZN(
        n11306) );
  OAI22_X1 U2564 ( .A1(n16632), .A2(n14846), .B1(n16629), .B2(n14392), .ZN(
        n11299) );
  OAI22_X1 U2565 ( .A1(n16644), .A2(n14620), .B1(n16641), .B2(n11896), .ZN(
        n11298) );
  OAI22_X1 U2566 ( .A1(n16584), .A2(n15168), .B1(n16581), .B2(n14393), .ZN(
        n11264) );
  OAI22_X1 U2567 ( .A1(n16572), .A2(n15052), .B1(n16569), .B2(n12188), .ZN(
        n11265) );
  OAI22_X1 U2568 ( .A1(n16596), .A2(n12326), .B1(n16593), .B2(n11860), .ZN(
        n11263) );
  OAI22_X1 U2569 ( .A1(n16632), .A2(n14847), .B1(n16629), .B2(n14394), .ZN(
        n11256) );
  OAI22_X1 U2570 ( .A1(n16644), .A2(n14621), .B1(n16641), .B2(n11897), .ZN(
        n11255) );
  OAI22_X1 U2571 ( .A1(n16584), .A2(n15170), .B1(n16581), .B2(n14395), .ZN(
        n11221) );
  OAI22_X1 U2572 ( .A1(n16572), .A2(n15053), .B1(n16569), .B2(n12189), .ZN(
        n11222) );
  OAI22_X1 U2573 ( .A1(n16596), .A2(n12327), .B1(n16593), .B2(n11862), .ZN(
        n11220) );
  OAI22_X1 U2574 ( .A1(n16632), .A2(n14848), .B1(n16629), .B2(n14408), .ZN(
        n11213) );
  OAI22_X1 U2575 ( .A1(n16644), .A2(n14622), .B1(n16641), .B2(n11898), .ZN(
        n11212) );
  OAI22_X1 U2576 ( .A1(n16584), .A2(n15171), .B1(n16581), .B2(n14398), .ZN(
        n11178) );
  OAI22_X1 U2577 ( .A1(n16572), .A2(n15055), .B1(n16569), .B2(n12190), .ZN(
        n11179) );
  OAI22_X1 U2578 ( .A1(n16596), .A2(n12328), .B1(n16593), .B2(n11863), .ZN(
        n11177) );
  OAI22_X1 U2579 ( .A1(n16632), .A2(n14849), .B1(n16629), .B2(n14409), .ZN(
        n11170) );
  OAI22_X1 U2580 ( .A1(n16644), .A2(n14623), .B1(n16641), .B2(n11899), .ZN(
        n11169) );
  OAI22_X1 U2581 ( .A1(n16584), .A2(n15172), .B1(n16581), .B2(n14399), .ZN(
        n11135) );
  OAI22_X1 U2582 ( .A1(n16572), .A2(n15056), .B1(n16569), .B2(n12191), .ZN(
        n11136) );
  OAI22_X1 U2583 ( .A1(n16596), .A2(n12329), .B1(n16593), .B2(n11864), .ZN(
        n11134) );
  OAI22_X1 U2584 ( .A1(n16632), .A2(n14850), .B1(n16629), .B2(n14410), .ZN(
        n11127) );
  OAI22_X1 U2585 ( .A1(n16644), .A2(n14624), .B1(n16641), .B2(n11900), .ZN(
        n11126) );
  OAI22_X1 U2586 ( .A1(n16584), .A2(n15173), .B1(n16581), .B2(n14400), .ZN(
        n11092) );
  OAI22_X1 U2587 ( .A1(n16572), .A2(n15057), .B1(n16569), .B2(n12192), .ZN(
        n11093) );
  OAI22_X1 U2588 ( .A1(n16596), .A2(n12330), .B1(n16593), .B2(n11865), .ZN(
        n11091) );
  OAI22_X1 U2589 ( .A1(n16632), .A2(n14851), .B1(n16629), .B2(n14411), .ZN(
        n11084) );
  OAI22_X1 U2590 ( .A1(n16644), .A2(n14625), .B1(n16641), .B2(n11901), .ZN(
        n11083) );
  OAI22_X1 U2591 ( .A1(n16584), .A2(n15174), .B1(n16581), .B2(n14401), .ZN(
        n11049) );
  OAI22_X1 U2592 ( .A1(n16572), .A2(n15058), .B1(n16569), .B2(n12193), .ZN(
        n11050) );
  OAI22_X1 U2593 ( .A1(n16596), .A2(n12331), .B1(n16593), .B2(n11866), .ZN(
        n11048) );
  OAI22_X1 U2594 ( .A1(n16632), .A2(n14852), .B1(n16629), .B2(n14412), .ZN(
        n11041) );
  OAI22_X1 U2595 ( .A1(n16644), .A2(n14626), .B1(n16641), .B2(n11902), .ZN(
        n11040) );
  OAI22_X1 U2596 ( .A1(n16584), .A2(n15175), .B1(n16581), .B2(n14402), .ZN(
        n11006) );
  OAI22_X1 U2597 ( .A1(n16572), .A2(n15059), .B1(n16569), .B2(n12164), .ZN(
        n11007) );
  OAI22_X1 U2598 ( .A1(n16596), .A2(n12332), .B1(n16593), .B2(n11867), .ZN(
        n11005) );
  OAI22_X1 U2599 ( .A1(n16632), .A2(n14824), .B1(n16629), .B2(n14413), .ZN(
        n10998) );
  OAI22_X1 U2600 ( .A1(n16644), .A2(n14598), .B1(n16641), .B2(n11874), .ZN(
        n10997) );
  OAI22_X1 U2601 ( .A1(n17727), .A2(n15575), .B1(n17724), .B2(n12309), .ZN(
        n12390) );
  OAI22_X1 U2602 ( .A1(n17763), .A2(n15369), .B1(n17760), .B2(n14484), .ZN(
        n12387) );
  OAI22_X1 U2603 ( .A1(n17751), .A2(n12356), .B1(n17748), .B2(n12018), .ZN(
        n12388) );
  OAI22_X1 U2604 ( .A1(n17679), .A2(n14547), .B1(n17676), .B2(n11951), .ZN(
        n12398) );
  OAI22_X1 U2605 ( .A1(n17715), .A2(n15576), .B1(n17712), .B2(n11713), .ZN(
        n12395) );
  OAI22_X1 U2606 ( .A1(n17703), .A2(n15574), .B1(n17700), .B2(n14669), .ZN(
        n12396) );
  OAI22_X1 U2607 ( .A1(n17727), .A2(n15577), .B1(n17724), .B2(n12310), .ZN(
        n12236) );
  OAI22_X1 U2608 ( .A1(n17763), .A2(n15370), .B1(n17760), .B2(n14485), .ZN(
        n12233) );
  OAI22_X1 U2609 ( .A1(n17751), .A2(n12358), .B1(n17748), .B2(n12019), .ZN(
        n12234) );
  OAI22_X1 U2610 ( .A1(n17679), .A2(n14548), .B1(n17676), .B2(n11952), .ZN(
        n12244) );
  OAI22_X1 U2611 ( .A1(n17715), .A2(n15580), .B1(n17712), .B2(n11756), .ZN(
        n12241) );
  OAI22_X1 U2612 ( .A1(n17703), .A2(n15661), .B1(n17700), .B2(n14645), .ZN(
        n12242) );
  OAI22_X1 U2613 ( .A1(n17727), .A2(n15586), .B1(n17724), .B2(n12311), .ZN(
        n12081) );
  OAI22_X1 U2614 ( .A1(n17763), .A2(n15401), .B1(n17760), .B2(n14486), .ZN(
        n12078) );
  OAI22_X1 U2615 ( .A1(n17751), .A2(n12360), .B1(n17748), .B2(n12020), .ZN(
        n12079) );
  OAI22_X1 U2616 ( .A1(n17679), .A2(n14549), .B1(n17676), .B2(n11995), .ZN(
        n12089) );
  OAI22_X1 U2617 ( .A1(n17715), .A2(n15581), .B1(n17712), .B2(n11799), .ZN(
        n12086) );
  OAI22_X1 U2618 ( .A1(n17703), .A2(n15578), .B1(n17700), .B2(n14643), .ZN(
        n12087) );
  OAI22_X1 U2619 ( .A1(n17727), .A2(n15587), .B1(n17724), .B2(n12312), .ZN(
        n11928) );
  OAI22_X1 U2620 ( .A1(n17763), .A2(n15402), .B1(n17760), .B2(n14487), .ZN(
        n11925) );
  OAI22_X1 U2621 ( .A1(n17751), .A2(n12340), .B1(n17748), .B2(n12016), .ZN(
        n11926) );
  OAI22_X1 U2622 ( .A1(n17679), .A2(n14536), .B1(n17676), .B2(n11905), .ZN(
        n11936) );
  OAI22_X1 U2623 ( .A1(n17715), .A2(n15582), .B1(n17712), .B2(n11842), .ZN(
        n11933) );
  OAI22_X1 U2624 ( .A1(n17703), .A2(n15361), .B1(n17700), .B2(n14635), .ZN(
        n11934) );
  OAI22_X1 U2625 ( .A1(n17727), .A2(n15588), .B1(n17724), .B2(n12313), .ZN(
        n10485) );
  OAI22_X1 U2626 ( .A1(n17763), .A2(n15351), .B1(n17760), .B2(n14294), .ZN(
        n10482) );
  OAI22_X1 U2627 ( .A1(n17751), .A2(n12341), .B1(n17748), .B2(n12017), .ZN(
        n10483) );
  OAI22_X1 U2628 ( .A1(n17679), .A2(n14550), .B1(n17676), .B2(n11997), .ZN(
        n10493) );
  OAI22_X1 U2629 ( .A1(n17715), .A2(n15583), .B1(n17712), .B2(n11844), .ZN(
        n10490) );
  OAI22_X1 U2630 ( .A1(n17703), .A2(n15362), .B1(n17700), .B2(n14636), .ZN(
        n10491) );
  OAI22_X1 U2631 ( .A1(n17727), .A2(n15363), .B1(n17724), .B2(n12308), .ZN(
        n10375) );
  OAI22_X1 U2632 ( .A1(n17763), .A2(n15352), .B1(n17760), .B2(n14295), .ZN(
        n10372) );
  OAI22_X1 U2633 ( .A1(n17751), .A2(n12364), .B1(n17748), .B2(n12021), .ZN(
        n10373) );
  OAI22_X1 U2634 ( .A1(n17679), .A2(n14537), .B1(n17676), .B2(n11906), .ZN(
        n10383) );
  OAI22_X1 U2635 ( .A1(n17715), .A2(n15584), .B1(n17712), .B2(n11584), .ZN(
        n10380) );
  OAI22_X1 U2636 ( .A1(n17703), .A2(n15364), .B1(n17700), .B2(n14637), .ZN(
        n10381) );
  OAI22_X1 U2637 ( .A1(n17727), .A2(n15589), .B1(n17724), .B2(n12315), .ZN(
        n10263) );
  OAI22_X1 U2638 ( .A1(n17763), .A2(n15403), .B1(n17760), .B2(n14488), .ZN(
        n10260) );
  OAI22_X1 U2639 ( .A1(n17751), .A2(n12366), .B1(n17748), .B2(n12022), .ZN(
        n10261) );
  OAI22_X1 U2640 ( .A1(n17679), .A2(n14551), .B1(n17676), .B2(n11998), .ZN(
        n10271) );
  OAI22_X1 U2641 ( .A1(n17715), .A2(n15579), .B1(n17712), .B2(n11846), .ZN(
        n10268) );
  OAI22_X1 U2642 ( .A1(n17703), .A2(n15637), .B1(n17700), .B2(n14646), .ZN(
        n10269) );
  OAI22_X1 U2643 ( .A1(n17727), .A2(n15591), .B1(n17724), .B2(n12316), .ZN(
        n7627) );
  OAI22_X1 U2644 ( .A1(n17763), .A2(n15404), .B1(n17760), .B2(n14489), .ZN(
        n7624) );
  OAI22_X1 U2645 ( .A1(n17751), .A2(n12368), .B1(n17748), .B2(n12023), .ZN(
        n7625) );
  OAI22_X1 U2646 ( .A1(n17679), .A2(n14552), .B1(n17676), .B2(n11999), .ZN(
        n7635) );
  OAI22_X1 U2647 ( .A1(n17715), .A2(n15592), .B1(n17712), .B2(n11847), .ZN(
        n7632) );
  OAI22_X1 U2648 ( .A1(n17703), .A2(n15638), .B1(n17700), .B2(n14647), .ZN(
        n7633) );
  OAI22_X1 U2649 ( .A1(n17727), .A2(n15593), .B1(n17724), .B2(n12317), .ZN(
        n7512) );
  OAI22_X1 U2650 ( .A1(n17763), .A2(n15405), .B1(n17760), .B2(n14490), .ZN(
        n7509) );
  OAI22_X1 U2651 ( .A1(n17751), .A2(n12407), .B1(n17748), .B2(n12024), .ZN(
        n7510) );
  OAI22_X1 U2652 ( .A1(n17679), .A2(n14553), .B1(n17676), .B2(n12000), .ZN(
        n7520) );
  OAI22_X1 U2653 ( .A1(n17715), .A2(n15594), .B1(n17712), .B2(n11849), .ZN(
        n7517) );
  OAI22_X1 U2654 ( .A1(n17703), .A2(n15639), .B1(n17700), .B2(n14648), .ZN(
        n7518) );
  OAI22_X1 U2655 ( .A1(n17727), .A2(n15595), .B1(n17724), .B2(n12318), .ZN(
        n7403) );
  OAI22_X1 U2656 ( .A1(n17763), .A2(n15406), .B1(n17760), .B2(n14491), .ZN(
        n7400) );
  OAI22_X1 U2657 ( .A1(n17751), .A2(n12409), .B1(n17748), .B2(n12025), .ZN(
        n7401) );
  OAI22_X1 U2658 ( .A1(n17679), .A2(n14554), .B1(n17676), .B2(n12001), .ZN(
        n7411) );
  OAI22_X1 U2659 ( .A1(n17715), .A2(n15596), .B1(n17712), .B2(n11850), .ZN(
        n7408) );
  OAI22_X1 U2660 ( .A1(n17703), .A2(n15640), .B1(n17700), .B2(n14649), .ZN(
        n7409) );
  OAI22_X1 U2661 ( .A1(n17727), .A2(n15597), .B1(n17724), .B2(n12319), .ZN(
        n7294) );
  OAI22_X1 U2662 ( .A1(n17763), .A2(n15407), .B1(n17760), .B2(n14492), .ZN(
        n7291) );
  OAI22_X1 U2663 ( .A1(n17751), .A2(n12411), .B1(n17748), .B2(n12026), .ZN(
        n7292) );
  OAI22_X1 U2664 ( .A1(n17679), .A2(n14555), .B1(n17676), .B2(n12002), .ZN(
        n7302) );
  OAI22_X1 U2665 ( .A1(n17715), .A2(n15598), .B1(n17712), .B2(n11851), .ZN(
        n7299) );
  OAI22_X1 U2666 ( .A1(n17703), .A2(n15641), .B1(n17700), .B2(n14650), .ZN(
        n7300) );
  OAI22_X1 U2667 ( .A1(n17728), .A2(n15599), .B1(n17725), .B2(n12320), .ZN(
        n7180) );
  OAI22_X1 U2668 ( .A1(n17764), .A2(n15408), .B1(n17761), .B2(n14493), .ZN(
        n7177) );
  OAI22_X1 U2669 ( .A1(n17752), .A2(n12600), .B1(n17749), .B2(n12027), .ZN(
        n7178) );
  OAI22_X1 U2670 ( .A1(n17680), .A2(n14556), .B1(n17677), .B2(n12003), .ZN(
        n7188) );
  OAI22_X1 U2671 ( .A1(n17716), .A2(n15600), .B1(n17713), .B2(n11852), .ZN(
        n7185) );
  OAI22_X1 U2672 ( .A1(n17704), .A2(n15642), .B1(n17701), .B2(n14651), .ZN(
        n7186) );
  OAI22_X1 U2673 ( .A1(n17728), .A2(n15601), .B1(n17725), .B2(n12321), .ZN(
        n7071) );
  OAI22_X1 U2674 ( .A1(n17764), .A2(n15409), .B1(n17761), .B2(n14494), .ZN(
        n7068) );
  OAI22_X1 U2675 ( .A1(n17752), .A2(n12652), .B1(n17749), .B2(n12028), .ZN(
        n7069) );
  OAI22_X1 U2676 ( .A1(n17680), .A2(n14557), .B1(n17677), .B2(n12004), .ZN(
        n7079) );
  OAI22_X1 U2677 ( .A1(n17716), .A2(n15602), .B1(n17713), .B2(n11854), .ZN(
        n7076) );
  OAI22_X1 U2678 ( .A1(n17704), .A2(n15643), .B1(n17701), .B2(n14652), .ZN(
        n7077) );
  OAI22_X1 U2679 ( .A1(n17728), .A2(n15603), .B1(n17725), .B2(n12322), .ZN(
        n6962) );
  OAI22_X1 U2680 ( .A1(n17764), .A2(n15410), .B1(n17761), .B2(n14495), .ZN(
        n6959) );
  OAI22_X1 U2681 ( .A1(n17752), .A2(n13996), .B1(n17749), .B2(n12030), .ZN(
        n6960) );
  OAI22_X1 U2682 ( .A1(n17680), .A2(n14558), .B1(n17677), .B2(n12005), .ZN(
        n6970) );
  OAI22_X1 U2683 ( .A1(n17716), .A2(n15604), .B1(n17713), .B2(n11855), .ZN(
        n6967) );
  OAI22_X1 U2684 ( .A1(n17704), .A2(n15644), .B1(n17701), .B2(n14653), .ZN(
        n6968) );
  OAI22_X1 U2685 ( .A1(n17728), .A2(n15605), .B1(n17725), .B2(n12323), .ZN(
        n6853) );
  OAI22_X1 U2686 ( .A1(n17764), .A2(n15411), .B1(n17761), .B2(n14496), .ZN(
        n6850) );
  OAI22_X1 U2687 ( .A1(n17752), .A2(n14008), .B1(n17749), .B2(n12031), .ZN(
        n6851) );
  OAI22_X1 U2688 ( .A1(n17680), .A2(n14559), .B1(n17677), .B2(n12006), .ZN(
        n6861) );
  OAI22_X1 U2689 ( .A1(n17716), .A2(n15606), .B1(n17713), .B2(n11856), .ZN(
        n6858) );
  OAI22_X1 U2690 ( .A1(n17704), .A2(n15645), .B1(n17701), .B2(n14654), .ZN(
        n6859) );
  OAI22_X1 U2691 ( .A1(n17728), .A2(n15607), .B1(n17725), .B2(n12324), .ZN(
        n6744) );
  OAI22_X1 U2692 ( .A1(n17764), .A2(n15412), .B1(n17761), .B2(n14497), .ZN(
        n6741) );
  OAI22_X1 U2693 ( .A1(n17752), .A2(n14015), .B1(n17749), .B2(n12032), .ZN(
        n6742) );
  OAI22_X1 U2694 ( .A1(n17680), .A2(n14560), .B1(n17677), .B2(n12007), .ZN(
        n6752) );
  OAI22_X1 U2695 ( .A1(n17716), .A2(n15608), .B1(n17713), .B2(n11857), .ZN(
        n6749) );
  OAI22_X1 U2696 ( .A1(n17704), .A2(n15646), .B1(n17701), .B2(n14655), .ZN(
        n6750) );
  OAI22_X1 U2697 ( .A1(n17728), .A2(n15609), .B1(n17725), .B2(n12325), .ZN(
        n6601) );
  OAI22_X1 U2698 ( .A1(n17764), .A2(n15413), .B1(n17761), .B2(n14498), .ZN(
        n6598) );
  OAI22_X1 U2699 ( .A1(n17752), .A2(n14035), .B1(n17749), .B2(n12033), .ZN(
        n6599) );
  OAI22_X1 U2700 ( .A1(n17680), .A2(n14561), .B1(n17677), .B2(n12008), .ZN(
        n6610) );
  OAI22_X1 U2701 ( .A1(n17716), .A2(n15610), .B1(n17713), .B2(n11858), .ZN(
        n6606) );
  OAI22_X1 U2702 ( .A1(n17704), .A2(n15647), .B1(n17701), .B2(n14656), .ZN(
        n6607) );
  OAI22_X1 U2703 ( .A1(n17728), .A2(n15611), .B1(n17725), .B2(n12326), .ZN(
        n6414) );
  OAI22_X1 U2704 ( .A1(n17764), .A2(n15414), .B1(n17761), .B2(n14499), .ZN(
        n6411) );
  OAI22_X1 U2705 ( .A1(n17752), .A2(n14037), .B1(n17749), .B2(n12034), .ZN(
        n6412) );
  OAI22_X1 U2706 ( .A1(n17680), .A2(n14562), .B1(n17677), .B2(n12009), .ZN(
        n6425) );
  OAI22_X1 U2707 ( .A1(n17716), .A2(n15612), .B1(n17713), .B2(n11860), .ZN(
        n6420) );
  OAI22_X1 U2708 ( .A1(n17704), .A2(n15648), .B1(n17701), .B2(n14657), .ZN(
        n6421) );
  OAI22_X1 U2709 ( .A1(n17728), .A2(n15613), .B1(n17725), .B2(n12327), .ZN(
        n6227) );
  OAI22_X1 U2710 ( .A1(n17764), .A2(n15415), .B1(n17761), .B2(n14500), .ZN(
        n6224) );
  OAI22_X1 U2711 ( .A1(n17752), .A2(n14039), .B1(n17749), .B2(n12035), .ZN(
        n6225) );
  OAI22_X1 U2712 ( .A1(n17680), .A2(n14563), .B1(n17677), .B2(n12010), .ZN(
        n6238) );
  OAI22_X1 U2713 ( .A1(n17716), .A2(n15626), .B1(n17713), .B2(n11862), .ZN(
        n6234) );
  OAI22_X1 U2714 ( .A1(n17704), .A2(n15649), .B1(n17701), .B2(n14658), .ZN(
        n6236) );
  OAI22_X1 U2715 ( .A1(n17728), .A2(n15616), .B1(n17725), .B2(n12328), .ZN(
        n6040) );
  OAI22_X1 U2716 ( .A1(n17764), .A2(n15416), .B1(n17761), .B2(n14501), .ZN(
        n6037) );
  OAI22_X1 U2717 ( .A1(n17752), .A2(n14041), .B1(n17749), .B2(n12036), .ZN(
        n6038) );
  OAI22_X1 U2718 ( .A1(n17680), .A2(n14564), .B1(n17677), .B2(n12011), .ZN(
        n6051) );
  OAI22_X1 U2719 ( .A1(n17716), .A2(n15627), .B1(n17713), .B2(n11863), .ZN(
        n6048) );
  OAI22_X1 U2720 ( .A1(n17704), .A2(n15650), .B1(n17701), .B2(n14659), .ZN(
        n6049) );
  OAI22_X1 U2721 ( .A1(n17728), .A2(n15617), .B1(n17725), .B2(n12329), .ZN(
        n5854) );
  OAI22_X1 U2722 ( .A1(n17764), .A2(n15417), .B1(n17761), .B2(n14502), .ZN(
        n5850) );
  OAI22_X1 U2723 ( .A1(n17752), .A2(n14043), .B1(n17749), .B2(n12037), .ZN(
        n5851) );
  OAI22_X1 U2724 ( .A1(n17680), .A2(n14565), .B1(n17677), .B2(n12012), .ZN(
        n5866) );
  OAI22_X1 U2725 ( .A1(n17716), .A2(n15628), .B1(n17713), .B2(n11864), .ZN(
        n5861) );
  OAI22_X1 U2726 ( .A1(n17704), .A2(n15651), .B1(n17701), .B2(n14660), .ZN(
        n5862) );
  OAI22_X1 U2727 ( .A1(n17728), .A2(n15618), .B1(n17725), .B2(n12330), .ZN(
        n5669) );
  OAI22_X1 U2728 ( .A1(n17764), .A2(n15418), .B1(n17761), .B2(n14503), .ZN(
        n5664) );
  OAI22_X1 U2729 ( .A1(n17752), .A2(n14045), .B1(n17749), .B2(n12038), .ZN(
        n5665) );
  OAI22_X1 U2730 ( .A1(n17680), .A2(n14566), .B1(n17677), .B2(n12013), .ZN(
        n5680) );
  OAI22_X1 U2731 ( .A1(n17716), .A2(n15629), .B1(n17713), .B2(n11865), .ZN(
        n5674) );
  OAI22_X1 U2732 ( .A1(n17704), .A2(n15652), .B1(n17701), .B2(n14661), .ZN(
        n5677) );
  OAI22_X1 U2733 ( .A1(n17728), .A2(n15619), .B1(n17725), .B2(n12331), .ZN(
        n5482) );
  OAI22_X1 U2734 ( .A1(n17764), .A2(n15419), .B1(n17761), .B2(n14504), .ZN(
        n5478) );
  OAI22_X1 U2735 ( .A1(n17752), .A2(n14047), .B1(n17749), .B2(n12039), .ZN(
        n5480) );
  OAI22_X1 U2736 ( .A1(n17680), .A2(n14567), .B1(n17677), .B2(n12014), .ZN(
        n5493) );
  OAI22_X1 U2737 ( .A1(n17716), .A2(n15630), .B1(n17713), .B2(n11866), .ZN(
        n5489) );
  OAI22_X1 U2738 ( .A1(n17704), .A2(n15653), .B1(n17701), .B2(n14662), .ZN(
        n5491) );
  OAI22_X1 U2739 ( .A1(n17727), .A2(n15590), .B1(n17724), .B2(n12314), .ZN(
        n14148) );
  OAI22_X1 U2740 ( .A1(n17763), .A2(n15427), .B1(n17760), .B2(n14477), .ZN(
        n14113) );
  OAI22_X1 U2741 ( .A1(n17751), .A2(n12355), .B1(n17748), .B2(n12047), .ZN(
        n14126) );
  OAI22_X1 U2742 ( .A1(n17679), .A2(n14546), .B1(n17676), .B2(n11950), .ZN(
        n14175) );
  OAI22_X1 U2743 ( .A1(n17715), .A2(n15585), .B1(n17712), .B2(n11845), .ZN(
        n14157) );
  OAI22_X1 U2744 ( .A1(n17703), .A2(n15317), .B1(n17700), .B2(n14634), .ZN(
        n14161) );
  OAI22_X1 U2745 ( .A1(n14960), .A2(n16427), .B1(n14284), .B2(n16424), .ZN(
        n13900) );
  OAI22_X1 U2746 ( .A1(n14961), .A2(n16427), .B1(n14285), .B2(n16424), .ZN(
        n13858) );
  OAI22_X1 U2747 ( .A1(n14962), .A2(n16427), .B1(n14286), .B2(n16424), .ZN(
        n13816) );
  OAI22_X1 U2748 ( .A1(n14980), .A2(n16427), .B1(n14287), .B2(n16424), .ZN(
        n13774) );
  OAI22_X1 U2749 ( .A1(n14963), .A2(n16427), .B1(n14071), .B2(n16424), .ZN(
        n13732) );
  OAI22_X1 U2750 ( .A1(n14964), .A2(n16427), .B1(n14212), .B2(n16424), .ZN(
        n13690) );
  OAI22_X1 U2751 ( .A1(n14868), .A2(n16427), .B1(n14053), .B2(n16424), .ZN(
        n13648) );
  OAI22_X1 U2752 ( .A1(n14965), .A2(n16427), .B1(n14216), .B2(n16424), .ZN(
        n13606) );
  OAI22_X1 U2753 ( .A1(n14966), .A2(n16427), .B1(n14219), .B2(n16424), .ZN(
        n13564) );
  OAI22_X1 U2754 ( .A1(n14967), .A2(n16427), .B1(n14225), .B2(n16424), .ZN(
        n13522) );
  OAI22_X1 U2755 ( .A1(n14968), .A2(n16427), .B1(n14227), .B2(n16424), .ZN(
        n13480) );
  OAI22_X1 U2756 ( .A1(n14969), .A2(n16427), .B1(n14230), .B2(n16424), .ZN(
        n13438) );
  OAI22_X1 U2757 ( .A1(n14970), .A2(n16428), .B1(n14235), .B2(n16425), .ZN(
        n13396) );
  OAI22_X1 U2758 ( .A1(n14971), .A2(n16428), .B1(n14242), .B2(n16425), .ZN(
        n13354) );
  OAI22_X1 U2759 ( .A1(n14972), .A2(n16428), .B1(n14243), .B2(n16425), .ZN(
        n13312) );
  OAI22_X1 U2760 ( .A1(n14973), .A2(n16428), .B1(n14246), .B2(n16425), .ZN(
        n13270) );
  OAI22_X1 U2761 ( .A1(n14974), .A2(n16428), .B1(n14255), .B2(n16425), .ZN(
        n13228) );
  OAI22_X1 U2762 ( .A1(n14975), .A2(n16428), .B1(n14261), .B2(n16425), .ZN(
        n13186) );
  OAI22_X1 U2763 ( .A1(n14976), .A2(n16428), .B1(n14264), .B2(n16425), .ZN(
        n13144) );
  OAI22_X1 U2764 ( .A1(n14977), .A2(n16428), .B1(n14269), .B2(n16425), .ZN(
        n13102) );
  OAI22_X1 U2765 ( .A1(n14978), .A2(n16428), .B1(n14270), .B2(n16425), .ZN(
        n13060) );
  OAI22_X1 U2766 ( .A1(n14981), .A2(n16428), .B1(n14271), .B2(n16425), .ZN(
        n13018) );
  OAI22_X1 U2767 ( .A1(n14982), .A2(n16428), .B1(n14268), .B2(n16425), .ZN(
        n12976) );
  OAI22_X1 U2768 ( .A1(n14979), .A2(n16428), .B1(n14272), .B2(n16425), .ZN(
        n12934) );
  OAI22_X1 U2769 ( .A1(n16680), .A2(n14965), .B1(n14216), .B2(n16677), .ZN(
        n11674) );
  OAI22_X1 U2770 ( .A1(n16680), .A2(n14966), .B1(n14219), .B2(n16677), .ZN(
        n11631) );
  OAI22_X1 U2771 ( .A1(n16680), .A2(n14967), .B1(n14225), .B2(n16677), .ZN(
        n11588) );
  OAI22_X1 U2772 ( .A1(n16680), .A2(n14968), .B1(n14227), .B2(n16677), .ZN(
        n11545) );
  OAI22_X1 U2773 ( .A1(n16680), .A2(n14969), .B1(n14230), .B2(n16677), .ZN(
        n11502) );
  OAI22_X1 U2774 ( .A1(n16680), .A2(n14970), .B1(n14235), .B2(n16677), .ZN(
        n11458) );
  OAI22_X1 U2775 ( .A1(n16680), .A2(n14971), .B1(n14242), .B2(n16677), .ZN(
        n11415) );
  OAI22_X1 U2776 ( .A1(n16680), .A2(n14972), .B1(n14243), .B2(n16677), .ZN(
        n11372) );
  OAI22_X1 U2777 ( .A1(n16680), .A2(n14973), .B1(n14246), .B2(n16677), .ZN(
        n11329) );
  OAI22_X1 U2778 ( .A1(n16680), .A2(n14974), .B1(n14255), .B2(n16677), .ZN(
        n11286) );
  OAI22_X1 U2779 ( .A1(n16680), .A2(n14975), .B1(n14261), .B2(n16677), .ZN(
        n11243) );
  OAI22_X1 U2780 ( .A1(n16680), .A2(n14976), .B1(n14264), .B2(n16676), .ZN(
        n11200) );
  OAI22_X1 U2781 ( .A1(n16679), .A2(n14977), .B1(n14269), .B2(n16676), .ZN(
        n11157) );
  OAI22_X1 U2782 ( .A1(n16679), .A2(n14978), .B1(n14270), .B2(n16676), .ZN(
        n11114) );
  OAI22_X1 U2783 ( .A1(n16679), .A2(n14981), .B1(n14271), .B2(n16676), .ZN(
        n11071) );
  OAI22_X1 U2784 ( .A1(n16679), .A2(n14982), .B1(n14268), .B2(n16676), .ZN(
        n11028) );
  OAI22_X1 U2785 ( .A1(n16679), .A2(n14979), .B1(n14272), .B2(n16677), .ZN(
        n10985) );
  OAI22_X1 U2786 ( .A1(n16679), .A2(n14983), .B1(n14273), .B2(n16676), .ZN(
        n10942) );
  OAI22_X1 U2787 ( .A1(n16679), .A2(n14984), .B1(n14274), .B2(n16676), .ZN(
        n10899) );
  OAI22_X1 U2788 ( .A1(n16679), .A2(n14985), .B1(n14275), .B2(n16676), .ZN(
        n10856) );
  OAI22_X1 U2789 ( .A1(n16679), .A2(n14986), .B1(n14276), .B2(n16676), .ZN(
        n10813) );
  OAI22_X1 U2790 ( .A1(n16679), .A2(n14987), .B1(n14277), .B2(n16676), .ZN(
        n10770) );
  OAI22_X1 U2791 ( .A1(n16679), .A2(n14988), .B1(n14278), .B2(n16676), .ZN(
        n10727) );
  OAI22_X1 U2792 ( .A1(n16679), .A2(n14860), .B1(n14052), .B2(n16676), .ZN(
        n10668) );
  NOR3_X1 U2793 ( .A1(N9908), .A2(n14178), .A3(N9910), .ZN(n14193) );
  INV_X1 U2794 ( .A(n14095), .ZN(n14090) );
  OAI22_X1 U2795 ( .A1(n16372), .A2(n15203), .B1(n16369), .B2(n12199), .ZN(
        n12906) );
  OAI22_X1 U2796 ( .A1(n16372), .A2(n15204), .B1(n16369), .B2(n12200), .ZN(
        n12864) );
  OAI22_X1 U2797 ( .A1(n16372), .A2(n15205), .B1(n16369), .B2(n12201), .ZN(
        n12822) );
  OAI22_X1 U2798 ( .A1(n16372), .A2(n15206), .B1(n16369), .B2(n12202), .ZN(
        n12780) );
  OAI22_X1 U2799 ( .A1(n16372), .A2(n15207), .B1(n16369), .B2(n12203), .ZN(
        n12738) );
  OAI22_X1 U2800 ( .A1(n16372), .A2(n15208), .B1(n16369), .B2(n12204), .ZN(
        n12696) );
  OAI22_X1 U2801 ( .A1(n16372), .A2(n14873), .B1(n16369), .B2(n12161), .ZN(
        n12653) );
  OAI22_X1 U2802 ( .A1(n16372), .A2(n15209), .B1(n16369), .B2(n12307), .ZN(
        n12554) );
  OAI22_X1 U2803 ( .A1(n16624), .A2(n15203), .B1(n16621), .B2(n12199), .ZN(
        n10956) );
  OAI22_X1 U2804 ( .A1(n16624), .A2(n15204), .B1(n16621), .B2(n12200), .ZN(
        n10913) );
  OAI22_X1 U2805 ( .A1(n16624), .A2(n15205), .B1(n16621), .B2(n12201), .ZN(
        n10870) );
  OAI22_X1 U2806 ( .A1(n16624), .A2(n15206), .B1(n16621), .B2(n12202), .ZN(
        n10827) );
  OAI22_X1 U2807 ( .A1(n16624), .A2(n15207), .B1(n16621), .B2(n12203), .ZN(
        n10784) );
  OAI22_X1 U2808 ( .A1(n16624), .A2(n15208), .B1(n16621), .B2(n12204), .ZN(
        n10741) );
  OAI22_X1 U2809 ( .A1(n16624), .A2(n14873), .B1(n16621), .B2(n12161), .ZN(
        n10685) );
  OAI22_X1 U2810 ( .A1(n16624), .A2(n15209), .B1(n16621), .B2(n12307), .ZN(
        n10557) );
  NAND2_X1 U2811 ( .A1(n14007), .A2(n14020), .ZN(n14009) );
  BUF_X1 U2812 ( .A(n4240), .Z(n17635) );
  BUF_X1 U2813 ( .A(n4240), .Z(n17634) );
  BUF_X1 U2814 ( .A(n12527), .Z(n16416) );
  BUF_X1 U2815 ( .A(n12527), .Z(n16415) );
  BUF_X1 U2816 ( .A(n10525), .Z(n16668) );
  BUF_X1 U2817 ( .A(n10525), .Z(n16667) );
  OAI22_X1 U2818 ( .A1(n16370), .A2(n15181), .B1(n16367), .B2(n12205), .ZN(
        n13934) );
  OAI22_X1 U2819 ( .A1(n16370), .A2(n15182), .B1(n16367), .B2(n12206), .ZN(
        n13872) );
  OAI22_X1 U2820 ( .A1(n16370), .A2(n15183), .B1(n16367), .B2(n12207), .ZN(
        n13830) );
  OAI22_X1 U2821 ( .A1(n16370), .A2(n15001), .B1(n16367), .B2(n12208), .ZN(
        n13788) );
  OAI22_X1 U2822 ( .A1(n16370), .A2(n15002), .B1(n16367), .B2(n12195), .ZN(
        n13746) );
  OAI22_X1 U2823 ( .A1(n16370), .A2(n15184), .B1(n16367), .B2(n12209), .ZN(
        n13704) );
  OAI22_X1 U2824 ( .A1(n16370), .A2(n15185), .B1(n16367), .B2(n12210), .ZN(
        n13662) );
  OAI22_X1 U2825 ( .A1(n16370), .A2(n15186), .B1(n16367), .B2(n12211), .ZN(
        n13620) );
  OAI22_X1 U2826 ( .A1(n16370), .A2(n15187), .B1(n16367), .B2(n12212), .ZN(
        n13578) );
  OAI22_X1 U2827 ( .A1(n16370), .A2(n15188), .B1(n16367), .B2(n12213), .ZN(
        n13536) );
  OAI22_X1 U2828 ( .A1(n16370), .A2(n15189), .B1(n16367), .B2(n12214), .ZN(
        n13494) );
  OAI22_X1 U2829 ( .A1(n16370), .A2(n15190), .B1(n16367), .B2(n12215), .ZN(
        n13452) );
  OAI22_X1 U2830 ( .A1(n16371), .A2(n15191), .B1(n16368), .B2(n12253), .ZN(
        n13410) );
  OAI22_X1 U2831 ( .A1(n16371), .A2(n15192), .B1(n16368), .B2(n12254), .ZN(
        n13368) );
  OAI22_X1 U2832 ( .A1(n16371), .A2(n15193), .B1(n16368), .B2(n12255), .ZN(
        n13326) );
  OAI22_X1 U2833 ( .A1(n16371), .A2(n15194), .B1(n16368), .B2(n12256), .ZN(
        n13284) );
  OAI22_X1 U2834 ( .A1(n16371), .A2(n15195), .B1(n16368), .B2(n12257), .ZN(
        n13242) );
  OAI22_X1 U2835 ( .A1(n16371), .A2(n15196), .B1(n16368), .B2(n12258), .ZN(
        n13200) );
  OAI22_X1 U2836 ( .A1(n16371), .A2(n15197), .B1(n16368), .B2(n12301), .ZN(
        n13158) );
  OAI22_X1 U2837 ( .A1(n16371), .A2(n15198), .B1(n16368), .B2(n12303), .ZN(
        n13116) );
  OAI22_X1 U2838 ( .A1(n16371), .A2(n15199), .B1(n16368), .B2(n12304), .ZN(
        n13074) );
  OAI22_X1 U2839 ( .A1(n16371), .A2(n15200), .B1(n16368), .B2(n12305), .ZN(
        n13032) );
  OAI22_X1 U2840 ( .A1(n16371), .A2(n15201), .B1(n16368), .B2(n12306), .ZN(
        n12990) );
  OAI22_X1 U2841 ( .A1(n16371), .A2(n15202), .B1(n16368), .B2(n12198), .ZN(
        n12948) );
  OAI22_X1 U2842 ( .A1(n16622), .A2(n15181), .B1(n16619), .B2(n12205), .ZN(
        n12453) );
  OAI22_X1 U2843 ( .A1(n16622), .A2(n15182), .B1(n16619), .B2(n12206), .ZN(
        n12276) );
  OAI22_X1 U2844 ( .A1(n16622), .A2(n15183), .B1(n16619), .B2(n12207), .ZN(
        n12123) );
  OAI22_X1 U2845 ( .A1(n16622), .A2(n15001), .B1(n16619), .B2(n12208), .ZN(
        n11970) );
  OAI22_X1 U2846 ( .A1(n16622), .A2(n15002), .B1(n16619), .B2(n12195), .ZN(
        n11817) );
  OAI22_X1 U2847 ( .A1(n16622), .A2(n15184), .B1(n16619), .B2(n12209), .ZN(
        n11774) );
  OAI22_X1 U2848 ( .A1(n16622), .A2(n15185), .B1(n16619), .B2(n12210), .ZN(
        n11731) );
  OAI22_X1 U2849 ( .A1(n16622), .A2(n15186), .B1(n16619), .B2(n12211), .ZN(
        n11688) );
  OAI22_X1 U2850 ( .A1(n16622), .A2(n15187), .B1(n16619), .B2(n12212), .ZN(
        n11645) );
  OAI22_X1 U2851 ( .A1(n16622), .A2(n15188), .B1(n16619), .B2(n12213), .ZN(
        n11602) );
  OAI22_X1 U2852 ( .A1(n16622), .A2(n15189), .B1(n16619), .B2(n12214), .ZN(
        n11559) );
  OAI22_X1 U2853 ( .A1(n16622), .A2(n15190), .B1(n16619), .B2(n12215), .ZN(
        n11516) );
  OAI22_X1 U2854 ( .A1(n16623), .A2(n15191), .B1(n16620), .B2(n12253), .ZN(
        n11473) );
  OAI22_X1 U2855 ( .A1(n16623), .A2(n15192), .B1(n16620), .B2(n12254), .ZN(
        n11429) );
  OAI22_X1 U2856 ( .A1(n16623), .A2(n15193), .B1(n16620), .B2(n12255), .ZN(
        n11386) );
  OAI22_X1 U2857 ( .A1(n16623), .A2(n15194), .B1(n16620), .B2(n12256), .ZN(
        n11343) );
  OAI22_X1 U2858 ( .A1(n16623), .A2(n15195), .B1(n16620), .B2(n12257), .ZN(
        n11300) );
  OAI22_X1 U2859 ( .A1(n16623), .A2(n15196), .B1(n16620), .B2(n12258), .ZN(
        n11257) );
  OAI22_X1 U2860 ( .A1(n16623), .A2(n15197), .B1(n16620), .B2(n12301), .ZN(
        n11214) );
  OAI22_X1 U2861 ( .A1(n16623), .A2(n15198), .B1(n16620), .B2(n12303), .ZN(
        n11171) );
  OAI22_X1 U2862 ( .A1(n16623), .A2(n15199), .B1(n16620), .B2(n12304), .ZN(
        n11128) );
  OAI22_X1 U2863 ( .A1(n16623), .A2(n15200), .B1(n16620), .B2(n12305), .ZN(
        n11085) );
  OAI22_X1 U2864 ( .A1(n16623), .A2(n15201), .B1(n16620), .B2(n12306), .ZN(
        n11042) );
  OAI22_X1 U2865 ( .A1(n16623), .A2(n15202), .B1(n16620), .B2(n12198), .ZN(
        n10999) );
  NOR2_X1 U2866 ( .A1(n12492), .A2(n12493), .ZN(n10649) );
  NAND2_X1 U2867 ( .A1(n14158), .A2(n14095), .ZN(n4184) );
  NAND2_X1 U2868 ( .A1(n14094), .A2(n14095), .ZN(n4119) );
  NAND2_X1 U2869 ( .A1(n14104), .A2(n14095), .ZN(n4126) );
  NAND2_X1 U2870 ( .A1(n14107), .A2(n14095), .ZN(n4135) );
  NAND2_X1 U2871 ( .A1(n14108), .A2(n14095), .ZN(n4133) );
  NOR2_X1 U2872 ( .A1(n14100), .A2(n14020), .ZN(n14180) );
  NAND2_X1 U2873 ( .A1(datain[6]), .A2(n18038), .ZN(n7652) );
  NAND2_X1 U2874 ( .A1(n14137), .A2(N9925), .ZN(n14131) );
  NAND2_X1 U2875 ( .A1(n14202), .A2(N9925), .ZN(n14145) );
  NAND2_X1 U2876 ( .A1(n14263), .A2(N273), .ZN(n14066) );
  NOR2_X1 U2877 ( .A1(n14172), .A2(n14020), .ZN(n14204) );
  BUF_X1 U2878 ( .A(n4223), .Z(n17665) );
  BUF_X1 U2879 ( .A(n4223), .Z(n17664) );
  BUF_X1 U2880 ( .A(n4202), .Z(n17689) );
  BUF_X1 U2881 ( .A(n4202), .Z(n17688) );
  BUF_X1 U2882 ( .A(n4240), .Z(n17636) );
  NOR2_X1 U2883 ( .A1(n13976), .A2(N46301), .ZN(n13937) );
  NOR2_X1 U2884 ( .A1(n12495), .A2(N45787), .ZN(n12456) );
  NOR2_X1 U2885 ( .A1(n13975), .A2(N46300), .ZN(n13961) );
  NOR2_X1 U2886 ( .A1(n12494), .A2(N45786), .ZN(n12480) );
  NOR2_X1 U2887 ( .A1(N46301), .A2(N46300), .ZN(n13958) );
  NOR2_X1 U2888 ( .A1(N45787), .A2(N45786), .ZN(n12475) );
  NOR2_X1 U2889 ( .A1(n14144), .A2(n14820), .ZN(n14179) );
  OAI22_X1 U2890 ( .A1(n16700), .A2(n14960), .B1(n16439), .B2(n16692), .ZN(
        n7759) );
  OAI22_X1 U2891 ( .A1(n17585), .A2(n14284), .B1(n16439), .B2(n17577), .ZN(
        n7798) );
  OAI22_X1 U2892 ( .A1(n17836), .A2(n14506), .B1(n16439), .B2(n17839), .ZN(
        n7800) );
  OAI22_X1 U2893 ( .A1(n17880), .A2(n15574), .B1(n16439), .B2(n17883), .ZN(
        n7801) );
  OAI22_X1 U2894 ( .A1(n17923), .A2(n15432), .B1(n16439), .B2(n17926), .ZN(
        n7802) );
  OAI22_X1 U2895 ( .A1(n17965), .A2(n15245), .B1(n16439), .B2(n17968), .ZN(
        n7803) );
  OAI22_X1 U2896 ( .A1(n18012), .A2(n12055), .B1(n16439), .B2(n18003), .ZN(
        n7804) );
  OAI22_X1 U2897 ( .A1(n16887), .A2(n15369), .B1(n16439), .B2(n16888), .ZN(
        n7806) );
  OAI22_X1 U2898 ( .A1(n16910), .A2(n14484), .B1(n16439), .B2(n16911), .ZN(
        n7807) );
  OAI22_X1 U2899 ( .A1(n16943), .A2(n14547), .B1(n16440), .B2(n16934), .ZN(
        n7808) );
  OAI22_X1 U2900 ( .A1(n16956), .A2(n14772), .B1(n16440), .B2(n16957), .ZN(
        n7809) );
  OAI22_X1 U2901 ( .A1(n16976), .A2(n14888), .B1(n16440), .B2(n16977), .ZN(
        n7810) );
  OAI22_X1 U2902 ( .A1(n16999), .A2(n14427), .B1(n16440), .B2(n17000), .ZN(
        n7811) );
  OAI22_X1 U2903 ( .A1(n17032), .A2(n12171), .B1(n16440), .B2(n17023), .ZN(
        n7812) );
  OAI22_X1 U2904 ( .A1(n17058), .A2(n14359), .B1(n16440), .B2(n17049), .ZN(
        n7813) );
  OAI22_X1 U2905 ( .A1(n17084), .A2(n15575), .B1(n16440), .B2(n17075), .ZN(
        n7814) );
  OAI22_X1 U2906 ( .A1(n17110), .A2(n11713), .B1(n16440), .B2(n17101), .ZN(
        n7815) );
  OAI22_X1 U2907 ( .A1(n17136), .A2(n15736), .B1(n16440), .B2(n17127), .ZN(
        n7816) );
  OAI22_X1 U2908 ( .A1(n17171), .A2(n12018), .B1(n16440), .B2(n17172), .ZN(
        n7818) );
  OAI22_X1 U2909 ( .A1(n17192), .A2(n14300), .B1(n16440), .B2(n17193), .ZN(
        n7819) );
  OAI22_X1 U2910 ( .A1(n17251), .A2(n12205), .B1(n16441), .B2(n17242), .ZN(
        n7821) );
  OAI22_X1 U2911 ( .A1(n17303), .A2(n14605), .B1(n16441), .B2(n17294), .ZN(
        n7823) );
  OAI22_X1 U2912 ( .A1(n17329), .A2(n15292), .B1(n16441), .B2(n17320), .ZN(
        n7824) );
  OAI22_X1 U2913 ( .A1(n17355), .A2(n15072), .B1(n16441), .B2(n17346), .ZN(
        n7825) );
  OAI22_X1 U2914 ( .A1(n17381), .A2(n14426), .B1(n16441), .B2(n17372), .ZN(
        n7826) );
  OAI22_X1 U2915 ( .A1(n17407), .A2(n14329), .B1(n16441), .B2(n17398), .ZN(
        n7827) );
  OAI22_X1 U2916 ( .A1(n17433), .A2(n15326), .B1(n16441), .B2(n17424), .ZN(
        n7828) );
  OAI22_X1 U2917 ( .A1(n17459), .A2(n14711), .B1(n16441), .B2(n17451), .ZN(
        n7829) );
  OAI22_X1 U2918 ( .A1(n17485), .A2(n15758), .B1(n16441), .B2(n17476), .ZN(
        n7830) );
  OAI22_X1 U2919 ( .A1(n17511), .A2(n15576), .B1(n16441), .B2(n17502), .ZN(
        n7831) );
  OAI22_X1 U2920 ( .A1(n16700), .A2(n14961), .B1(n16445), .B2(n16692), .ZN(
        n7833) );
  OAI22_X1 U2921 ( .A1(n17585), .A2(n14285), .B1(n16445), .B2(n17577), .ZN(
        n7872) );
  OAI22_X1 U2922 ( .A1(n17838), .A2(n14507), .B1(n16445), .B2(n17839), .ZN(
        n7874) );
  OAI22_X1 U2923 ( .A1(n17860), .A2(n15124), .B1(n16445), .B2(n17861), .ZN(
        n7875) );
  OAI22_X1 U2924 ( .A1(n17925), .A2(n15433), .B1(n16445), .B2(n17926), .ZN(
        n7876) );
  OAI22_X1 U2925 ( .A1(n17946), .A2(n14911), .B1(n16445), .B2(n17947), .ZN(
        n7877) );
  OAI22_X1 U2926 ( .A1(n18012), .A2(n12052), .B1(n16445), .B2(n18003), .ZN(
        n7878) );
  OAI22_X1 U2927 ( .A1(n18025), .A2(n14570), .B1(n16445), .B2(n18016), .ZN(
        n7879) );
  OAI22_X1 U2928 ( .A1(n16887), .A2(n15370), .B1(n16445), .B2(n16888), .ZN(
        n7880) );
  OAI22_X1 U2929 ( .A1(n16943), .A2(n14548), .B1(n16446), .B2(n16934), .ZN(
        n7882) );
  OAI22_X1 U2930 ( .A1(n16945), .A2(n11952), .B1(n16446), .B2(n16946), .ZN(
        n7883) );
  OAI22_X1 U2931 ( .A1(n16976), .A2(n14889), .B1(n16446), .B2(n16977), .ZN(
        n7884) );
  OAI22_X1 U2932 ( .A1(n17032), .A2(n12172), .B1(n16446), .B2(n17023), .ZN(
        n7886) );
  OAI22_X1 U2933 ( .A1(n17045), .A2(n15035), .B1(n16446), .B2(n17036), .ZN(
        n7887) );
  OAI22_X1 U2934 ( .A1(n17084), .A2(n15577), .B1(n16446), .B2(n17075), .ZN(
        n7888) );
  OAI22_X1 U2935 ( .A1(n17097), .A2(n15496), .B1(n16446), .B2(n17088), .ZN(
        n7889) );
  OAI22_X1 U2936 ( .A1(n17136), .A2(n15737), .B1(n16446), .B2(n17127), .ZN(
        n7890) );
  OAI22_X1 U2937 ( .A1(n17137), .A2(n14679), .B1(n16446), .B2(n17138), .ZN(
        n7891) );
  OAI22_X1 U2938 ( .A1(n17171), .A2(n12019), .B1(n16446), .B2(n17172), .ZN(
        n7892) );
  OAI22_X1 U2939 ( .A1(n17182), .A2(n12358), .B1(n16446), .B2(n17183), .ZN(
        n7893) );
  OAI22_X1 U2940 ( .A1(n17238), .A2(n15371), .B1(n16447), .B2(n17229), .ZN(
        n7895) );
  OAI22_X1 U2941 ( .A1(n17290), .A2(n14360), .B1(n16447), .B2(n17281), .ZN(
        n7897) );
  OAI22_X1 U2942 ( .A1(n17329), .A2(n15293), .B1(n16447), .B2(n17320), .ZN(
        n7898) );
  OAI22_X1 U2943 ( .A1(n17342), .A2(n11882), .B1(n16447), .B2(n17333), .ZN(
        n7899) );
  OAI22_X1 U2944 ( .A1(n17381), .A2(n14428), .B1(n16447), .B2(n17372), .ZN(
        n7900) );
  OAI22_X1 U2945 ( .A1(n17394), .A2(n14714), .B1(n16447), .B2(n17385), .ZN(
        n7901) );
  OAI22_X1 U2946 ( .A1(n17433), .A2(n15327), .B1(n16447), .B2(n17424), .ZN(
        n7902) );
  OAI22_X1 U2947 ( .A1(n17446), .A2(n12359), .B1(n16447), .B2(n17437), .ZN(
        n7903) );
  OAI22_X1 U2948 ( .A1(n17485), .A2(n15759), .B1(n16447), .B2(n17476), .ZN(
        n7904) );
  OAI22_X1 U2949 ( .A1(n17498), .A2(n14773), .B1(n16447), .B2(n17489), .ZN(
        n7905) );
  OAI22_X1 U2950 ( .A1(n16700), .A2(n14962), .B1(n16451), .B2(n16692), .ZN(
        n7907) );
  OAI22_X1 U2951 ( .A1(n17838), .A2(n14508), .B1(n16451), .B2(n17840), .ZN(
        n7948) );
  OAI22_X1 U2952 ( .A1(n17860), .A2(n15125), .B1(n16451), .B2(n17861), .ZN(
        n7949) );
  OAI22_X1 U2953 ( .A1(n17882), .A2(n15578), .B1(n16451), .B2(n17883), .ZN(
        n7950) );
  OAI22_X1 U2954 ( .A1(n17904), .A2(n14643), .B1(n16451), .B2(n17905), .ZN(
        n7951) );
  OAI22_X1 U2955 ( .A1(n18012), .A2(n12053), .B1(n16451), .B2(n18003), .ZN(
        n7952) );
  OAI22_X1 U2956 ( .A1(n18025), .A2(n14571), .B1(n16451), .B2(n18016), .ZN(
        n7953) );
  OAI22_X1 U2957 ( .A1(n16877), .A2(n14940), .B1(n16451), .B2(n16878), .ZN(
        n7955) );
  OAI22_X1 U2958 ( .A1(n16943), .A2(n14549), .B1(n16452), .B2(n16934), .ZN(
        n7956) );
  OAI22_X1 U2959 ( .A1(n16945), .A2(n11995), .B1(n16452), .B2(n16946), .ZN(
        n7957) );
  OAI22_X1 U2960 ( .A1(n16956), .A2(n14776), .B1(n16452), .B2(n16957), .ZN(
        n7958) );
  OAI22_X1 U2961 ( .A1(n16966), .A2(n15468), .B1(n16452), .B2(n16967), .ZN(
        n7959) );
  OAI22_X1 U2962 ( .A1(n17032), .A2(n12173), .B1(n16452), .B2(n17023), .ZN(
        n7960) );
  OAI22_X1 U2963 ( .A1(n17045), .A2(n15036), .B1(n16452), .B2(n17036), .ZN(
        n7961) );
  OAI22_X1 U2964 ( .A1(n17058), .A2(n14361), .B1(n16452), .B2(n17049), .ZN(
        n7962) );
  OAI22_X1 U2965 ( .A1(n17071), .A2(n15151), .B1(n16452), .B2(n17062), .ZN(
        n7963) );
  OAI22_X1 U2966 ( .A1(n17136), .A2(n15738), .B1(n16452), .B2(n17127), .ZN(
        n7964) );
  OAI22_X1 U2967 ( .A1(n17137), .A2(n14680), .B1(n16452), .B2(n17138), .ZN(
        n7965) );
  OAI22_X1 U2968 ( .A1(n17160), .A2(n15006), .B1(n16452), .B2(n17161), .ZN(
        n7967) );
  OAI22_X1 U2969 ( .A1(n17238), .A2(n15372), .B1(n16453), .B2(n17229), .ZN(
        n7969) );
  OAI22_X1 U2970 ( .A1(n17251), .A2(n12207), .B1(n16453), .B2(n17242), .ZN(
        n7970) );
  OAI22_X1 U2971 ( .A1(n17264), .A2(n14833), .B1(n16453), .B2(n17255), .ZN(
        n7971) );
  OAI22_X1 U2972 ( .A1(n17329), .A2(n15294), .B1(n16453), .B2(n17320), .ZN(
        n7972) );
  OAI22_X1 U2973 ( .A1(n17342), .A2(n11883), .B1(n16453), .B2(n17333), .ZN(
        n7973) );
  OAI22_X1 U2974 ( .A1(n17355), .A2(n15076), .B1(n16453), .B2(n17346), .ZN(
        n7974) );
  OAI22_X1 U2975 ( .A1(n17368), .A2(n15671), .B1(n16453), .B2(n17359), .ZN(
        n7975) );
  OAI22_X1 U2976 ( .A1(n17433), .A2(n15328), .B1(n16453), .B2(n17424), .ZN(
        n7976) );
  OAI22_X1 U2977 ( .A1(n17446), .A2(n12361), .B1(n16453), .B2(n17437), .ZN(
        n7977) );
  OAI22_X1 U2978 ( .A1(n17459), .A2(n14715), .B1(n16453), .B2(n17451), .ZN(
        n7978) );
  OAI22_X1 U2979 ( .A1(n17472), .A2(n15523), .B1(n16453), .B2(n17463), .ZN(
        n7979) );
  OAI22_X1 U2980 ( .A1(n17123), .A2(n12309), .B1(n17115), .B2(n16437), .ZN(
        n7780) );
  OAI22_X1 U2981 ( .A1(n17316), .A2(n15699), .B1(n17308), .B2(n16438), .ZN(
        n7788) );
  OAI22_X1 U2982 ( .A1(n17420), .A2(n15210), .B1(n17412), .B2(n16438), .ZN(
        n7792) );
  OAI22_X1 U2983 ( .A1(n17123), .A2(n12310), .B1(n17114), .B2(n16443), .ZN(
        n7855) );
  OAI22_X1 U2984 ( .A1(n17316), .A2(n15700), .B1(n17307), .B2(n16444), .ZN(
        n7863) );
  OAI22_X1 U2985 ( .A1(n17420), .A2(n15211), .B1(n17411), .B2(n16444), .ZN(
        n7867) );
  OAI22_X1 U2986 ( .A1(n17123), .A2(n12311), .B1(n17114), .B2(n16449), .ZN(
        n7931) );
  OAI22_X1 U2987 ( .A1(n17316), .A2(n15701), .B1(n17307), .B2(n16450), .ZN(
        n7939) );
  OAI22_X1 U2988 ( .A1(n17420), .A2(n15212), .B1(n17411), .B2(n16450), .ZN(
        n7943) );
  OAI22_X1 U2989 ( .A1(n17122), .A2(n12312), .B1(n17114), .B2(n16457), .ZN(
        n8005) );
  OAI22_X1 U2990 ( .A1(n17315), .A2(n15702), .B1(n17307), .B2(n16458), .ZN(
        n8013) );
  OAI22_X1 U2991 ( .A1(n17122), .A2(n12313), .B1(n17115), .B2(n16710), .ZN(
        n8133) );
  OAI22_X1 U2992 ( .A1(n17419), .A2(n15213), .B1(n17411), .B2(n16711), .ZN(
        n8149) );
  OAI22_X1 U2993 ( .A1(n17315), .A2(n15703), .B1(n17308), .B2(n16719), .ZN(
        n8213) );
  OAI22_X1 U2994 ( .A1(n17419), .A2(n15214), .B1(n17412), .B2(n16720), .ZN(
        n8221) );
  OAI22_X1 U2995 ( .A1(n17123), .A2(n12314), .B1(n17115), .B2(n16705), .ZN(
        n10093) );
  OAI22_X1 U2996 ( .A1(n17316), .A2(n15721), .B1(n17308), .B2(n16703), .ZN(
        n10109) );
  OAI22_X1 U2997 ( .A1(n17420), .A2(n15239), .B1(n17412), .B2(n16703), .ZN(
        n10117) );
  NOR2_X1 U2998 ( .A1(n13981), .A2(n13982), .ZN(n13962) );
  INV_X1 U2999 ( .A(n13983), .ZN(n13982) );
  NOR2_X1 U3000 ( .A1(n12500), .A2(n12501), .ZN(n12481) );
  INV_X1 U3001 ( .A(n12502), .ZN(n12501) );
  OAI22_X1 U3002 ( .A1(n17484), .A2(n15764), .B1(n17476), .B2(n16730), .ZN(
        n8322) );
  OAI22_X1 U3003 ( .A1(n17497), .A2(n14781), .B1(n17490), .B2(n16730), .ZN(
        n8323) );
  OAI22_X1 U3004 ( .A1(n17510), .A2(n15579), .B1(n17503), .B2(n16730), .ZN(
        n8324) );
  OAI22_X1 U3005 ( .A1(n17446), .A2(n12357), .B1(n17438), .B2(n16438), .ZN(
        n7793) );
  OAI22_X1 U3006 ( .A1(n17472), .A2(n15521), .B1(n17464), .B2(n16438), .ZN(
        n7794) );
  OAI22_X1 U3007 ( .A1(n17498), .A2(n14771), .B1(n17490), .B2(n16438), .ZN(
        n7795) );
  OAI22_X1 U3008 ( .A1(n17459), .A2(n14713), .B1(n17451), .B2(n16444), .ZN(
        n7868) );
  OAI22_X1 U3009 ( .A1(n17472), .A2(n15522), .B1(n17463), .B2(n16444), .ZN(
        n7869) );
  OAI22_X1 U3010 ( .A1(n17511), .A2(n15580), .B1(n17503), .B2(n16444), .ZN(
        n7870) );
  OAI22_X1 U3011 ( .A1(n17485), .A2(n15760), .B1(n17476), .B2(n16450), .ZN(
        n7944) );
  OAI22_X1 U3012 ( .A1(n17498), .A2(n14775), .B1(n17489), .B2(n16450), .ZN(
        n7945) );
  OAI22_X1 U3013 ( .A1(n17511), .A2(n15581), .B1(n17502), .B2(n16450), .ZN(
        n7946) );
  OAI22_X1 U3014 ( .A1(n17432), .A2(n15329), .B1(n17425), .B2(n16458), .ZN(
        n8022) );
  OAI22_X1 U3015 ( .A1(n17445), .A2(n12362), .B1(n17437), .B2(n16458), .ZN(
        n8023) );
  OAI22_X1 U3016 ( .A1(n17458), .A2(n14717), .B1(n17451), .B2(n16458), .ZN(
        n8024) );
  OAI22_X1 U3017 ( .A1(n17471), .A2(n15524), .B1(n17464), .B2(n16458), .ZN(
        n8025) );
  OAI22_X1 U3018 ( .A1(n17484), .A2(n15761), .B1(n17476), .B2(n16459), .ZN(
        n8026) );
  OAI22_X1 U3019 ( .A1(n17497), .A2(n14777), .B1(n17489), .B2(n16459), .ZN(
        n8027) );
  OAI22_X1 U3020 ( .A1(n17510), .A2(n15582), .B1(n17502), .B2(n16459), .ZN(
        n8028) );
  OAI22_X1 U3021 ( .A1(n17432), .A2(n15330), .B1(n17425), .B2(n16711), .ZN(
        n8150) );
  OAI22_X1 U3022 ( .A1(n17445), .A2(n12363), .B1(n17438), .B2(n16711), .ZN(
        n8151) );
  OAI22_X1 U3023 ( .A1(n17458), .A2(n14718), .B1(n17451), .B2(n16711), .ZN(
        n8152) );
  OAI22_X1 U3024 ( .A1(n17471), .A2(n15525), .B1(n17463), .B2(n16711), .ZN(
        n8153) );
  OAI22_X1 U3025 ( .A1(n17484), .A2(n15762), .B1(n17477), .B2(n16712), .ZN(
        n8154) );
  OAI22_X1 U3026 ( .A1(n17497), .A2(n14778), .B1(n17490), .B2(n16712), .ZN(
        n8155) );
  OAI22_X1 U3027 ( .A1(n17510), .A2(n15583), .B1(n17503), .B2(n16712), .ZN(
        n8156) );
  OAI22_X1 U3028 ( .A1(n17432), .A2(n15331), .B1(n17424), .B2(n16720), .ZN(
        n8222) );
  OAI22_X1 U3029 ( .A1(n17445), .A2(n12365), .B1(n17437), .B2(n16720), .ZN(
        n8223) );
  OAI22_X1 U3030 ( .A1(n17458), .A2(n14720), .B1(n17451), .B2(n16720), .ZN(
        n8224) );
  OAI22_X1 U3031 ( .A1(n17471), .A2(n15526), .B1(n17463), .B2(n16720), .ZN(
        n8225) );
  OAI22_X1 U3032 ( .A1(n17484), .A2(n15763), .B1(n17477), .B2(n16721), .ZN(
        n8226) );
  OAI22_X1 U3033 ( .A1(n17497), .A2(n14780), .B1(n17490), .B2(n16721), .ZN(
        n8227) );
  OAI22_X1 U3034 ( .A1(n17510), .A2(n15584), .B1(n17503), .B2(n16721), .ZN(
        n8228) );
  OAI22_X1 U3035 ( .A1(n17432), .A2(n15332), .B1(n17424), .B2(n16729), .ZN(
        n8318) );
  OAI22_X1 U3036 ( .A1(n17445), .A2(n12367), .B1(n17437), .B2(n16729), .ZN(
        n8319) );
  OAI22_X1 U3037 ( .A1(n17458), .A2(n14722), .B1(n17451), .B2(n16729), .ZN(
        n8320) );
  OAI22_X1 U3038 ( .A1(n17431), .A2(n15333), .B1(n17424), .B2(n16736), .ZN(
        n8390) );
  OAI22_X1 U3039 ( .A1(n17433), .A2(n15349), .B1(n17425), .B2(n16703), .ZN(
        n10118) );
  OAI22_X1 U3040 ( .A1(n17446), .A2(n12348), .B1(n17438), .B2(n16702), .ZN(
        n10119) );
  OAI22_X1 U3041 ( .A1(n17459), .A2(n15318), .B1(n17451), .B2(n16703), .ZN(
        n10120) );
  OAI22_X1 U3042 ( .A1(n17472), .A2(n15458), .B1(n17464), .B2(n16702), .ZN(
        n10121) );
  OAI22_X1 U3043 ( .A1(n17485), .A2(n15781), .B1(n17477), .B2(n16702), .ZN(
        n10122) );
  OAI22_X1 U3044 ( .A1(n17498), .A2(n14815), .B1(n17489), .B2(n16702), .ZN(
        n10123) );
  OAI22_X1 U3045 ( .A1(n17511), .A2(n15585), .B1(n17502), .B2(n16702), .ZN(
        n10124) );
  OAI22_X1 U3046 ( .A1(n17045), .A2(n15037), .B1(n17036), .B2(n16437), .ZN(
        n7777) );
  OAI22_X1 U3047 ( .A1(n17071), .A2(n15152), .B1(n17062), .B2(n16437), .ZN(
        n7778) );
  OAI22_X1 U3048 ( .A1(n17097), .A2(n15495), .B1(n17088), .B2(n16437), .ZN(
        n7779) );
  OAI22_X1 U3049 ( .A1(n17238), .A2(n15373), .B1(n17229), .B2(n16438), .ZN(
        n7785) );
  OAI22_X1 U3050 ( .A1(n17264), .A2(n14831), .B1(n17255), .B2(n16438), .ZN(
        n7786) );
  OAI22_X1 U3051 ( .A1(n17290), .A2(n14362), .B1(n17281), .B2(n16438), .ZN(
        n7787) );
  OAI22_X1 U3052 ( .A1(n17342), .A2(n11881), .B1(n17333), .B2(n16438), .ZN(
        n7789) );
  OAI22_X1 U3053 ( .A1(n17368), .A2(n15669), .B1(n17359), .B2(n16438), .ZN(
        n7790) );
  OAI22_X1 U3054 ( .A1(n17394), .A2(n14712), .B1(n17385), .B2(n16438), .ZN(
        n7791) );
  OAI22_X1 U3055 ( .A1(n17058), .A2(n14363), .B1(n17049), .B2(n16443), .ZN(
        n7852) );
  OAI22_X1 U3056 ( .A1(n17071), .A2(n15153), .B1(n17063), .B2(n16443), .ZN(
        n7853) );
  OAI22_X1 U3057 ( .A1(n17110), .A2(n11756), .B1(n17101), .B2(n16443), .ZN(
        n7854) );
  OAI22_X1 U3058 ( .A1(n17251), .A2(n12206), .B1(n17242), .B2(n16444), .ZN(
        n7860) );
  OAI22_X1 U3059 ( .A1(n17264), .A2(n14832), .B1(n17256), .B2(n16444), .ZN(
        n7861) );
  OAI22_X1 U3060 ( .A1(n17303), .A2(n14606), .B1(n17294), .B2(n16444), .ZN(
        n7862) );
  OAI22_X1 U3061 ( .A1(n17355), .A2(n15074), .B1(n17346), .B2(n16444), .ZN(
        n7864) );
  OAI22_X1 U3062 ( .A1(n17368), .A2(n15670), .B1(n17360), .B2(n16444), .ZN(
        n7865) );
  OAI22_X1 U3063 ( .A1(n17407), .A2(n14330), .B1(n17398), .B2(n16444), .ZN(
        n7866) );
  OAI22_X1 U3064 ( .A1(n17084), .A2(n15586), .B1(n17075), .B2(n16449), .ZN(
        n7928) );
  OAI22_X1 U3065 ( .A1(n17097), .A2(n15497), .B1(n17089), .B2(n16449), .ZN(
        n7929) );
  OAI22_X1 U3066 ( .A1(n17110), .A2(n11799), .B1(n17102), .B2(n16449), .ZN(
        n7930) );
  OAI22_X1 U3067 ( .A1(n17290), .A2(n14364), .B1(n17282), .B2(n16450), .ZN(
        n7937) );
  OAI22_X1 U3068 ( .A1(n17303), .A2(n14607), .B1(n17295), .B2(n16450), .ZN(
        n7938) );
  OAI22_X1 U3069 ( .A1(n17381), .A2(n14430), .B1(n17372), .B2(n16450), .ZN(
        n7940) );
  OAI22_X1 U3070 ( .A1(n17394), .A2(n14716), .B1(n17386), .B2(n16450), .ZN(
        n7941) );
  OAI22_X1 U3071 ( .A1(n17407), .A2(n14331), .B1(n17399), .B2(n16450), .ZN(
        n7942) );
  OAI22_X1 U3072 ( .A1(n17031), .A2(n12174), .B1(n17024), .B2(n16457), .ZN(
        n7998) );
  OAI22_X1 U3073 ( .A1(n17044), .A2(n15038), .B1(n17037), .B2(n16457), .ZN(
        n7999) );
  OAI22_X1 U3074 ( .A1(n17057), .A2(n14365), .B1(n17050), .B2(n16457), .ZN(
        n8000) );
  OAI22_X1 U3075 ( .A1(n17070), .A2(n15154), .B1(n17062), .B2(n16457), .ZN(
        n8001) );
  OAI22_X1 U3076 ( .A1(n17083), .A2(n15587), .B1(n17076), .B2(n16457), .ZN(
        n8002) );
  OAI22_X1 U3077 ( .A1(n17096), .A2(n15498), .B1(n17088), .B2(n16457), .ZN(
        n8003) );
  OAI22_X1 U3078 ( .A1(n17109), .A2(n11842), .B1(n17101), .B2(n16457), .ZN(
        n8004) );
  OAI22_X1 U3079 ( .A1(n17237), .A2(n15374), .B1(n17230), .B2(n16458), .ZN(
        n8007) );
  OAI22_X1 U3080 ( .A1(n17250), .A2(n12208), .B1(n17243), .B2(n16458), .ZN(
        n8008) );
  OAI22_X1 U3081 ( .A1(n17263), .A2(n14834), .B1(n17255), .B2(n16458), .ZN(
        n8009) );
  OAI22_X1 U3082 ( .A1(n17289), .A2(n14366), .B1(n17281), .B2(n16458), .ZN(
        n8011) );
  OAI22_X1 U3083 ( .A1(n17302), .A2(n14608), .B1(n17294), .B2(n16458), .ZN(
        n8012) );
  OAI22_X1 U3084 ( .A1(n17031), .A2(n12175), .B1(n17023), .B2(n16710), .ZN(
        n8126) );
  OAI22_X1 U3085 ( .A1(n17044), .A2(n15039), .B1(n17036), .B2(n16710), .ZN(
        n8127) );
  OAI22_X1 U3086 ( .A1(n17057), .A2(n14367), .B1(n17049), .B2(n16710), .ZN(
        n8128) );
  OAI22_X1 U3087 ( .A1(n17070), .A2(n15155), .B1(n17063), .B2(n16710), .ZN(
        n8129) );
  OAI22_X1 U3088 ( .A1(n17083), .A2(n15588), .B1(n17075), .B2(n16710), .ZN(
        n8130) );
  OAI22_X1 U3089 ( .A1(n17096), .A2(n15499), .B1(n17089), .B2(n16710), .ZN(
        n8131) );
  OAI22_X1 U3090 ( .A1(n17109), .A2(n11844), .B1(n17102), .B2(n16710), .ZN(
        n8132) );
  OAI22_X1 U3091 ( .A1(n17328), .A2(n15295), .B1(n17321), .B2(n16711), .ZN(
        n8142) );
  OAI22_X1 U3092 ( .A1(n17341), .A2(n11884), .B1(n17334), .B2(n16711), .ZN(
        n8143) );
  OAI22_X1 U3093 ( .A1(n17354), .A2(n15078), .B1(n17347), .B2(n16711), .ZN(
        n8144) );
  OAI22_X1 U3094 ( .A1(n17367), .A2(n15672), .B1(n17359), .B2(n16711), .ZN(
        n8145) );
  OAI22_X1 U3095 ( .A1(n17380), .A2(n14432), .B1(n17373), .B2(n16711), .ZN(
        n8146) );
  OAI22_X1 U3096 ( .A1(n17393), .A2(n14719), .B1(n17385), .B2(n16711), .ZN(
        n8147) );
  OAI22_X1 U3097 ( .A1(n17406), .A2(n14332), .B1(n17398), .B2(n16711), .ZN(
        n8148) );
  OAI22_X1 U3098 ( .A1(n17237), .A2(n15375), .B1(n17229), .B2(n16719), .ZN(
        n8207) );
  OAI22_X1 U3099 ( .A1(n17250), .A2(n12209), .B1(n17242), .B2(n16719), .ZN(
        n8208) );
  OAI22_X1 U3100 ( .A1(n17263), .A2(n14835), .B1(n17256), .B2(n16719), .ZN(
        n8209) );
  OAI22_X1 U3101 ( .A1(n17289), .A2(n14368), .B1(n17282), .B2(n16719), .ZN(
        n8211) );
  OAI22_X1 U3102 ( .A1(n17302), .A2(n14609), .B1(n17295), .B2(n16719), .ZN(
        n8212) );
  OAI22_X1 U3103 ( .A1(n17328), .A2(n15296), .B1(n17320), .B2(n16720), .ZN(
        n8214) );
  OAI22_X1 U3104 ( .A1(n17341), .A2(n11885), .B1(n17333), .B2(n16720), .ZN(
        n8215) );
  OAI22_X1 U3105 ( .A1(n17354), .A2(n15080), .B1(n17346), .B2(n16720), .ZN(
        n8216) );
  OAI22_X1 U3106 ( .A1(n17367), .A2(n15673), .B1(n17360), .B2(n16720), .ZN(
        n8217) );
  OAI22_X1 U3107 ( .A1(n17380), .A2(n14434), .B1(n17372), .B2(n16720), .ZN(
        n8218) );
  OAI22_X1 U3108 ( .A1(n17393), .A2(n14721), .B1(n17386), .B2(n16720), .ZN(
        n8219) );
  OAI22_X1 U3109 ( .A1(n17406), .A2(n14333), .B1(n17399), .B2(n16720), .ZN(
        n8220) );
  OAI22_X1 U3110 ( .A1(n17031), .A2(n12176), .B1(n17023), .B2(n16727), .ZN(
        n8286) );
  OAI22_X1 U3111 ( .A1(n17044), .A2(n15040), .B1(n17036), .B2(n16727), .ZN(
        n8287) );
  OAI22_X1 U3112 ( .A1(n17057), .A2(n14369), .B1(n17049), .B2(n16727), .ZN(
        n8288) );
  OAI22_X1 U3113 ( .A1(n17083), .A2(n15589), .B1(n17075), .B2(n16727), .ZN(
        n8290) );
  OAI22_X1 U3114 ( .A1(n17237), .A2(n15376), .B1(n17229), .B2(n16728), .ZN(
        n8303) );
  OAI22_X1 U3115 ( .A1(n17250), .A2(n12210), .B1(n17242), .B2(n16728), .ZN(
        n8304) );
  OAI22_X1 U3116 ( .A1(n17328), .A2(n15297), .B1(n17320), .B2(n16729), .ZN(
        n8310) );
  OAI22_X1 U3117 ( .A1(n17341), .A2(n11886), .B1(n17333), .B2(n16729), .ZN(
        n8311) );
  OAI22_X1 U3118 ( .A1(n17354), .A2(n15081), .B1(n17346), .B2(n16729), .ZN(
        n8312) );
  OAI22_X1 U3119 ( .A1(n17380), .A2(n14435), .B1(n17372), .B2(n16729), .ZN(
        n8314) );
  OAI22_X1 U3120 ( .A1(n17031), .A2(n12177), .B1(n17023), .B2(n16733), .ZN(
        n8358) );
  OAI22_X1 U3121 ( .A1(n17328), .A2(n15298), .B1(n17320), .B2(n16735), .ZN(
        n8382) );
  OAI22_X1 U3122 ( .A1(n17032), .A2(n12194), .B1(n17024), .B2(n16705), .ZN(
        n10086) );
  OAI22_X1 U3123 ( .A1(n17045), .A2(n15041), .B1(n17037), .B2(n16705), .ZN(
        n10087) );
  OAI22_X1 U3124 ( .A1(n17058), .A2(n14370), .B1(n17050), .B2(n16705), .ZN(
        n10088) );
  OAI22_X1 U3125 ( .A1(n17071), .A2(n15156), .B1(n17062), .B2(n16705), .ZN(
        n10089) );
  OAI22_X1 U3126 ( .A1(n17084), .A2(n15590), .B1(n17076), .B2(n16705), .ZN(
        n10090) );
  OAI22_X1 U3127 ( .A1(n17097), .A2(n15517), .B1(n17088), .B2(n16705), .ZN(
        n10091) );
  OAI22_X1 U3128 ( .A1(n17110), .A2(n11845), .B1(n17101), .B2(n16705), .ZN(
        n10092) );
  OAI22_X1 U3129 ( .A1(n17238), .A2(n15377), .B1(n17230), .B2(n16704), .ZN(
        n10103) );
  OAI22_X1 U3130 ( .A1(n17251), .A2(n12307), .B1(n17243), .B2(n16704), .ZN(
        n10104) );
  OAI22_X1 U3131 ( .A1(n17264), .A2(n14853), .B1(n17255), .B2(n16704), .ZN(
        n10105) );
  OAI22_X1 U3132 ( .A1(n17290), .A2(n14371), .B1(n17281), .B2(n16703), .ZN(
        n10107) );
  OAI22_X1 U3133 ( .A1(n17303), .A2(n14627), .B1(n17294), .B2(n16704), .ZN(
        n10108) );
  OAI22_X1 U3134 ( .A1(n17329), .A2(n15314), .B1(n17321), .B2(n16703), .ZN(
        n10110) );
  OAI22_X1 U3135 ( .A1(n17342), .A2(n11903), .B1(n17334), .B2(n16703), .ZN(
        n10111) );
  OAI22_X1 U3136 ( .A1(n17355), .A2(n15071), .B1(n17347), .B2(n16703), .ZN(
        n10112) );
  OAI22_X1 U3137 ( .A1(n17368), .A2(n15691), .B1(n17359), .B2(n16703), .ZN(
        n10113) );
  OAI22_X1 U3138 ( .A1(n17381), .A2(n14425), .B1(n17373), .B2(n16703), .ZN(
        n10114) );
  OAI22_X1 U3139 ( .A1(n17394), .A2(n14756), .B1(n17385), .B2(n16703), .ZN(
        n10115) );
  OAI22_X1 U3140 ( .A1(n17407), .A2(n14358), .B1(n17398), .B2(n16703), .ZN(
        n10116) );
  OAI22_X1 U3141 ( .A1(n17585), .A2(n14286), .B1(n17577), .B2(n16448), .ZN(
        n7911) );
  OAI22_X1 U3142 ( .A1(n17585), .A2(n14287), .B1(n17577), .B2(n16456), .ZN(
        n7985) );
  OAI22_X1 U3143 ( .A1(n16699), .A2(n14963), .B1(n16692), .B2(n16709), .ZN(
        n8055) );
  OAI22_X1 U3144 ( .A1(n16699), .A2(n14964), .B1(n16692), .B2(n16718), .ZN(
        n8057) );
  OAI22_X1 U3145 ( .A1(n16699), .A2(n14965), .B1(n16692), .B2(n16731), .ZN(
        n8061) );
  OAI22_X1 U3146 ( .A1(n16699), .A2(n14966), .B1(n16692), .B2(n16737), .ZN(
        n8063) );
  OAI22_X1 U3147 ( .A1(n17584), .A2(n14071), .B1(n17577), .B2(n16709), .ZN(
        n8113) );
  OAI22_X1 U3148 ( .A1(n17584), .A2(n14212), .B1(n17577), .B2(n16718), .ZN(
        n8185) );
  OAI22_X1 U3149 ( .A1(n16942), .A2(n14550), .B1(n16935), .B2(n16709), .ZN(
        n8118) );
  OAI22_X1 U3150 ( .A1(n17135), .A2(n15739), .B1(n17128), .B2(n16718), .ZN(
        n8198) );
  OAI22_X1 U3151 ( .A1(n16942), .A2(n14551), .B1(n16934), .B2(n16726), .ZN(
        n8278) );
  OAI22_X1 U3152 ( .A1(n17135), .A2(n15740), .B1(n17127), .B2(n16727), .ZN(
        n8294) );
  OAI22_X1 U3153 ( .A1(n16942), .A2(n14552), .B1(n16935), .B2(n16733), .ZN(
        n8350) );
  OAI22_X1 U3154 ( .A1(n17135), .A2(n15741), .B1(n17128), .B2(n16734), .ZN(
        n8366) );
  OAI22_X1 U3155 ( .A1(n16943), .A2(n14546), .B1(n16934), .B2(n16706), .ZN(
        n10078) );
  OAI22_X1 U3156 ( .A1(n17136), .A2(n15757), .B1(n17127), .B2(n16705), .ZN(
        n10094) );
  OAI22_X1 U3157 ( .A1(n18025), .A2(n14573), .B1(n18017), .B2(n16436), .ZN(
        n7769) );
  OAI22_X1 U3158 ( .A1(n18012), .A2(n12054), .B1(n18003), .B2(n16456), .ZN(
        n7990) );
  OAI22_X1 U3159 ( .A1(n18025), .A2(n14572), .B1(n18016), .B2(n16456), .ZN(
        n7991) );
  OAI22_X1 U3160 ( .A1(n18011), .A2(n12056), .B1(n18003), .B2(n16725), .ZN(
        n8270) );
  OAI22_X1 U3161 ( .A1(n18024), .A2(n14574), .B1(n18016), .B2(n16725), .ZN(
        n8271) );
  OAI22_X1 U3162 ( .A1(n18011), .A2(n12057), .B1(n18004), .B2(n16732), .ZN(
        n8342) );
  OAI22_X1 U3163 ( .A1(n17852), .A2(n18026), .B1(n17836), .B2(n14280), .ZN(
        n9990) );
  OAI22_X1 U3164 ( .A1(n17874), .A2(n18026), .B1(n17858), .B2(n14991), .ZN(
        n9991) );
  OAI22_X1 U3165 ( .A1(n17896), .A2(n18026), .B1(n17880), .B2(n15316), .ZN(
        n9992) );
  OAI22_X1 U3166 ( .A1(n17918), .A2(n18026), .B1(n17902), .B2(n14633), .ZN(
        n9993) );
  OAI22_X1 U3167 ( .A1(n17939), .A2(n18026), .B1(n17923), .B2(n15315), .ZN(
        n9994) );
  OAI22_X1 U3168 ( .A1(n17960), .A2(n18026), .B1(n17944), .B2(n14858), .ZN(
        n9995) );
  OAI22_X1 U3169 ( .A1(n17981), .A2(n18026), .B1(n17965), .B2(n15033), .ZN(
        n9996) );
  OAI22_X1 U3170 ( .A1(n17853), .A2(n16701), .B1(n17836), .B2(n14281), .ZN(
        n10062) );
  OAI22_X1 U3171 ( .A1(n17875), .A2(n16701), .B1(n17858), .B2(n14992), .ZN(
        n10063) );
  OAI22_X1 U3172 ( .A1(n17897), .A2(n16701), .B1(n17880), .B2(n15317), .ZN(
        n10064) );
  OAI22_X1 U3173 ( .A1(n17919), .A2(n16701), .B1(n17902), .B2(n14634), .ZN(
        n10065) );
  OAI22_X1 U3174 ( .A1(n17940), .A2(n16701), .B1(n17923), .B2(n14670), .ZN(
        n10066) );
  OAI22_X1 U3175 ( .A1(n17961), .A2(n16701), .B1(n17944), .B2(n14859), .ZN(
        n10067) );
  OAI22_X1 U3176 ( .A1(n17982), .A2(n16702), .B1(n17965), .B2(n15034), .ZN(
        n10068) );
  OAI22_X1 U3177 ( .A1(n16698), .A2(n14967), .B1(n16691), .B2(n16743), .ZN(
        n8065) );
  OAI22_X1 U3178 ( .A1(n16698), .A2(n14968), .B1(n16691), .B2(n16749), .ZN(
        n8067) );
  OAI22_X1 U3179 ( .A1(n16698), .A2(n14969), .B1(n16691), .B2(n16755), .ZN(
        n8069) );
  OAI22_X1 U3180 ( .A1(n16698), .A2(n14970), .B1(n16691), .B2(n16761), .ZN(
        n8071) );
  OAI22_X1 U3181 ( .A1(n16697), .A2(n14971), .B1(n16691), .B2(n16767), .ZN(
        n8073) );
  OAI22_X1 U3182 ( .A1(n16697), .A2(n14972), .B1(n16691), .B2(n16773), .ZN(
        n8075) );
  OAI22_X1 U3183 ( .A1(n16697), .A2(n14973), .B1(n16691), .B2(n16779), .ZN(
        n8077) );
  OAI22_X1 U3184 ( .A1(n16696), .A2(n14974), .B1(n16691), .B2(n16785), .ZN(
        n8079) );
  OAI22_X1 U3185 ( .A1(n16696), .A2(n14975), .B1(n16691), .B2(n16791), .ZN(
        n8081) );
  OAI22_X1 U3186 ( .A1(n16696), .A2(n14976), .B1(n16691), .B2(n16797), .ZN(
        n8083) );
  OAI22_X1 U3187 ( .A1(n16696), .A2(n14977), .B1(n16691), .B2(n16803), .ZN(
        n8085) );
  OAI22_X1 U3188 ( .A1(n16695), .A2(n14978), .B1(n16691), .B2(n16809), .ZN(
        n8087) );
  OAI22_X1 U3189 ( .A1(n16697), .A2(n14979), .B1(n16691), .B2(n16827), .ZN(
        n8093) );
  OAI22_X1 U3190 ( .A1(n17070), .A2(n15157), .B1(n17063), .B2(n16727), .ZN(
        n8289) );
  OAI22_X1 U3191 ( .A1(n17096), .A2(n15500), .B1(n17089), .B2(n16727), .ZN(
        n8291) );
  OAI22_X1 U3192 ( .A1(n17109), .A2(n11846), .B1(n17102), .B2(n16727), .ZN(
        n8292) );
  OAI22_X1 U3193 ( .A1(n17263), .A2(n14836), .B1(n17256), .B2(n16728), .ZN(
        n8305) );
  OAI22_X1 U3194 ( .A1(n17289), .A2(n14372), .B1(n17282), .B2(n16728), .ZN(
        n8307) );
  OAI22_X1 U3195 ( .A1(n17302), .A2(n14610), .B1(n17295), .B2(n16728), .ZN(
        n8308) );
  OAI22_X1 U3196 ( .A1(n17367), .A2(n15674), .B1(n17360), .B2(n16729), .ZN(
        n8313) );
  OAI22_X1 U3197 ( .A1(n17393), .A2(n14723), .B1(n17386), .B2(n16729), .ZN(
        n8315) );
  OAI22_X1 U3198 ( .A1(n17406), .A2(n14334), .B1(n17399), .B2(n16729), .ZN(
        n8316) );
  OAI22_X1 U3199 ( .A1(n17471), .A2(n15527), .B1(n17464), .B2(n16729), .ZN(
        n8321) );
  OAI22_X1 U3200 ( .A1(n17584), .A2(n14216), .B1(n17576), .B2(n16731), .ZN(
        n8329) );
  OAI22_X1 U3201 ( .A1(n18024), .A2(n14575), .B1(n18017), .B2(n16732), .ZN(
        n8343) );
  OAI22_X1 U3202 ( .A1(n17044), .A2(n15042), .B1(n17037), .B2(n16733), .ZN(
        n8359) );
  OAI22_X1 U3203 ( .A1(n17057), .A2(n14373), .B1(n17050), .B2(n16733), .ZN(
        n8360) );
  OAI22_X1 U3204 ( .A1(n17070), .A2(n15158), .B1(n17063), .B2(n16733), .ZN(
        n8361) );
  OAI22_X1 U3205 ( .A1(n17083), .A2(n15591), .B1(n17076), .B2(n16734), .ZN(
        n8362) );
  OAI22_X1 U3206 ( .A1(n17096), .A2(n15501), .B1(n17089), .B2(n16734), .ZN(
        n8363) );
  OAI22_X1 U3207 ( .A1(n17109), .A2(n11847), .B1(n17102), .B2(n16734), .ZN(
        n8364) );
  OAI22_X1 U3208 ( .A1(n17237), .A2(n15378), .B1(n17230), .B2(n16735), .ZN(
        n8375) );
  OAI22_X1 U3209 ( .A1(n17250), .A2(n12211), .B1(n17243), .B2(n16735), .ZN(
        n8376) );
  OAI22_X1 U3210 ( .A1(n17263), .A2(n14837), .B1(n17256), .B2(n16735), .ZN(
        n8377) );
  OAI22_X1 U3211 ( .A1(n17289), .A2(n14374), .B1(n17282), .B2(n16735), .ZN(
        n8379) );
  OAI22_X1 U3212 ( .A1(n17302), .A2(n14611), .B1(n17295), .B2(n16735), .ZN(
        n8380) );
  OAI22_X1 U3213 ( .A1(n17341), .A2(n11887), .B1(n17334), .B2(n16735), .ZN(
        n8383) );
  OAI22_X1 U3214 ( .A1(n17354), .A2(n15083), .B1(n17347), .B2(n16735), .ZN(
        n8384) );
  OAI22_X1 U3215 ( .A1(n17367), .A2(n15675), .B1(n17360), .B2(n16735), .ZN(
        n8385) );
  OAI22_X1 U3216 ( .A1(n17380), .A2(n14437), .B1(n17373), .B2(n16736), .ZN(
        n8386) );
  OAI22_X1 U3217 ( .A1(n17393), .A2(n14725), .B1(n17386), .B2(n16736), .ZN(
        n8387) );
  OAI22_X1 U3218 ( .A1(n17406), .A2(n14335), .B1(n17399), .B2(n16736), .ZN(
        n8388) );
  OAI22_X1 U3219 ( .A1(n17444), .A2(n12369), .B1(n17438), .B2(n16736), .ZN(
        n8391) );
  OAI22_X1 U3220 ( .A1(n17457), .A2(n14724), .B1(n17450), .B2(n16736), .ZN(
        n8392) );
  OAI22_X1 U3221 ( .A1(n17470), .A2(n15528), .B1(n17464), .B2(n16736), .ZN(
        n8393) );
  OAI22_X1 U3222 ( .A1(n17483), .A2(n15765), .B1(n17477), .B2(n16736), .ZN(
        n8394) );
  OAI22_X1 U3223 ( .A1(n17496), .A2(n14783), .B1(n17490), .B2(n16736), .ZN(
        n8395) );
  OAI22_X1 U3224 ( .A1(n17509), .A2(n15592), .B1(n17503), .B2(n16736), .ZN(
        n8396) );
  OAI22_X1 U3225 ( .A1(n17584), .A2(n14219), .B1(n17576), .B2(n16737), .ZN(
        n8401) );
  OAI22_X1 U3226 ( .A1(n18011), .A2(n12058), .B1(n18004), .B2(n16738), .ZN(
        n8414) );
  OAI22_X1 U3227 ( .A1(n18024), .A2(n14576), .B1(n18017), .B2(n16738), .ZN(
        n8415) );
  OAI22_X1 U3228 ( .A1(n16942), .A2(n14553), .B1(n16935), .B2(n16739), .ZN(
        n8422) );
  OAI22_X1 U3229 ( .A1(n17030), .A2(n12178), .B1(n17024), .B2(n16739), .ZN(
        n8430) );
  OAI22_X1 U3230 ( .A1(n17043), .A2(n15043), .B1(n17037), .B2(n16739), .ZN(
        n8431) );
  OAI22_X1 U3231 ( .A1(n17056), .A2(n14375), .B1(n17050), .B2(n16739), .ZN(
        n8432) );
  OAI22_X1 U3232 ( .A1(n17069), .A2(n15159), .B1(n17063), .B2(n16739), .ZN(
        n8433) );
  OAI22_X1 U3233 ( .A1(n17082), .A2(n15593), .B1(n17076), .B2(n16740), .ZN(
        n8434) );
  OAI22_X1 U3234 ( .A1(n17095), .A2(n15502), .B1(n17089), .B2(n16740), .ZN(
        n8435) );
  OAI22_X1 U3235 ( .A1(n17108), .A2(n11849), .B1(n17102), .B2(n16740), .ZN(
        n8436) );
  OAI22_X1 U3236 ( .A1(n17135), .A2(n15742), .B1(n17128), .B2(n16740), .ZN(
        n8438) );
  OAI22_X1 U3237 ( .A1(n17236), .A2(n15379), .B1(n17230), .B2(n16741), .ZN(
        n8447) );
  OAI22_X1 U3238 ( .A1(n17249), .A2(n12212), .B1(n17243), .B2(n16741), .ZN(
        n8448) );
  OAI22_X1 U3239 ( .A1(n17262), .A2(n14838), .B1(n17256), .B2(n16741), .ZN(
        n8449) );
  OAI22_X1 U3240 ( .A1(n17288), .A2(n14376), .B1(n17282), .B2(n16741), .ZN(
        n8451) );
  OAI22_X1 U3241 ( .A1(n17301), .A2(n14612), .B1(n17295), .B2(n16741), .ZN(
        n8452) );
  OAI22_X1 U3242 ( .A1(n17327), .A2(n15299), .B1(n17321), .B2(n16741), .ZN(
        n8454) );
  OAI22_X1 U3243 ( .A1(n17340), .A2(n11888), .B1(n17334), .B2(n16741), .ZN(
        n8455) );
  OAI22_X1 U3244 ( .A1(n17353), .A2(n15085), .B1(n17347), .B2(n16741), .ZN(
        n8456) );
  OAI22_X1 U3245 ( .A1(n17366), .A2(n15676), .B1(n17360), .B2(n16741), .ZN(
        n8457) );
  OAI22_X1 U3246 ( .A1(n17379), .A2(n14439), .B1(n17373), .B2(n16742), .ZN(
        n8458) );
  OAI22_X1 U3247 ( .A1(n17392), .A2(n14727), .B1(n17386), .B2(n16742), .ZN(
        n8459) );
  OAI22_X1 U3248 ( .A1(n17405), .A2(n14336), .B1(n17399), .B2(n16742), .ZN(
        n8460) );
  OAI22_X1 U3249 ( .A1(n17431), .A2(n15334), .B1(n17425), .B2(n16742), .ZN(
        n8462) );
  OAI22_X1 U3250 ( .A1(n17444), .A2(n12408), .B1(n17438), .B2(n16742), .ZN(
        n8463) );
  OAI22_X1 U3251 ( .A1(n17457), .A2(n14726), .B1(n17450), .B2(n16742), .ZN(
        n8464) );
  OAI22_X1 U3252 ( .A1(n17470), .A2(n15529), .B1(n17464), .B2(n16742), .ZN(
        n8465) );
  OAI22_X1 U3253 ( .A1(n17483), .A2(n15766), .B1(n17477), .B2(n16742), .ZN(
        n8466) );
  OAI22_X1 U3254 ( .A1(n17496), .A2(n14785), .B1(n17490), .B2(n16742), .ZN(
        n8467) );
  OAI22_X1 U3255 ( .A1(n17509), .A2(n15594), .B1(n17503), .B2(n16742), .ZN(
        n8468) );
  OAI22_X1 U3256 ( .A1(n17583), .A2(n14225), .B1(n17576), .B2(n16743), .ZN(
        n8473) );
  OAI22_X1 U3257 ( .A1(n18011), .A2(n12059), .B1(n18004), .B2(n16744), .ZN(
        n8486) );
  OAI22_X1 U3258 ( .A1(n18024), .A2(n14577), .B1(n18017), .B2(n16744), .ZN(
        n8487) );
  OAI22_X1 U3259 ( .A1(n16941), .A2(n14554), .B1(n16935), .B2(n16745), .ZN(
        n8494) );
  OAI22_X1 U3260 ( .A1(n17030), .A2(n12179), .B1(n17024), .B2(n16745), .ZN(
        n8502) );
  OAI22_X1 U3261 ( .A1(n17043), .A2(n15044), .B1(n17037), .B2(n16745), .ZN(
        n8503) );
  OAI22_X1 U3262 ( .A1(n17056), .A2(n14377), .B1(n17050), .B2(n16745), .ZN(
        n8504) );
  OAI22_X1 U3263 ( .A1(n17069), .A2(n15160), .B1(n17063), .B2(n16745), .ZN(
        n8505) );
  OAI22_X1 U3264 ( .A1(n17082), .A2(n15595), .B1(n17076), .B2(n16746), .ZN(
        n8506) );
  OAI22_X1 U3265 ( .A1(n17095), .A2(n15503), .B1(n17089), .B2(n16746), .ZN(
        n8507) );
  OAI22_X1 U3266 ( .A1(n17108), .A2(n11850), .B1(n17102), .B2(n16746), .ZN(
        n8508) );
  OAI22_X1 U3267 ( .A1(n17134), .A2(n15743), .B1(n17128), .B2(n16746), .ZN(
        n8510) );
  OAI22_X1 U3268 ( .A1(n17236), .A2(n15380), .B1(n17230), .B2(n16747), .ZN(
        n8519) );
  OAI22_X1 U3269 ( .A1(n17249), .A2(n12213), .B1(n17243), .B2(n16747), .ZN(
        n8520) );
  OAI22_X1 U3270 ( .A1(n17262), .A2(n14839), .B1(n17256), .B2(n16747), .ZN(
        n8521) );
  OAI22_X1 U3271 ( .A1(n17288), .A2(n14378), .B1(n17282), .B2(n16747), .ZN(
        n8523) );
  OAI22_X1 U3272 ( .A1(n17301), .A2(n14613), .B1(n17295), .B2(n16747), .ZN(
        n8524) );
  OAI22_X1 U3273 ( .A1(n17327), .A2(n15300), .B1(n17321), .B2(n16747), .ZN(
        n8526) );
  OAI22_X1 U3274 ( .A1(n17340), .A2(n11889), .B1(n17334), .B2(n16747), .ZN(
        n8527) );
  OAI22_X1 U3275 ( .A1(n17353), .A2(n15087), .B1(n17347), .B2(n16747), .ZN(
        n8528) );
  OAI22_X1 U3276 ( .A1(n17366), .A2(n15677), .B1(n17360), .B2(n16747), .ZN(
        n8529) );
  OAI22_X1 U3277 ( .A1(n17379), .A2(n14441), .B1(n17373), .B2(n16748), .ZN(
        n8530) );
  OAI22_X1 U3278 ( .A1(n17392), .A2(n14729), .B1(n17386), .B2(n16748), .ZN(
        n8531) );
  OAI22_X1 U3279 ( .A1(n17405), .A2(n14337), .B1(n17399), .B2(n16748), .ZN(
        n8532) );
  OAI22_X1 U3280 ( .A1(n17431), .A2(n15335), .B1(n17425), .B2(n16748), .ZN(
        n8534) );
  OAI22_X1 U3281 ( .A1(n17444), .A2(n12410), .B1(n17438), .B2(n16748), .ZN(
        n8535) );
  OAI22_X1 U3282 ( .A1(n17457), .A2(n14728), .B1(n17450), .B2(n16748), .ZN(
        n8536) );
  OAI22_X1 U3283 ( .A1(n17470), .A2(n15530), .B1(n17464), .B2(n16748), .ZN(
        n8537) );
  OAI22_X1 U3284 ( .A1(n17483), .A2(n15767), .B1(n17477), .B2(n16748), .ZN(
        n8538) );
  OAI22_X1 U3285 ( .A1(n17496), .A2(n14787), .B1(n17490), .B2(n16748), .ZN(
        n8539) );
  OAI22_X1 U3286 ( .A1(n17509), .A2(n15596), .B1(n17503), .B2(n16748), .ZN(
        n8540) );
  OAI22_X1 U3287 ( .A1(n17583), .A2(n14227), .B1(n17576), .B2(n16749), .ZN(
        n8545) );
  OAI22_X1 U3288 ( .A1(n18010), .A2(n12060), .B1(n18004), .B2(n16750), .ZN(
        n8558) );
  OAI22_X1 U3289 ( .A1(n18023), .A2(n14578), .B1(n18017), .B2(n16750), .ZN(
        n8559) );
  OAI22_X1 U3290 ( .A1(n16941), .A2(n14555), .B1(n16935), .B2(n16751), .ZN(
        n8566) );
  OAI22_X1 U3291 ( .A1(n17030), .A2(n12180), .B1(n17024), .B2(n16751), .ZN(
        n8574) );
  OAI22_X1 U3292 ( .A1(n17043), .A2(n15045), .B1(n17037), .B2(n16751), .ZN(
        n8575) );
  OAI22_X1 U3293 ( .A1(n17056), .A2(n14379), .B1(n17050), .B2(n16751), .ZN(
        n8576) );
  OAI22_X1 U3294 ( .A1(n17069), .A2(n15161), .B1(n17063), .B2(n16751), .ZN(
        n8577) );
  OAI22_X1 U3295 ( .A1(n17082), .A2(n15597), .B1(n17076), .B2(n16752), .ZN(
        n8578) );
  OAI22_X1 U3296 ( .A1(n17095), .A2(n15504), .B1(n17089), .B2(n16752), .ZN(
        n8579) );
  OAI22_X1 U3297 ( .A1(n17108), .A2(n11851), .B1(n17102), .B2(n16752), .ZN(
        n8580) );
  OAI22_X1 U3298 ( .A1(n17134), .A2(n15744), .B1(n17128), .B2(n16752), .ZN(
        n8582) );
  OAI22_X1 U3299 ( .A1(n17236), .A2(n15381), .B1(n17230), .B2(n16753), .ZN(
        n8591) );
  OAI22_X1 U3300 ( .A1(n17249), .A2(n12214), .B1(n17243), .B2(n16753), .ZN(
        n8592) );
  OAI22_X1 U3301 ( .A1(n17262), .A2(n14840), .B1(n17256), .B2(n16753), .ZN(
        n8593) );
  OAI22_X1 U3302 ( .A1(n17288), .A2(n14380), .B1(n17282), .B2(n16753), .ZN(
        n8595) );
  OAI22_X1 U3303 ( .A1(n17301), .A2(n14614), .B1(n17295), .B2(n16753), .ZN(
        n8596) );
  OAI22_X1 U3304 ( .A1(n17327), .A2(n15301), .B1(n17321), .B2(n16753), .ZN(
        n8598) );
  OAI22_X1 U3305 ( .A1(n17340), .A2(n11890), .B1(n17334), .B2(n16753), .ZN(
        n8599) );
  OAI22_X1 U3306 ( .A1(n17353), .A2(n15089), .B1(n17347), .B2(n16753), .ZN(
        n8600) );
  OAI22_X1 U3307 ( .A1(n17366), .A2(n15678), .B1(n17360), .B2(n16753), .ZN(
        n8601) );
  OAI22_X1 U3308 ( .A1(n17379), .A2(n14443), .B1(n17373), .B2(n16754), .ZN(
        n8602) );
  OAI22_X1 U3309 ( .A1(n17392), .A2(n14731), .B1(n17386), .B2(n16754), .ZN(
        n8603) );
  OAI22_X1 U3310 ( .A1(n17405), .A2(n14338), .B1(n17399), .B2(n16754), .ZN(
        n8604) );
  OAI22_X1 U3311 ( .A1(n17431), .A2(n15336), .B1(n17425), .B2(n16754), .ZN(
        n8606) );
  OAI22_X1 U3312 ( .A1(n17444), .A2(n12551), .B1(n17438), .B2(n16754), .ZN(
        n8607) );
  OAI22_X1 U3313 ( .A1(n17457), .A2(n14730), .B1(n17450), .B2(n16754), .ZN(
        n8608) );
  OAI22_X1 U3314 ( .A1(n17470), .A2(n15531), .B1(n17464), .B2(n16754), .ZN(
        n8609) );
  OAI22_X1 U3315 ( .A1(n17483), .A2(n15768), .B1(n17477), .B2(n16754), .ZN(
        n8610) );
  OAI22_X1 U3316 ( .A1(n17496), .A2(n14789), .B1(n17490), .B2(n16754), .ZN(
        n8611) );
  OAI22_X1 U3317 ( .A1(n17509), .A2(n15598), .B1(n17503), .B2(n16754), .ZN(
        n8612) );
  OAI22_X1 U3318 ( .A1(n17583), .A2(n14230), .B1(n17576), .B2(n16755), .ZN(
        n8617) );
  OAI22_X1 U3319 ( .A1(n18010), .A2(n12098), .B1(n18004), .B2(n16756), .ZN(
        n8630) );
  OAI22_X1 U3320 ( .A1(n18023), .A2(n14579), .B1(n18017), .B2(n16756), .ZN(
        n8631) );
  OAI22_X1 U3321 ( .A1(n16941), .A2(n14556), .B1(n16935), .B2(n16757), .ZN(
        n8638) );
  OAI22_X1 U3322 ( .A1(n17030), .A2(n12181), .B1(n17024), .B2(n16757), .ZN(
        n8646) );
  OAI22_X1 U3323 ( .A1(n17043), .A2(n15046), .B1(n17037), .B2(n16757), .ZN(
        n8647) );
  OAI22_X1 U3324 ( .A1(n17056), .A2(n14381), .B1(n17050), .B2(n16757), .ZN(
        n8648) );
  OAI22_X1 U3325 ( .A1(n17069), .A2(n15162), .B1(n17063), .B2(n16757), .ZN(
        n8649) );
  OAI22_X1 U3326 ( .A1(n17082), .A2(n15599), .B1(n17076), .B2(n16758), .ZN(
        n8650) );
  OAI22_X1 U3327 ( .A1(n17095), .A2(n15505), .B1(n17089), .B2(n16758), .ZN(
        n8651) );
  OAI22_X1 U3328 ( .A1(n17108), .A2(n11852), .B1(n17102), .B2(n16758), .ZN(
        n8652) );
  OAI22_X1 U3329 ( .A1(n17134), .A2(n15745), .B1(n17128), .B2(n16758), .ZN(
        n8654) );
  OAI22_X1 U3330 ( .A1(n17236), .A2(n15382), .B1(n17230), .B2(n16759), .ZN(
        n8663) );
  OAI22_X1 U3331 ( .A1(n17249), .A2(n12215), .B1(n17243), .B2(n16759), .ZN(
        n8664) );
  OAI22_X1 U3332 ( .A1(n17262), .A2(n14841), .B1(n17256), .B2(n16759), .ZN(
        n8665) );
  OAI22_X1 U3333 ( .A1(n17288), .A2(n14382), .B1(n17282), .B2(n16759), .ZN(
        n8667) );
  OAI22_X1 U3334 ( .A1(n17301), .A2(n14615), .B1(n17295), .B2(n16759), .ZN(
        n8668) );
  OAI22_X1 U3335 ( .A1(n17327), .A2(n15302), .B1(n17321), .B2(n16759), .ZN(
        n8670) );
  OAI22_X1 U3336 ( .A1(n17340), .A2(n11891), .B1(n17334), .B2(n16759), .ZN(
        n8671) );
  OAI22_X1 U3337 ( .A1(n17353), .A2(n15091), .B1(n17347), .B2(n16759), .ZN(
        n8672) );
  OAI22_X1 U3338 ( .A1(n17366), .A2(n15679), .B1(n17360), .B2(n16759), .ZN(
        n8673) );
  OAI22_X1 U3339 ( .A1(n17379), .A2(n14445), .B1(n17373), .B2(n16760), .ZN(
        n8674) );
  OAI22_X1 U3340 ( .A1(n17392), .A2(n14733), .B1(n17386), .B2(n16760), .ZN(
        n8675) );
  OAI22_X1 U3341 ( .A1(n17405), .A2(n14339), .B1(n17399), .B2(n16760), .ZN(
        n8676) );
  OAI22_X1 U3342 ( .A1(n17430), .A2(n15337), .B1(n17425), .B2(n16760), .ZN(
        n8678) );
  OAI22_X1 U3343 ( .A1(n17443), .A2(n12602), .B1(n17438), .B2(n16760), .ZN(
        n8679) );
  OAI22_X1 U3344 ( .A1(n17456), .A2(n14732), .B1(n17450), .B2(n16760), .ZN(
        n8680) );
  OAI22_X1 U3345 ( .A1(n17469), .A2(n15532), .B1(n17464), .B2(n16760), .ZN(
        n8681) );
  OAI22_X1 U3346 ( .A1(n17482), .A2(n15769), .B1(n17477), .B2(n16760), .ZN(
        n8682) );
  OAI22_X1 U3347 ( .A1(n17495), .A2(n14791), .B1(n17490), .B2(n16760), .ZN(
        n8683) );
  OAI22_X1 U3348 ( .A1(n17508), .A2(n15600), .B1(n17503), .B2(n16760), .ZN(
        n8684) );
  OAI22_X1 U3349 ( .A1(n17583), .A2(n14235), .B1(n17576), .B2(n16761), .ZN(
        n8689) );
  OAI22_X1 U3350 ( .A1(n18010), .A2(n12099), .B1(n18004), .B2(n16762), .ZN(
        n8702) );
  OAI22_X1 U3351 ( .A1(n18023), .A2(n14580), .B1(n18017), .B2(n16762), .ZN(
        n8703) );
  OAI22_X1 U3352 ( .A1(n16941), .A2(n14557), .B1(n16935), .B2(n16763), .ZN(
        n8710) );
  OAI22_X1 U3353 ( .A1(n17029), .A2(n12182), .B1(n17024), .B2(n16763), .ZN(
        n8718) );
  OAI22_X1 U3354 ( .A1(n17042), .A2(n15047), .B1(n17037), .B2(n16763), .ZN(
        n8719) );
  OAI22_X1 U3355 ( .A1(n17055), .A2(n14383), .B1(n17050), .B2(n16763), .ZN(
        n8720) );
  OAI22_X1 U3356 ( .A1(n17068), .A2(n15163), .B1(n17063), .B2(n16763), .ZN(
        n8721) );
  OAI22_X1 U3357 ( .A1(n17081), .A2(n15601), .B1(n17076), .B2(n16764), .ZN(
        n8722) );
  OAI22_X1 U3358 ( .A1(n17094), .A2(n15506), .B1(n17089), .B2(n16764), .ZN(
        n8723) );
  OAI22_X1 U3359 ( .A1(n17107), .A2(n11854), .B1(n17102), .B2(n16764), .ZN(
        n8724) );
  OAI22_X1 U3360 ( .A1(n17134), .A2(n15746), .B1(n17128), .B2(n16764), .ZN(
        n8726) );
  OAI22_X1 U3361 ( .A1(n17235), .A2(n15383), .B1(n17230), .B2(n16765), .ZN(
        n8735) );
  OAI22_X1 U3362 ( .A1(n17248), .A2(n12253), .B1(n17243), .B2(n16765), .ZN(
        n8736) );
  OAI22_X1 U3363 ( .A1(n17261), .A2(n14842), .B1(n17256), .B2(n16765), .ZN(
        n8737) );
  OAI22_X1 U3364 ( .A1(n17287), .A2(n14384), .B1(n17282), .B2(n16765), .ZN(
        n8739) );
  OAI22_X1 U3365 ( .A1(n17300), .A2(n14616), .B1(n17295), .B2(n16765), .ZN(
        n8740) );
  OAI22_X1 U3366 ( .A1(n17326), .A2(n15303), .B1(n17321), .B2(n16765), .ZN(
        n8742) );
  OAI22_X1 U3367 ( .A1(n17339), .A2(n11892), .B1(n17334), .B2(n16765), .ZN(
        n8743) );
  OAI22_X1 U3368 ( .A1(n17352), .A2(n15093), .B1(n17347), .B2(n16765), .ZN(
        n8744) );
  OAI22_X1 U3369 ( .A1(n17365), .A2(n15680), .B1(n17360), .B2(n16765), .ZN(
        n8745) );
  OAI22_X1 U3370 ( .A1(n17378), .A2(n14447), .B1(n17373), .B2(n16766), .ZN(
        n8746) );
  OAI22_X1 U3371 ( .A1(n17391), .A2(n14735), .B1(n17386), .B2(n16766), .ZN(
        n8747) );
  OAI22_X1 U3372 ( .A1(n17404), .A2(n14340), .B1(n17399), .B2(n16766), .ZN(
        n8748) );
  OAI22_X1 U3373 ( .A1(n17430), .A2(n15338), .B1(n17425), .B2(n16766), .ZN(
        n8750) );
  OAI22_X1 U3374 ( .A1(n17443), .A2(n12669), .B1(n17438), .B2(n16766), .ZN(
        n8751) );
  OAI22_X1 U3375 ( .A1(n17456), .A2(n14734), .B1(n17450), .B2(n16766), .ZN(
        n8752) );
  OAI22_X1 U3376 ( .A1(n17469), .A2(n15533), .B1(n17464), .B2(n16766), .ZN(
        n8753) );
  OAI22_X1 U3377 ( .A1(n17482), .A2(n15770), .B1(n17477), .B2(n16766), .ZN(
        n8754) );
  OAI22_X1 U3378 ( .A1(n17495), .A2(n14793), .B1(n17490), .B2(n16766), .ZN(
        n8755) );
  OAI22_X1 U3379 ( .A1(n17508), .A2(n15602), .B1(n17503), .B2(n16766), .ZN(
        n8756) );
  OAI22_X1 U3380 ( .A1(n17582), .A2(n14242), .B1(n17576), .B2(n16767), .ZN(
        n8761) );
  OAI22_X1 U3381 ( .A1(n18010), .A2(n12100), .B1(n18004), .B2(n16768), .ZN(
        n8774) );
  OAI22_X1 U3382 ( .A1(n18023), .A2(n14581), .B1(n18017), .B2(n16768), .ZN(
        n8775) );
  OAI22_X1 U3383 ( .A1(n16940), .A2(n14558), .B1(n16935), .B2(n16769), .ZN(
        n8782) );
  OAI22_X1 U3384 ( .A1(n17029), .A2(n12183), .B1(n17024), .B2(n16769), .ZN(
        n8790) );
  OAI22_X1 U3385 ( .A1(n17042), .A2(n15048), .B1(n17037), .B2(n16769), .ZN(
        n8791) );
  OAI22_X1 U3386 ( .A1(n17055), .A2(n14385), .B1(n17050), .B2(n16769), .ZN(
        n8792) );
  OAI22_X1 U3387 ( .A1(n17068), .A2(n15164), .B1(n17063), .B2(n16769), .ZN(
        n8793) );
  OAI22_X1 U3388 ( .A1(n17081), .A2(n15603), .B1(n17076), .B2(n16770), .ZN(
        n8794) );
  OAI22_X1 U3389 ( .A1(n17094), .A2(n15507), .B1(n17089), .B2(n16770), .ZN(
        n8795) );
  OAI22_X1 U3390 ( .A1(n17107), .A2(n11855), .B1(n17102), .B2(n16770), .ZN(
        n8796) );
  OAI22_X1 U3391 ( .A1(n17133), .A2(n15747), .B1(n17128), .B2(n16770), .ZN(
        n8798) );
  OAI22_X1 U3392 ( .A1(n17235), .A2(n15384), .B1(n17230), .B2(n16771), .ZN(
        n8807) );
  OAI22_X1 U3393 ( .A1(n17248), .A2(n12254), .B1(n17243), .B2(n16771), .ZN(
        n8808) );
  OAI22_X1 U3394 ( .A1(n17261), .A2(n14843), .B1(n17256), .B2(n16771), .ZN(
        n8809) );
  OAI22_X1 U3395 ( .A1(n17287), .A2(n14386), .B1(n17282), .B2(n16771), .ZN(
        n8811) );
  OAI22_X1 U3396 ( .A1(n17300), .A2(n14617), .B1(n17295), .B2(n16771), .ZN(
        n8812) );
  OAI22_X1 U3397 ( .A1(n17326), .A2(n15304), .B1(n17321), .B2(n16771), .ZN(
        n8814) );
  OAI22_X1 U3398 ( .A1(n17339), .A2(n11893), .B1(n17334), .B2(n16771), .ZN(
        n8815) );
  OAI22_X1 U3399 ( .A1(n17352), .A2(n15095), .B1(n17347), .B2(n16771), .ZN(
        n8816) );
  OAI22_X1 U3400 ( .A1(n17365), .A2(n15681), .B1(n17360), .B2(n16771), .ZN(
        n8817) );
  OAI22_X1 U3401 ( .A1(n17378), .A2(n14449), .B1(n17373), .B2(n16772), .ZN(
        n8818) );
  OAI22_X1 U3402 ( .A1(n17391), .A2(n14737), .B1(n17386), .B2(n16772), .ZN(
        n8819) );
  OAI22_X1 U3403 ( .A1(n17404), .A2(n14341), .B1(n17399), .B2(n16772), .ZN(
        n8820) );
  OAI22_X1 U3404 ( .A1(n17430), .A2(n15339), .B1(n17425), .B2(n16772), .ZN(
        n8822) );
  OAI22_X1 U3405 ( .A1(n17443), .A2(n13999), .B1(n17438), .B2(n16772), .ZN(
        n8823) );
  OAI22_X1 U3406 ( .A1(n17456), .A2(n14736), .B1(n17450), .B2(n16772), .ZN(
        n8824) );
  OAI22_X1 U3407 ( .A1(n17469), .A2(n15534), .B1(n17464), .B2(n16772), .ZN(
        n8825) );
  OAI22_X1 U3408 ( .A1(n17482), .A2(n15771), .B1(n17477), .B2(n16772), .ZN(
        n8826) );
  OAI22_X1 U3409 ( .A1(n17495), .A2(n14795), .B1(n17490), .B2(n16772), .ZN(
        n8827) );
  OAI22_X1 U3410 ( .A1(n17508), .A2(n15604), .B1(n17503), .B2(n16772), .ZN(
        n8828) );
  OAI22_X1 U3411 ( .A1(n17582), .A2(n14243), .B1(n17576), .B2(n16773), .ZN(
        n8833) );
  OAI22_X1 U3412 ( .A1(n18009), .A2(n12101), .B1(n18004), .B2(n16774), .ZN(
        n8846) );
  OAI22_X1 U3413 ( .A1(n18022), .A2(n14582), .B1(n18017), .B2(n16774), .ZN(
        n8847) );
  OAI22_X1 U3414 ( .A1(n16940), .A2(n14559), .B1(n16935), .B2(n16775), .ZN(
        n8854) );
  OAI22_X1 U3415 ( .A1(n17029), .A2(n12185), .B1(n17024), .B2(n16775), .ZN(
        n8862) );
  OAI22_X1 U3416 ( .A1(n17042), .A2(n15049), .B1(n17037), .B2(n16775), .ZN(
        n8863) );
  OAI22_X1 U3417 ( .A1(n17055), .A2(n14387), .B1(n17050), .B2(n16775), .ZN(
        n8864) );
  OAI22_X1 U3418 ( .A1(n17068), .A2(n15165), .B1(n17063), .B2(n16775), .ZN(
        n8865) );
  OAI22_X1 U3419 ( .A1(n17081), .A2(n15605), .B1(n17076), .B2(n16776), .ZN(
        n8866) );
  OAI22_X1 U3420 ( .A1(n17094), .A2(n15508), .B1(n17089), .B2(n16776), .ZN(
        n8867) );
  OAI22_X1 U3421 ( .A1(n17107), .A2(n11856), .B1(n17102), .B2(n16776), .ZN(
        n8868) );
  OAI22_X1 U3422 ( .A1(n17133), .A2(n15748), .B1(n17128), .B2(n16776), .ZN(
        n8870) );
  OAI22_X1 U3423 ( .A1(n17235), .A2(n15385), .B1(n17230), .B2(n16777), .ZN(
        n8879) );
  OAI22_X1 U3424 ( .A1(n17248), .A2(n12255), .B1(n17243), .B2(n16777), .ZN(
        n8880) );
  OAI22_X1 U3425 ( .A1(n17261), .A2(n14844), .B1(n17256), .B2(n16777), .ZN(
        n8881) );
  OAI22_X1 U3426 ( .A1(n17287), .A2(n14388), .B1(n17282), .B2(n16777), .ZN(
        n8883) );
  OAI22_X1 U3427 ( .A1(n17300), .A2(n14618), .B1(n17295), .B2(n16777), .ZN(
        n8884) );
  OAI22_X1 U3428 ( .A1(n17326), .A2(n15305), .B1(n17321), .B2(n16777), .ZN(
        n8886) );
  OAI22_X1 U3429 ( .A1(n17339), .A2(n11894), .B1(n17334), .B2(n16777), .ZN(
        n8887) );
  OAI22_X1 U3430 ( .A1(n17352), .A2(n15097), .B1(n17347), .B2(n16777), .ZN(
        n8888) );
  OAI22_X1 U3431 ( .A1(n17365), .A2(n15682), .B1(n17360), .B2(n16777), .ZN(
        n8889) );
  OAI22_X1 U3432 ( .A1(n17378), .A2(n14451), .B1(n17373), .B2(n16778), .ZN(
        n8890) );
  OAI22_X1 U3433 ( .A1(n17391), .A2(n14739), .B1(n17386), .B2(n16778), .ZN(
        n8891) );
  OAI22_X1 U3434 ( .A1(n17404), .A2(n14342), .B1(n17399), .B2(n16778), .ZN(
        n8892) );
  OAI22_X1 U3435 ( .A1(n17429), .A2(n15340), .B1(n17425), .B2(n16778), .ZN(
        n8894) );
  OAI22_X1 U3436 ( .A1(n17442), .A2(n14014), .B1(n17438), .B2(n16778), .ZN(
        n8895) );
  OAI22_X1 U3437 ( .A1(n17455), .A2(n14738), .B1(n17450), .B2(n16778), .ZN(
        n8896) );
  OAI22_X1 U3438 ( .A1(n17468), .A2(n15535), .B1(n17464), .B2(n16778), .ZN(
        n8897) );
  OAI22_X1 U3439 ( .A1(n17481), .A2(n15772), .B1(n17477), .B2(n16778), .ZN(
        n8898) );
  OAI22_X1 U3440 ( .A1(n17494), .A2(n14797), .B1(n17490), .B2(n16778), .ZN(
        n8899) );
  OAI22_X1 U3441 ( .A1(n17507), .A2(n15606), .B1(n17503), .B2(n16778), .ZN(
        n8900) );
  OAI22_X1 U3442 ( .A1(n17582), .A2(n14246), .B1(n17576), .B2(n16779), .ZN(
        n8905) );
  OAI22_X1 U3443 ( .A1(n18009), .A2(n12102), .B1(n18004), .B2(n16780), .ZN(
        n8918) );
  OAI22_X1 U3444 ( .A1(n18022), .A2(n14583), .B1(n18017), .B2(n16780), .ZN(
        n8919) );
  OAI22_X1 U3445 ( .A1(n16940), .A2(n14560), .B1(n16935), .B2(n16781), .ZN(
        n8926) );
  OAI22_X1 U3446 ( .A1(n17028), .A2(n12186), .B1(n17024), .B2(n16781), .ZN(
        n8934) );
  OAI22_X1 U3447 ( .A1(n17041), .A2(n15050), .B1(n17037), .B2(n16781), .ZN(
        n8935) );
  OAI22_X1 U3448 ( .A1(n17054), .A2(n14389), .B1(n17050), .B2(n16781), .ZN(
        n8936) );
  OAI22_X1 U3449 ( .A1(n17067), .A2(n15166), .B1(n17063), .B2(n16781), .ZN(
        n8937) );
  OAI22_X1 U3450 ( .A1(n17080), .A2(n15607), .B1(n17076), .B2(n16782), .ZN(
        n8938) );
  OAI22_X1 U3451 ( .A1(n17093), .A2(n15509), .B1(n17089), .B2(n16782), .ZN(
        n8939) );
  OAI22_X1 U3452 ( .A1(n17106), .A2(n11857), .B1(n17102), .B2(n16782), .ZN(
        n8940) );
  OAI22_X1 U3453 ( .A1(n17133), .A2(n15749), .B1(n17128), .B2(n16782), .ZN(
        n8942) );
  OAI22_X1 U3454 ( .A1(n17234), .A2(n15386), .B1(n17230), .B2(n16783), .ZN(
        n8951) );
  OAI22_X1 U3455 ( .A1(n17247), .A2(n12256), .B1(n17243), .B2(n16783), .ZN(
        n8952) );
  OAI22_X1 U3456 ( .A1(n17260), .A2(n14845), .B1(n17256), .B2(n16783), .ZN(
        n8953) );
  OAI22_X1 U3457 ( .A1(n17286), .A2(n14390), .B1(n17282), .B2(n16783), .ZN(
        n8955) );
  OAI22_X1 U3458 ( .A1(n17299), .A2(n14619), .B1(n17295), .B2(n16783), .ZN(
        n8956) );
  OAI22_X1 U3459 ( .A1(n17325), .A2(n15306), .B1(n17321), .B2(n16783), .ZN(
        n8958) );
  OAI22_X1 U3460 ( .A1(n17338), .A2(n11895), .B1(n17334), .B2(n16783), .ZN(
        n8959) );
  OAI22_X1 U3461 ( .A1(n17351), .A2(n15099), .B1(n17347), .B2(n16783), .ZN(
        n8960) );
  OAI22_X1 U3462 ( .A1(n17364), .A2(n15683), .B1(n17360), .B2(n16783), .ZN(
        n8961) );
  OAI22_X1 U3463 ( .A1(n17377), .A2(n14453), .B1(n17373), .B2(n16784), .ZN(
        n8962) );
  OAI22_X1 U3464 ( .A1(n17390), .A2(n14741), .B1(n17386), .B2(n16784), .ZN(
        n8963) );
  OAI22_X1 U3465 ( .A1(n17403), .A2(n14343), .B1(n17399), .B2(n16784), .ZN(
        n8964) );
  OAI22_X1 U3466 ( .A1(n17429), .A2(n15341), .B1(n17425), .B2(n16784), .ZN(
        n8966) );
  OAI22_X1 U3467 ( .A1(n17442), .A2(n14032), .B1(n17438), .B2(n16784), .ZN(
        n8967) );
  OAI22_X1 U3468 ( .A1(n17455), .A2(n14740), .B1(n17450), .B2(n16784), .ZN(
        n8968) );
  OAI22_X1 U3469 ( .A1(n17468), .A2(n15536), .B1(n17464), .B2(n16784), .ZN(
        n8969) );
  OAI22_X1 U3470 ( .A1(n17481), .A2(n15773), .B1(n17477), .B2(n16784), .ZN(
        n8970) );
  OAI22_X1 U3471 ( .A1(n17494), .A2(n14799), .B1(n17490), .B2(n16784), .ZN(
        n8971) );
  OAI22_X1 U3472 ( .A1(n17507), .A2(n15608), .B1(n17503), .B2(n16784), .ZN(
        n8972) );
  OAI22_X1 U3473 ( .A1(n17581), .A2(n14255), .B1(n17576), .B2(n16785), .ZN(
        n8977) );
  OAI22_X1 U3474 ( .A1(n18009), .A2(n12103), .B1(n18004), .B2(n16786), .ZN(
        n8990) );
  OAI22_X1 U3475 ( .A1(n18022), .A2(n14584), .B1(n18017), .B2(n16786), .ZN(
        n8991) );
  OAI22_X1 U3476 ( .A1(n16939), .A2(n14561), .B1(n16935), .B2(n16787), .ZN(
        n8998) );
  OAI22_X1 U3477 ( .A1(n17028), .A2(n12187), .B1(n17024), .B2(n16787), .ZN(
        n9006) );
  OAI22_X1 U3478 ( .A1(n17041), .A2(n15051), .B1(n17037), .B2(n16787), .ZN(
        n9007) );
  OAI22_X1 U3479 ( .A1(n17054), .A2(n14391), .B1(n17050), .B2(n16787), .ZN(
        n9008) );
  OAI22_X1 U3480 ( .A1(n17067), .A2(n15167), .B1(n17063), .B2(n16787), .ZN(
        n9009) );
  OAI22_X1 U3481 ( .A1(n17080), .A2(n15609), .B1(n17076), .B2(n16788), .ZN(
        n9010) );
  OAI22_X1 U3482 ( .A1(n17093), .A2(n15510), .B1(n17089), .B2(n16788), .ZN(
        n9011) );
  OAI22_X1 U3483 ( .A1(n17106), .A2(n11858), .B1(n17102), .B2(n16788), .ZN(
        n9012) );
  OAI22_X1 U3484 ( .A1(n17132), .A2(n15750), .B1(n17128), .B2(n16788), .ZN(
        n9014) );
  OAI22_X1 U3485 ( .A1(n17234), .A2(n15387), .B1(n17230), .B2(n16789), .ZN(
        n9023) );
  OAI22_X1 U3486 ( .A1(n17247), .A2(n12257), .B1(n17243), .B2(n16789), .ZN(
        n9024) );
  OAI22_X1 U3487 ( .A1(n17260), .A2(n14846), .B1(n17256), .B2(n16789), .ZN(
        n9025) );
  OAI22_X1 U3488 ( .A1(n17286), .A2(n14392), .B1(n17282), .B2(n16789), .ZN(
        n9027) );
  OAI22_X1 U3489 ( .A1(n17299), .A2(n14620), .B1(n17295), .B2(n16789), .ZN(
        n9028) );
  OAI22_X1 U3490 ( .A1(n17325), .A2(n15307), .B1(n17321), .B2(n16789), .ZN(
        n9030) );
  OAI22_X1 U3491 ( .A1(n17338), .A2(n11896), .B1(n17334), .B2(n16789), .ZN(
        n9031) );
  OAI22_X1 U3492 ( .A1(n17351), .A2(n15101), .B1(n17347), .B2(n16789), .ZN(
        n9032) );
  OAI22_X1 U3493 ( .A1(n17364), .A2(n15684), .B1(n17360), .B2(n16789), .ZN(
        n9033) );
  OAI22_X1 U3494 ( .A1(n17377), .A2(n14455), .B1(n17373), .B2(n16790), .ZN(
        n9034) );
  OAI22_X1 U3495 ( .A1(n17390), .A2(n14743), .B1(n17386), .B2(n16790), .ZN(
        n9035) );
  OAI22_X1 U3496 ( .A1(n17403), .A2(n14344), .B1(n17399), .B2(n16790), .ZN(
        n9036) );
  OAI22_X1 U3497 ( .A1(n17429), .A2(n15342), .B1(n17425), .B2(n16790), .ZN(
        n9038) );
  OAI22_X1 U3498 ( .A1(n17442), .A2(n14036), .B1(n17438), .B2(n16790), .ZN(
        n9039) );
  OAI22_X1 U3499 ( .A1(n17455), .A2(n14742), .B1(n17450), .B2(n16790), .ZN(
        n9040) );
  OAI22_X1 U3500 ( .A1(n17468), .A2(n15537), .B1(n17464), .B2(n16790), .ZN(
        n9041) );
  OAI22_X1 U3501 ( .A1(n17481), .A2(n15774), .B1(n17477), .B2(n16790), .ZN(
        n9042) );
  OAI22_X1 U3502 ( .A1(n17494), .A2(n14801), .B1(n17490), .B2(n16790), .ZN(
        n9043) );
  OAI22_X1 U3503 ( .A1(n17507), .A2(n15610), .B1(n17503), .B2(n16790), .ZN(
        n9044) );
  OAI22_X1 U3504 ( .A1(n17581), .A2(n14261), .B1(n17576), .B2(n16791), .ZN(
        n9049) );
  OAI22_X1 U3505 ( .A1(n18008), .A2(n12104), .B1(n18004), .B2(n16792), .ZN(
        n9062) );
  OAI22_X1 U3506 ( .A1(n18021), .A2(n14585), .B1(n18017), .B2(n16792), .ZN(
        n9063) );
  OAI22_X1 U3507 ( .A1(n16939), .A2(n14562), .B1(n16935), .B2(n16793), .ZN(
        n9070) );
  OAI22_X1 U3508 ( .A1(n17028), .A2(n12188), .B1(n17024), .B2(n16793), .ZN(
        n9078) );
  OAI22_X1 U3509 ( .A1(n17041), .A2(n15052), .B1(n17037), .B2(n16793), .ZN(
        n9079) );
  OAI22_X1 U3510 ( .A1(n17054), .A2(n14393), .B1(n17050), .B2(n16793), .ZN(
        n9080) );
  OAI22_X1 U3511 ( .A1(n17067), .A2(n15168), .B1(n17063), .B2(n16793), .ZN(
        n9081) );
  OAI22_X1 U3512 ( .A1(n17080), .A2(n15611), .B1(n17076), .B2(n16794), .ZN(
        n9082) );
  OAI22_X1 U3513 ( .A1(n17093), .A2(n15511), .B1(n17089), .B2(n16794), .ZN(
        n9083) );
  OAI22_X1 U3514 ( .A1(n17106), .A2(n11860), .B1(n17102), .B2(n16794), .ZN(
        n9084) );
  OAI22_X1 U3515 ( .A1(n17132), .A2(n15751), .B1(n17128), .B2(n16794), .ZN(
        n9086) );
  OAI22_X1 U3516 ( .A1(n17234), .A2(n15388), .B1(n17230), .B2(n16795), .ZN(
        n9095) );
  OAI22_X1 U3517 ( .A1(n17247), .A2(n12258), .B1(n17243), .B2(n16795), .ZN(
        n9096) );
  OAI22_X1 U3518 ( .A1(n17260), .A2(n14847), .B1(n17256), .B2(n16795), .ZN(
        n9097) );
  OAI22_X1 U3519 ( .A1(n17286), .A2(n14394), .B1(n17282), .B2(n16795), .ZN(
        n9099) );
  OAI22_X1 U3520 ( .A1(n17299), .A2(n14621), .B1(n17295), .B2(n16795), .ZN(
        n9100) );
  OAI22_X1 U3521 ( .A1(n17325), .A2(n15308), .B1(n17321), .B2(n16795), .ZN(
        n9102) );
  OAI22_X1 U3522 ( .A1(n17338), .A2(n11897), .B1(n17334), .B2(n16795), .ZN(
        n9103) );
  OAI22_X1 U3523 ( .A1(n17351), .A2(n15103), .B1(n17347), .B2(n16795), .ZN(
        n9104) );
  OAI22_X1 U3524 ( .A1(n17364), .A2(n15685), .B1(n17360), .B2(n16795), .ZN(
        n9105) );
  OAI22_X1 U3525 ( .A1(n17377), .A2(n14457), .B1(n17373), .B2(n16796), .ZN(
        n9106) );
  OAI22_X1 U3526 ( .A1(n17390), .A2(n14745), .B1(n17386), .B2(n16796), .ZN(
        n9107) );
  OAI22_X1 U3527 ( .A1(n17403), .A2(n14345), .B1(n17399), .B2(n16796), .ZN(
        n9108) );
  OAI22_X1 U3528 ( .A1(n17429), .A2(n15343), .B1(n17425), .B2(n16796), .ZN(
        n9110) );
  OAI22_X1 U3529 ( .A1(n17442), .A2(n14038), .B1(n17438), .B2(n16796), .ZN(
        n9111) );
  OAI22_X1 U3530 ( .A1(n17455), .A2(n14744), .B1(n17450), .B2(n16796), .ZN(
        n9112) );
  OAI22_X1 U3531 ( .A1(n17468), .A2(n15538), .B1(n17464), .B2(n16796), .ZN(
        n9113) );
  OAI22_X1 U3532 ( .A1(n17481), .A2(n15775), .B1(n17477), .B2(n16796), .ZN(
        n9114) );
  OAI22_X1 U3533 ( .A1(n17494), .A2(n14803), .B1(n17490), .B2(n16796), .ZN(
        n9115) );
  OAI22_X1 U3534 ( .A1(n17507), .A2(n15612), .B1(n17503), .B2(n16796), .ZN(
        n9116) );
  OAI22_X1 U3535 ( .A1(n17581), .A2(n14264), .B1(n17576), .B2(n16797), .ZN(
        n9121) );
  OAI22_X1 U3536 ( .A1(n18008), .A2(n12105), .B1(n18004), .B2(n16798), .ZN(
        n9134) );
  OAI22_X1 U3537 ( .A1(n18021), .A2(n14586), .B1(n18017), .B2(n16798), .ZN(
        n9135) );
  OAI22_X1 U3538 ( .A1(n16939), .A2(n14563), .B1(n16935), .B2(n16799), .ZN(
        n9142) );
  OAI22_X1 U3539 ( .A1(n17028), .A2(n12189), .B1(n17024), .B2(n16799), .ZN(
        n9150) );
  OAI22_X1 U3540 ( .A1(n17041), .A2(n15053), .B1(n17037), .B2(n16799), .ZN(
        n9151) );
  OAI22_X1 U3541 ( .A1(n17054), .A2(n14395), .B1(n17050), .B2(n16799), .ZN(
        n9152) );
  OAI22_X1 U3542 ( .A1(n17080), .A2(n15613), .B1(n17076), .B2(n16800), .ZN(
        n9154) );
  OAI22_X1 U3543 ( .A1(n17132), .A2(n15752), .B1(n17128), .B2(n16800), .ZN(
        n9158) );
  OAI22_X1 U3544 ( .A1(n17234), .A2(n15389), .B1(n17230), .B2(n16801), .ZN(
        n9167) );
  OAI22_X1 U3545 ( .A1(n17247), .A2(n12301), .B1(n17243), .B2(n16801), .ZN(
        n9168) );
  OAI22_X1 U3546 ( .A1(n17325), .A2(n15309), .B1(n17321), .B2(n16801), .ZN(
        n9174) );
  OAI22_X1 U3547 ( .A1(n17338), .A2(n11898), .B1(n17334), .B2(n16801), .ZN(
        n9175) );
  OAI22_X1 U3548 ( .A1(n17351), .A2(n15105), .B1(n17347), .B2(n16801), .ZN(
        n9176) );
  OAI22_X1 U3549 ( .A1(n17377), .A2(n14459), .B1(n17373), .B2(n16802), .ZN(
        n9178) );
  OAI22_X1 U3550 ( .A1(n17428), .A2(n15344), .B1(n17425), .B2(n16802), .ZN(
        n9182) );
  OAI22_X1 U3551 ( .A1(n17441), .A2(n14040), .B1(n17438), .B2(n16802), .ZN(
        n9183) );
  OAI22_X1 U3552 ( .A1(n17454), .A2(n14746), .B1(n17450), .B2(n16802), .ZN(
        n9184) );
  OAI22_X1 U3553 ( .A1(n17480), .A2(n15776), .B1(n17477), .B2(n16802), .ZN(
        n9186) );
  OAI22_X1 U3554 ( .A1(n18008), .A2(n12148), .B1(n18004), .B2(n16804), .ZN(
        n9206) );
  OAI22_X1 U3555 ( .A1(n16939), .A2(n14564), .B1(n16935), .B2(n16805), .ZN(
        n9214) );
  OAI22_X1 U3556 ( .A1(n17027), .A2(n12190), .B1(n17024), .B2(n16805), .ZN(
        n9222) );
  OAI22_X1 U3557 ( .A1(n17132), .A2(n15753), .B1(n17128), .B2(n16806), .ZN(
        n9230) );
  OAI22_X1 U3558 ( .A1(n17324), .A2(n15310), .B1(n17321), .B2(n16807), .ZN(
        n9246) );
  OAI22_X1 U3559 ( .A1(n17428), .A2(n15345), .B1(n17425), .B2(n16808), .ZN(
        n9254) );
  OAI22_X1 U3560 ( .A1(n17582), .A2(n14268), .B1(n17576), .B2(n16821), .ZN(
        n9409) );
  OAI22_X1 U3561 ( .A1(n18009), .A2(n12152), .B1(n18004), .B2(n16822), .ZN(
        n9422) );
  OAI22_X1 U3562 ( .A1(n18022), .A2(n14590), .B1(n18017), .B2(n16822), .ZN(
        n9423) );
  OAI22_X1 U3563 ( .A1(n16940), .A2(n14545), .B1(n16935), .B2(n17514), .ZN(
        n9934) );
  OAI22_X1 U3564 ( .A1(n17029), .A2(n12170), .B1(n17024), .B2(n17514), .ZN(
        n9942) );
  OAI22_X1 U3565 ( .A1(n17042), .A2(n15054), .B1(n17037), .B2(n17514), .ZN(
        n9943) );
  OAI22_X1 U3566 ( .A1(n17055), .A2(n14396), .B1(n17050), .B2(n17514), .ZN(
        n9944) );
  OAI22_X1 U3567 ( .A1(n17068), .A2(n15169), .B1(n17063), .B2(n17514), .ZN(
        n9945) );
  OAI22_X1 U3568 ( .A1(n17081), .A2(n15614), .B1(n17076), .B2(n17515), .ZN(
        n9946) );
  OAI22_X1 U3569 ( .A1(n17094), .A2(n15494), .B1(n17089), .B2(n17515), .ZN(
        n9947) );
  OAI22_X1 U3570 ( .A1(n17107), .A2(n11861), .B1(n17102), .B2(n17515), .ZN(
        n9948) );
  OAI22_X1 U3571 ( .A1(n17133), .A2(n15734), .B1(n17128), .B2(n17515), .ZN(
        n9950) );
  OAI22_X1 U3572 ( .A1(n17235), .A2(n15390), .B1(n17230), .B2(n17516), .ZN(
        n9959) );
  OAI22_X1 U3573 ( .A1(n17248), .A2(n12204), .B1(n17243), .B2(n17516), .ZN(
        n9960) );
  OAI22_X1 U3574 ( .A1(n17261), .A2(n14830), .B1(n17256), .B2(n17516), .ZN(
        n9961) );
  OAI22_X1 U3575 ( .A1(n17287), .A2(n14397), .B1(n17282), .B2(n17516), .ZN(
        n9963) );
  OAI22_X1 U3576 ( .A1(n17300), .A2(n14604), .B1(n17295), .B2(n17516), .ZN(
        n9964) );
  OAI22_X1 U3577 ( .A1(n17326), .A2(n15291), .B1(n17321), .B2(n17516), .ZN(
        n9966) );
  OAI22_X1 U3578 ( .A1(n17339), .A2(n11880), .B1(n17334), .B2(n17516), .ZN(
        n9967) );
  OAI22_X1 U3579 ( .A1(n17352), .A2(n15070), .B1(n17347), .B2(n17516), .ZN(
        n9968) );
  OAI22_X1 U3580 ( .A1(n17365), .A2(n15668), .B1(n17360), .B2(n17516), .ZN(
        n9969) );
  OAI22_X1 U3581 ( .A1(n17378), .A2(n14424), .B1(n17373), .B2(n17517), .ZN(
        n9970) );
  OAI22_X1 U3582 ( .A1(n17391), .A2(n14710), .B1(n17386), .B2(n17517), .ZN(
        n9971) );
  OAI22_X1 U3583 ( .A1(n17404), .A2(n14357), .B1(n17399), .B2(n17517), .ZN(
        n9972) );
  OAI22_X1 U3584 ( .A1(n17430), .A2(n15325), .B1(n17425), .B2(n17517), .ZN(
        n9974) );
  OAI22_X1 U3585 ( .A1(n17443), .A2(n12347), .B1(n17438), .B2(n17517), .ZN(
        n9975) );
  OAI22_X1 U3586 ( .A1(n17456), .A2(n14709), .B1(n17450), .B2(n17517), .ZN(
        n9976) );
  OAI22_X1 U3587 ( .A1(n17469), .A2(n15457), .B1(n17464), .B2(n17517), .ZN(
        n9977) );
  OAI22_X1 U3588 ( .A1(n17482), .A2(n15735), .B1(n17477), .B2(n17517), .ZN(
        n9978) );
  OAI22_X1 U3589 ( .A1(n17495), .A2(n14769), .B1(n17490), .B2(n17517), .ZN(
        n9979) );
  OAI22_X1 U3590 ( .A1(n17508), .A2(n15615), .B1(n17503), .B2(n17517), .ZN(
        n9980) );
  BUF_X1 U3591 ( .A(n4223), .Z(n17666) );
  BUF_X1 U3592 ( .A(n4202), .Z(n17690) );
  NAND2_X1 U3593 ( .A1(N273), .A2(n14262), .ZN(n14064) );
  OAI22_X1 U3594 ( .A1(n16700), .A2(n14980), .B1(n16692), .B2(n16456), .ZN(
        n7981) );
  OAI22_X1 U3595 ( .A1(n16695), .A2(n14981), .B1(n16691), .B2(n16815), .ZN(
        n8089) );
  OAI22_X1 U3596 ( .A1(n16695), .A2(n14982), .B1(n16692), .B2(n16821), .ZN(
        n8091) );
  OAI22_X1 U3597 ( .A1(n16694), .A2(n14983), .B1(n16692), .B2(n16833), .ZN(
        n8095) );
  OAI22_X1 U3598 ( .A1(n16694), .A2(n14984), .B1(n16691), .B2(n16839), .ZN(
        n8097) );
  OAI22_X1 U3599 ( .A1(n16694), .A2(n14985), .B1(n16692), .B2(n16845), .ZN(
        n8099) );
  OAI22_X1 U3600 ( .A1(n16693), .A2(n14986), .B1(n16692), .B2(n16851), .ZN(
        n8101) );
  OAI22_X1 U3601 ( .A1(n16695), .A2(n14987), .B1(n16691), .B2(n16857), .ZN(
        n8103) );
  OAI22_X1 U3602 ( .A1(n16694), .A2(n14988), .B1(n16692), .B2(n17512), .ZN(
        n8105) );
  OAI22_X1 U3603 ( .A1(n18008), .A2(n12150), .B1(n18003), .B2(n16810), .ZN(
        n9278) );
  OAI22_X1 U3604 ( .A1(n16938), .A2(n14565), .B1(n16934), .B2(n16811), .ZN(
        n9286) );
  OAI22_X1 U3605 ( .A1(n17027), .A2(n12191), .B1(n17023), .B2(n16811), .ZN(
        n9294) );
  OAI22_X1 U3606 ( .A1(n17131), .A2(n15754), .B1(n17127), .B2(n16812), .ZN(
        n9302) );
  OAI22_X1 U3607 ( .A1(n17324), .A2(n15311), .B1(n17320), .B2(n16813), .ZN(
        n9318) );
  OAI22_X1 U3608 ( .A1(n17428), .A2(n15346), .B1(n17424), .B2(n16814), .ZN(
        n9326) );
  OAI22_X1 U3609 ( .A1(n18007), .A2(n12151), .B1(n18003), .B2(n16816), .ZN(
        n9350) );
  OAI22_X1 U3610 ( .A1(n16938), .A2(n14566), .B1(n16934), .B2(n16817), .ZN(
        n9358) );
  OAI22_X1 U3611 ( .A1(n17027), .A2(n12192), .B1(n17023), .B2(n16817), .ZN(
        n9366) );
  OAI22_X1 U3612 ( .A1(n17131), .A2(n15755), .B1(n17127), .B2(n16818), .ZN(
        n9374) );
  OAI22_X1 U3613 ( .A1(n17324), .A2(n15312), .B1(n17320), .B2(n16819), .ZN(
        n9390) );
  OAI22_X1 U3614 ( .A1(n17428), .A2(n15347), .B1(n17424), .B2(n16820), .ZN(
        n9398) );
  OAI22_X1 U3615 ( .A1(n16938), .A2(n14567), .B1(n16934), .B2(n16823), .ZN(
        n9430) );
  OAI22_X1 U3616 ( .A1(n17027), .A2(n12193), .B1(n17023), .B2(n16823), .ZN(
        n9438) );
  OAI22_X1 U3617 ( .A1(n17131), .A2(n15756), .B1(n17127), .B2(n16824), .ZN(
        n9446) );
  OAI22_X1 U3618 ( .A1(n17323), .A2(n15313), .B1(n17320), .B2(n16825), .ZN(
        n9462) );
  OAI22_X1 U3619 ( .A1(n17427), .A2(n15348), .B1(n17424), .B2(n16826), .ZN(
        n9470) );
  OAI22_X1 U3620 ( .A1(n18007), .A2(n12153), .B1(n18003), .B2(n16828), .ZN(
        n9494) );
  OAI22_X1 U3621 ( .A1(n16937), .A2(n14568), .B1(n16934), .B2(n16829), .ZN(
        n9502) );
  OAI22_X1 U3622 ( .A1(n17026), .A2(n12164), .B1(n17023), .B2(n16829), .ZN(
        n9510) );
  OAI22_X1 U3623 ( .A1(n17130), .A2(n15722), .B1(n17127), .B2(n16830), .ZN(
        n9518) );
  OAI22_X1 U3624 ( .A1(n17323), .A2(n15285), .B1(n17320), .B2(n16831), .ZN(
        n9534) );
  OAI22_X1 U3625 ( .A1(n17427), .A2(n15319), .B1(n17424), .B2(n16832), .ZN(
        n9542) );
  OAI22_X1 U3626 ( .A1(n18007), .A2(n12154), .B1(n18003), .B2(n16834), .ZN(
        n9566) );
  OAI22_X1 U3627 ( .A1(n16938), .A2(n14540), .B1(n16934), .B2(n16835), .ZN(
        n9574) );
  OAI22_X1 U3628 ( .A1(n17026), .A2(n12165), .B1(n17023), .B2(n16835), .ZN(
        n9582) );
  OAI22_X1 U3629 ( .A1(n17131), .A2(n15724), .B1(n17127), .B2(n16836), .ZN(
        n9590) );
  OAI22_X1 U3630 ( .A1(n17324), .A2(n15286), .B1(n17320), .B2(n16837), .ZN(
        n9606) );
  OAI22_X1 U3631 ( .A1(n17427), .A2(n15320), .B1(n17424), .B2(n16838), .ZN(
        n9614) );
  OAI22_X1 U3632 ( .A1(n18007), .A2(n12155), .B1(n18003), .B2(n16840), .ZN(
        n9638) );
  OAI22_X1 U3633 ( .A1(n16937), .A2(n14541), .B1(n16934), .B2(n16841), .ZN(
        n9646) );
  OAI22_X1 U3634 ( .A1(n17026), .A2(n12166), .B1(n17023), .B2(n16841), .ZN(
        n9654) );
  OAI22_X1 U3635 ( .A1(n17130), .A2(n15726), .B1(n17127), .B2(n16842), .ZN(
        n9662) );
  OAI22_X1 U3636 ( .A1(n17323), .A2(n15287), .B1(n17320), .B2(n16843), .ZN(
        n9678) );
  OAI22_X1 U3637 ( .A1(n17427), .A2(n15321), .B1(n17424), .B2(n16844), .ZN(
        n9686) );
  OAI22_X1 U3638 ( .A1(n18006), .A2(n12156), .B1(n18003), .B2(n16846), .ZN(
        n9710) );
  OAI22_X1 U3639 ( .A1(n16937), .A2(n14542), .B1(n16934), .B2(n16847), .ZN(
        n9718) );
  OAI22_X1 U3640 ( .A1(n17026), .A2(n12167), .B1(n17023), .B2(n16847), .ZN(
        n9726) );
  OAI22_X1 U3641 ( .A1(n17130), .A2(n15728), .B1(n17127), .B2(n16848), .ZN(
        n9734) );
  OAI22_X1 U3642 ( .A1(n17323), .A2(n15288), .B1(n17320), .B2(n16849), .ZN(
        n9750) );
  OAI22_X1 U3643 ( .A1(n17426), .A2(n15322), .B1(n17424), .B2(n16850), .ZN(
        n9758) );
  OAI22_X1 U3644 ( .A1(n18006), .A2(n12157), .B1(n18003), .B2(n16852), .ZN(
        n9782) );
  OAI22_X1 U3645 ( .A1(n16937), .A2(n14543), .B1(n16934), .B2(n16853), .ZN(
        n9790) );
  OAI22_X1 U3646 ( .A1(n17025), .A2(n12168), .B1(n17023), .B2(n16853), .ZN(
        n9798) );
  OAI22_X1 U3647 ( .A1(n17130), .A2(n15730), .B1(n17127), .B2(n16854), .ZN(
        n9806) );
  OAI22_X1 U3648 ( .A1(n17322), .A2(n15289), .B1(n17320), .B2(n16855), .ZN(
        n9822) );
  OAI22_X1 U3649 ( .A1(n17426), .A2(n15323), .B1(n17424), .B2(n16856), .ZN(
        n9830) );
  OAI22_X1 U3650 ( .A1(n18006), .A2(n12158), .B1(n18003), .B2(n16858), .ZN(
        n9854) );
  OAI22_X1 U3651 ( .A1(n16936), .A2(n14544), .B1(n16934), .B2(n16859), .ZN(
        n9862) );
  OAI22_X1 U3652 ( .A1(n17025), .A2(n12169), .B1(n17023), .B2(n16859), .ZN(
        n9870) );
  OAI22_X1 U3653 ( .A1(n17129), .A2(n15732), .B1(n17127), .B2(n16860), .ZN(
        n9878) );
  OAI22_X1 U3654 ( .A1(n17322), .A2(n15290), .B1(n17320), .B2(n16861), .ZN(
        n9894) );
  OAI22_X1 U3655 ( .A1(n17426), .A2(n15324), .B1(n17424), .B2(n16862), .ZN(
        n9902) );
  OAI22_X1 U3656 ( .A1(n18006), .A2(n12159), .B1(n18003), .B2(n17513), .ZN(
        n9926) );
  OAI22_X1 U3657 ( .A1(n17581), .A2(n14269), .B1(n17576), .B2(n16803), .ZN(
        n9193) );
  OAI22_X1 U3658 ( .A1(n18021), .A2(n14587), .B1(n18016), .B2(n16804), .ZN(
        n9207) );
  OAI22_X1 U3659 ( .A1(n17040), .A2(n15055), .B1(n17036), .B2(n16805), .ZN(
        n9223) );
  OAI22_X1 U3660 ( .A1(n17053), .A2(n14398), .B1(n17049), .B2(n16805), .ZN(
        n9224) );
  OAI22_X1 U3661 ( .A1(n17079), .A2(n15616), .B1(n17075), .B2(n16806), .ZN(
        n9226) );
  OAI22_X1 U3662 ( .A1(n17233), .A2(n15391), .B1(n17229), .B2(n16807), .ZN(
        n9239) );
  OAI22_X1 U3663 ( .A1(n17246), .A2(n12303), .B1(n17242), .B2(n16807), .ZN(
        n9240) );
  OAI22_X1 U3664 ( .A1(n17337), .A2(n11899), .B1(n17333), .B2(n16807), .ZN(
        n9247) );
  OAI22_X1 U3665 ( .A1(n17350), .A2(n15107), .B1(n17346), .B2(n16807), .ZN(
        n9248) );
  OAI22_X1 U3666 ( .A1(n17376), .A2(n14461), .B1(n17372), .B2(n16808), .ZN(
        n9250) );
  OAI22_X1 U3667 ( .A1(n17441), .A2(n14042), .B1(n17437), .B2(n16808), .ZN(
        n9255) );
  OAI22_X1 U3668 ( .A1(n17454), .A2(n14748), .B1(n17450), .B2(n16808), .ZN(
        n9256) );
  OAI22_X1 U3669 ( .A1(n17480), .A2(n15777), .B1(n17476), .B2(n16808), .ZN(
        n9258) );
  OAI22_X1 U3670 ( .A1(n17580), .A2(n14270), .B1(n17576), .B2(n16809), .ZN(
        n9265) );
  OAI22_X1 U3671 ( .A1(n18021), .A2(n14588), .B1(n18016), .B2(n16810), .ZN(
        n9279) );
  OAI22_X1 U3672 ( .A1(n17040), .A2(n15056), .B1(n17036), .B2(n16811), .ZN(
        n9295) );
  OAI22_X1 U3673 ( .A1(n17053), .A2(n14399), .B1(n17049), .B2(n16811), .ZN(
        n9296) );
  OAI22_X1 U3674 ( .A1(n17079), .A2(n15617), .B1(n17075), .B2(n16812), .ZN(
        n9298) );
  OAI22_X1 U3675 ( .A1(n17233), .A2(n15392), .B1(n17229), .B2(n16813), .ZN(
        n9311) );
  OAI22_X1 U3676 ( .A1(n17246), .A2(n12304), .B1(n17242), .B2(n16813), .ZN(
        n9312) );
  OAI22_X1 U3677 ( .A1(n17337), .A2(n11900), .B1(n17333), .B2(n16813), .ZN(
        n9319) );
  OAI22_X1 U3678 ( .A1(n17350), .A2(n15109), .B1(n17346), .B2(n16813), .ZN(
        n9320) );
  OAI22_X1 U3679 ( .A1(n17376), .A2(n14463), .B1(n17372), .B2(n16814), .ZN(
        n9322) );
  OAI22_X1 U3680 ( .A1(n17441), .A2(n14044), .B1(n17437), .B2(n16814), .ZN(
        n9327) );
  OAI22_X1 U3681 ( .A1(n17454), .A2(n14750), .B1(n17450), .B2(n16814), .ZN(
        n9328) );
  OAI22_X1 U3682 ( .A1(n17480), .A2(n15778), .B1(n17476), .B2(n16814), .ZN(
        n9330) );
  OAI22_X1 U3683 ( .A1(n17580), .A2(n14271), .B1(n17577), .B2(n16815), .ZN(
        n9337) );
  OAI22_X1 U3684 ( .A1(n18020), .A2(n14589), .B1(n18016), .B2(n16816), .ZN(
        n9351) );
  OAI22_X1 U3685 ( .A1(n17040), .A2(n15057), .B1(n17036), .B2(n16817), .ZN(
        n9367) );
  OAI22_X1 U3686 ( .A1(n17053), .A2(n14400), .B1(n17049), .B2(n16817), .ZN(
        n9368) );
  OAI22_X1 U3687 ( .A1(n17079), .A2(n15618), .B1(n17075), .B2(n16818), .ZN(
        n9370) );
  OAI22_X1 U3688 ( .A1(n17233), .A2(n15393), .B1(n17229), .B2(n16819), .ZN(
        n9383) );
  OAI22_X1 U3689 ( .A1(n17246), .A2(n12305), .B1(n17242), .B2(n16819), .ZN(
        n9384) );
  OAI22_X1 U3690 ( .A1(n17337), .A2(n11901), .B1(n17333), .B2(n16819), .ZN(
        n9391) );
  OAI22_X1 U3691 ( .A1(n17350), .A2(n15111), .B1(n17346), .B2(n16819), .ZN(
        n9392) );
  OAI22_X1 U3692 ( .A1(n17376), .A2(n14465), .B1(n17372), .B2(n16820), .ZN(
        n9394) );
  OAI22_X1 U3693 ( .A1(n17441), .A2(n14046), .B1(n17437), .B2(n16820), .ZN(
        n9399) );
  OAI22_X1 U3694 ( .A1(n17454), .A2(n14752), .B1(n17451), .B2(n16820), .ZN(
        n9400) );
  OAI22_X1 U3695 ( .A1(n17480), .A2(n15779), .B1(n17476), .B2(n16820), .ZN(
        n9402) );
  OAI22_X1 U3696 ( .A1(n17040), .A2(n15058), .B1(n17036), .B2(n16823), .ZN(
        n9439) );
  OAI22_X1 U3697 ( .A1(n17053), .A2(n14401), .B1(n17049), .B2(n16823), .ZN(
        n9440) );
  OAI22_X1 U3698 ( .A1(n17079), .A2(n15619), .B1(n17075), .B2(n16824), .ZN(
        n9442) );
  OAI22_X1 U3699 ( .A1(n17233), .A2(n15394), .B1(n17229), .B2(n16825), .ZN(
        n9455) );
  OAI22_X1 U3700 ( .A1(n17246), .A2(n12306), .B1(n17242), .B2(n16825), .ZN(
        n9456) );
  OAI22_X1 U3701 ( .A1(n17336), .A2(n11902), .B1(n17333), .B2(n16825), .ZN(
        n9463) );
  OAI22_X1 U3702 ( .A1(n17349), .A2(n15113), .B1(n17346), .B2(n16825), .ZN(
        n9464) );
  OAI22_X1 U3703 ( .A1(n17375), .A2(n14467), .B1(n17372), .B2(n16826), .ZN(
        n9466) );
  OAI22_X1 U3704 ( .A1(n17440), .A2(n14048), .B1(n17437), .B2(n16826), .ZN(
        n9471) );
  OAI22_X1 U3705 ( .A1(n17453), .A2(n14754), .B1(n17451), .B2(n16826), .ZN(
        n9472) );
  OAI22_X1 U3706 ( .A1(n17479), .A2(n15780), .B1(n17476), .B2(n16826), .ZN(
        n9474) );
  OAI22_X1 U3707 ( .A1(n17580), .A2(n14272), .B1(n17577), .B2(n16827), .ZN(
        n9481) );
  OAI22_X1 U3708 ( .A1(n18020), .A2(n14591), .B1(n18016), .B2(n16828), .ZN(
        n9495) );
  OAI22_X1 U3709 ( .A1(n17039), .A2(n15059), .B1(n17036), .B2(n16829), .ZN(
        n9511) );
  OAI22_X1 U3710 ( .A1(n17052), .A2(n14402), .B1(n17049), .B2(n16829), .ZN(
        n9512) );
  OAI22_X1 U3711 ( .A1(n17078), .A2(n15620), .B1(n17075), .B2(n16830), .ZN(
        n9514) );
  OAI22_X1 U3712 ( .A1(n17232), .A2(n15395), .B1(n17229), .B2(n16831), .ZN(
        n9527) );
  OAI22_X1 U3713 ( .A1(n17245), .A2(n12198), .B1(n17242), .B2(n16831), .ZN(
        n9528) );
  OAI22_X1 U3714 ( .A1(n17336), .A2(n11874), .B1(n17333), .B2(n16831), .ZN(
        n9535) );
  OAI22_X1 U3715 ( .A1(n17349), .A2(n15115), .B1(n17346), .B2(n16831), .ZN(
        n9536) );
  OAI22_X1 U3716 ( .A1(n17375), .A2(n14469), .B1(n17372), .B2(n16832), .ZN(
        n9538) );
  OAI22_X1 U3717 ( .A1(n17440), .A2(n14050), .B1(n17437), .B2(n16832), .ZN(
        n9543) );
  OAI22_X1 U3718 ( .A1(n17453), .A2(n14817), .B1(n17451), .B2(n16832), .ZN(
        n9544) );
  OAI22_X1 U3719 ( .A1(n17479), .A2(n15723), .B1(n17476), .B2(n16832), .ZN(
        n9546) );
  OAI22_X1 U3720 ( .A1(n17579), .A2(n14273), .B1(n17577), .B2(n16833), .ZN(
        n9553) );
  OAI22_X1 U3721 ( .A1(n18020), .A2(n14592), .B1(n18016), .B2(n16834), .ZN(
        n9567) );
  OAI22_X1 U3722 ( .A1(n17039), .A2(n15060), .B1(n17036), .B2(n16835), .ZN(
        n9583) );
  OAI22_X1 U3723 ( .A1(n17052), .A2(n14403), .B1(n17049), .B2(n16835), .ZN(
        n9584) );
  OAI22_X1 U3724 ( .A1(n17078), .A2(n15621), .B1(n17075), .B2(n16836), .ZN(
        n9586) );
  OAI22_X1 U3725 ( .A1(n17232), .A2(n15396), .B1(n17229), .B2(n16837), .ZN(
        n9599) );
  OAI22_X1 U3726 ( .A1(n17245), .A2(n12199), .B1(n17242), .B2(n16837), .ZN(
        n9600) );
  OAI22_X1 U3727 ( .A1(n17337), .A2(n11875), .B1(n17333), .B2(n16837), .ZN(
        n9607) );
  OAI22_X1 U3728 ( .A1(n17350), .A2(n15065), .B1(n17346), .B2(n16837), .ZN(
        n9608) );
  OAI22_X1 U3729 ( .A1(n17376), .A2(n14419), .B1(n17372), .B2(n16838), .ZN(
        n9610) );
  OAI22_X1 U3730 ( .A1(n17440), .A2(n12342), .B1(n17437), .B2(n16838), .ZN(
        n9615) );
  OAI22_X1 U3731 ( .A1(n17453), .A2(n14818), .B1(n17451), .B2(n16838), .ZN(
        n9616) );
  OAI22_X1 U3732 ( .A1(n17479), .A2(n15725), .B1(n17476), .B2(n16838), .ZN(
        n9618) );
  OAI22_X1 U3733 ( .A1(n17580), .A2(n14274), .B1(n17577), .B2(n16839), .ZN(
        n9625) );
  OAI22_X1 U3734 ( .A1(n18020), .A2(n14593), .B1(n18016), .B2(n16840), .ZN(
        n9639) );
  OAI22_X1 U3735 ( .A1(n17039), .A2(n15061), .B1(n17036), .B2(n16841), .ZN(
        n9655) );
  OAI22_X1 U3736 ( .A1(n17052), .A2(n14404), .B1(n17049), .B2(n16841), .ZN(
        n9656) );
  OAI22_X1 U3737 ( .A1(n17078), .A2(n15622), .B1(n17075), .B2(n16842), .ZN(
        n9658) );
  OAI22_X1 U3738 ( .A1(n17232), .A2(n15397), .B1(n17229), .B2(n16843), .ZN(
        n9671) );
  OAI22_X1 U3739 ( .A1(n17245), .A2(n12200), .B1(n17242), .B2(n16843), .ZN(
        n9672) );
  OAI22_X1 U3740 ( .A1(n17336), .A2(n11876), .B1(n17333), .B2(n16843), .ZN(
        n9679) );
  OAI22_X1 U3741 ( .A1(n17349), .A2(n15066), .B1(n17346), .B2(n16843), .ZN(
        n9680) );
  OAI22_X1 U3742 ( .A1(n17375), .A2(n14420), .B1(n17372), .B2(n16844), .ZN(
        n9682) );
  OAI22_X1 U3743 ( .A1(n17440), .A2(n12343), .B1(n17437), .B2(n16844), .ZN(
        n9687) );
  OAI22_X1 U3744 ( .A1(n17453), .A2(n14819), .B1(n17451), .B2(n16844), .ZN(
        n9688) );
  OAI22_X1 U3745 ( .A1(n17479), .A2(n15727), .B1(n17476), .B2(n16844), .ZN(
        n9690) );
  OAI22_X1 U3746 ( .A1(n17579), .A2(n14275), .B1(n17577), .B2(n16845), .ZN(
        n9697) );
  OAI22_X1 U3747 ( .A1(n18019), .A2(n14594), .B1(n18016), .B2(n16846), .ZN(
        n9711) );
  OAI22_X1 U3748 ( .A1(n17039), .A2(n15062), .B1(n17036), .B2(n16847), .ZN(
        n9727) );
  OAI22_X1 U3749 ( .A1(n17052), .A2(n14405), .B1(n17049), .B2(n16847), .ZN(
        n9728) );
  OAI22_X1 U3750 ( .A1(n17078), .A2(n15623), .B1(n17075), .B2(n16848), .ZN(
        n9730) );
  OAI22_X1 U3751 ( .A1(n17232), .A2(n15398), .B1(n17229), .B2(n16849), .ZN(
        n9743) );
  OAI22_X1 U3752 ( .A1(n17245), .A2(n12201), .B1(n17242), .B2(n16849), .ZN(
        n9744) );
  OAI22_X1 U3753 ( .A1(n17336), .A2(n11877), .B1(n17333), .B2(n16849), .ZN(
        n9751) );
  OAI22_X1 U3754 ( .A1(n17349), .A2(n15067), .B1(n17346), .B2(n16849), .ZN(
        n9752) );
  OAI22_X1 U3755 ( .A1(n17375), .A2(n14421), .B1(n17372), .B2(n16850), .ZN(
        n9754) );
  OAI22_X1 U3756 ( .A1(n17439), .A2(n12344), .B1(n17437), .B2(n16850), .ZN(
        n9759) );
  OAI22_X1 U3757 ( .A1(n17452), .A2(n14703), .B1(n17451), .B2(n16850), .ZN(
        n9760) );
  OAI22_X1 U3758 ( .A1(n17478), .A2(n15729), .B1(n17476), .B2(n16850), .ZN(
        n9762) );
  OAI22_X1 U3759 ( .A1(n17579), .A2(n14276), .B1(n17577), .B2(n16851), .ZN(
        n9769) );
  OAI22_X1 U3760 ( .A1(n18019), .A2(n14595), .B1(n18016), .B2(n16852), .ZN(
        n9783) );
  OAI22_X1 U3761 ( .A1(n17038), .A2(n15063), .B1(n17036), .B2(n16853), .ZN(
        n9799) );
  OAI22_X1 U3762 ( .A1(n17051), .A2(n14406), .B1(n17049), .B2(n16853), .ZN(
        n9800) );
  OAI22_X1 U3763 ( .A1(n17077), .A2(n15624), .B1(n17075), .B2(n16854), .ZN(
        n9802) );
  OAI22_X1 U3764 ( .A1(n17231), .A2(n15399), .B1(n17229), .B2(n16855), .ZN(
        n9815) );
  OAI22_X1 U3765 ( .A1(n17244), .A2(n12202), .B1(n17242), .B2(n16855), .ZN(
        n9816) );
  OAI22_X1 U3766 ( .A1(n17335), .A2(n11878), .B1(n17333), .B2(n16855), .ZN(
        n9823) );
  OAI22_X1 U3767 ( .A1(n17348), .A2(n15068), .B1(n17346), .B2(n16855), .ZN(
        n9824) );
  OAI22_X1 U3768 ( .A1(n17374), .A2(n14422), .B1(n17372), .B2(n16856), .ZN(
        n9826) );
  OAI22_X1 U3769 ( .A1(n17439), .A2(n12345), .B1(n17437), .B2(n16856), .ZN(
        n9831) );
  OAI22_X1 U3770 ( .A1(n17452), .A2(n14705), .B1(n17450), .B2(n16856), .ZN(
        n9832) );
  OAI22_X1 U3771 ( .A1(n17478), .A2(n15731), .B1(n17476), .B2(n16856), .ZN(
        n9834) );
  OAI22_X1 U3772 ( .A1(n17579), .A2(n14277), .B1(n17576), .B2(n16857), .ZN(
        n9841) );
  OAI22_X1 U3773 ( .A1(n18019), .A2(n14596), .B1(n18016), .B2(n16858), .ZN(
        n9855) );
  OAI22_X1 U3774 ( .A1(n17038), .A2(n15064), .B1(n17036), .B2(n16859), .ZN(
        n9871) );
  OAI22_X1 U3775 ( .A1(n17051), .A2(n14407), .B1(n17049), .B2(n16859), .ZN(
        n9872) );
  OAI22_X1 U3776 ( .A1(n17077), .A2(n15625), .B1(n17075), .B2(n16860), .ZN(
        n9874) );
  OAI22_X1 U3777 ( .A1(n17231), .A2(n15400), .B1(n17229), .B2(n16861), .ZN(
        n9887) );
  OAI22_X1 U3778 ( .A1(n17244), .A2(n12203), .B1(n17242), .B2(n16861), .ZN(
        n9888) );
  OAI22_X1 U3779 ( .A1(n17335), .A2(n11879), .B1(n17333), .B2(n16861), .ZN(
        n9895) );
  OAI22_X1 U3780 ( .A1(n17348), .A2(n15069), .B1(n17346), .B2(n16861), .ZN(
        n9896) );
  OAI22_X1 U3781 ( .A1(n17374), .A2(n14423), .B1(n17372), .B2(n16862), .ZN(
        n9898) );
  OAI22_X1 U3782 ( .A1(n17439), .A2(n12346), .B1(n17437), .B2(n16862), .ZN(
        n9903) );
  OAI22_X1 U3783 ( .A1(n17452), .A2(n14707), .B1(n17451), .B2(n16862), .ZN(
        n9904) );
  OAI22_X1 U3784 ( .A1(n17478), .A2(n15733), .B1(n17476), .B2(n16862), .ZN(
        n9906) );
  OAI22_X1 U3785 ( .A1(n17578), .A2(n14278), .B1(n17577), .B2(n17512), .ZN(
        n9913) );
  OAI22_X1 U3786 ( .A1(n18019), .A2(n14597), .B1(n18016), .B2(n17513), .ZN(
        n9927) );
  OAI22_X1 U3787 ( .A1(n17067), .A2(n15170), .B1(n17062), .B2(n16799), .ZN(
        n9153) );
  OAI22_X1 U3788 ( .A1(n17093), .A2(n15512), .B1(n17088), .B2(n16800), .ZN(
        n9155) );
  OAI22_X1 U3789 ( .A1(n17106), .A2(n11862), .B1(n17101), .B2(n16800), .ZN(
        n9156) );
  OAI22_X1 U3790 ( .A1(n17260), .A2(n14848), .B1(n17255), .B2(n16801), .ZN(
        n9169) );
  OAI22_X1 U3791 ( .A1(n17286), .A2(n14408), .B1(n17281), .B2(n16801), .ZN(
        n9171) );
  OAI22_X1 U3792 ( .A1(n17299), .A2(n14622), .B1(n17294), .B2(n16801), .ZN(
        n9172) );
  OAI22_X1 U3793 ( .A1(n17364), .A2(n15686), .B1(n17359), .B2(n16801), .ZN(
        n9177) );
  OAI22_X1 U3794 ( .A1(n17390), .A2(n14747), .B1(n17385), .B2(n16802), .ZN(
        n9179) );
  OAI22_X1 U3795 ( .A1(n17403), .A2(n14346), .B1(n17398), .B2(n16802), .ZN(
        n9180) );
  OAI22_X1 U3796 ( .A1(n17467), .A2(n15539), .B1(n17463), .B2(n16802), .ZN(
        n9185) );
  OAI22_X1 U3797 ( .A1(n17493), .A2(n14805), .B1(n17489), .B2(n16802), .ZN(
        n9187) );
  OAI22_X1 U3798 ( .A1(n17506), .A2(n15626), .B1(n17502), .B2(n16802), .ZN(
        n9188) );
  OAI22_X1 U3799 ( .A1(n17066), .A2(n15171), .B1(n17062), .B2(n16805), .ZN(
        n9225) );
  OAI22_X1 U3800 ( .A1(n17092), .A2(n15513), .B1(n17088), .B2(n16806), .ZN(
        n9227) );
  OAI22_X1 U3801 ( .A1(n17105), .A2(n11863), .B1(n17101), .B2(n16806), .ZN(
        n9228) );
  OAI22_X1 U3802 ( .A1(n17259), .A2(n14849), .B1(n17255), .B2(n16807), .ZN(
        n9241) );
  OAI22_X1 U3803 ( .A1(n17285), .A2(n14409), .B1(n17281), .B2(n16807), .ZN(
        n9243) );
  OAI22_X1 U3804 ( .A1(n17298), .A2(n14623), .B1(n17294), .B2(n16807), .ZN(
        n9244) );
  OAI22_X1 U3805 ( .A1(n17363), .A2(n15687), .B1(n17359), .B2(n16807), .ZN(
        n9249) );
  OAI22_X1 U3806 ( .A1(n17389), .A2(n14749), .B1(n17385), .B2(n16808), .ZN(
        n9251) );
  OAI22_X1 U3807 ( .A1(n17402), .A2(n14347), .B1(n17398), .B2(n16808), .ZN(
        n9252) );
  OAI22_X1 U3808 ( .A1(n17467), .A2(n15540), .B1(n17463), .B2(n16808), .ZN(
        n9257) );
  OAI22_X1 U3809 ( .A1(n17493), .A2(n14807), .B1(n17489), .B2(n16808), .ZN(
        n9259) );
  OAI22_X1 U3810 ( .A1(n17506), .A2(n15627), .B1(n17502), .B2(n16808), .ZN(
        n9260) );
  OAI22_X1 U3811 ( .A1(n17066), .A2(n15172), .B1(n17062), .B2(n16811), .ZN(
        n9297) );
  OAI22_X1 U3812 ( .A1(n17092), .A2(n15514), .B1(n17088), .B2(n16812), .ZN(
        n9299) );
  OAI22_X1 U3813 ( .A1(n17105), .A2(n11864), .B1(n17101), .B2(n16812), .ZN(
        n9300) );
  OAI22_X1 U3814 ( .A1(n17259), .A2(n14850), .B1(n17255), .B2(n16813), .ZN(
        n9313) );
  OAI22_X1 U3815 ( .A1(n17285), .A2(n14410), .B1(n17281), .B2(n16813), .ZN(
        n9315) );
  OAI22_X1 U3816 ( .A1(n17298), .A2(n14624), .B1(n17294), .B2(n16813), .ZN(
        n9316) );
  OAI22_X1 U3817 ( .A1(n17363), .A2(n15688), .B1(n17359), .B2(n16813), .ZN(
        n9321) );
  OAI22_X1 U3818 ( .A1(n17389), .A2(n14751), .B1(n17385), .B2(n16814), .ZN(
        n9323) );
  OAI22_X1 U3819 ( .A1(n17402), .A2(n14348), .B1(n17398), .B2(n16814), .ZN(
        n9324) );
  OAI22_X1 U3820 ( .A1(n17467), .A2(n15541), .B1(n17463), .B2(n16814), .ZN(
        n9329) );
  OAI22_X1 U3821 ( .A1(n17493), .A2(n14809), .B1(n17489), .B2(n16814), .ZN(
        n9331) );
  OAI22_X1 U3822 ( .A1(n17506), .A2(n15628), .B1(n17502), .B2(n16814), .ZN(
        n9332) );
  OAI22_X1 U3823 ( .A1(n17066), .A2(n15173), .B1(n17062), .B2(n16817), .ZN(
        n9369) );
  OAI22_X1 U3824 ( .A1(n17092), .A2(n15515), .B1(n17088), .B2(n16818), .ZN(
        n9371) );
  OAI22_X1 U3825 ( .A1(n17105), .A2(n11865), .B1(n17101), .B2(n16818), .ZN(
        n9372) );
  OAI22_X1 U3826 ( .A1(n17259), .A2(n14851), .B1(n17255), .B2(n16819), .ZN(
        n9385) );
  OAI22_X1 U3827 ( .A1(n17285), .A2(n14411), .B1(n17281), .B2(n16819), .ZN(
        n9387) );
  OAI22_X1 U3828 ( .A1(n17298), .A2(n14625), .B1(n17294), .B2(n16819), .ZN(
        n9388) );
  OAI22_X1 U3829 ( .A1(n17363), .A2(n15689), .B1(n17359), .B2(n16819), .ZN(
        n9393) );
  OAI22_X1 U3830 ( .A1(n17389), .A2(n14753), .B1(n17385), .B2(n16820), .ZN(
        n9395) );
  OAI22_X1 U3831 ( .A1(n17402), .A2(n14349), .B1(n17398), .B2(n16820), .ZN(
        n9396) );
  OAI22_X1 U3832 ( .A1(n17467), .A2(n15542), .B1(n17463), .B2(n16820), .ZN(
        n9401) );
  OAI22_X1 U3833 ( .A1(n17493), .A2(n14811), .B1(n17489), .B2(n16820), .ZN(
        n9403) );
  OAI22_X1 U3834 ( .A1(n17506), .A2(n15629), .B1(n17502), .B2(n16820), .ZN(
        n9404) );
  OAI22_X1 U3835 ( .A1(n17066), .A2(n15174), .B1(n17062), .B2(n16823), .ZN(
        n9441) );
  OAI22_X1 U3836 ( .A1(n17092), .A2(n15516), .B1(n17088), .B2(n16824), .ZN(
        n9443) );
  OAI22_X1 U3837 ( .A1(n17105), .A2(n11866), .B1(n17101), .B2(n16824), .ZN(
        n9444) );
  OAI22_X1 U3838 ( .A1(n17259), .A2(n14852), .B1(n17255), .B2(n16825), .ZN(
        n9457) );
  OAI22_X1 U3839 ( .A1(n17285), .A2(n14412), .B1(n17281), .B2(n16825), .ZN(
        n9459) );
  OAI22_X1 U3840 ( .A1(n17298), .A2(n14626), .B1(n17294), .B2(n16825), .ZN(
        n9460) );
  OAI22_X1 U3841 ( .A1(n17362), .A2(n15690), .B1(n17359), .B2(n16825), .ZN(
        n9465) );
  OAI22_X1 U3842 ( .A1(n17388), .A2(n14755), .B1(n17385), .B2(n16826), .ZN(
        n9467) );
  OAI22_X1 U3843 ( .A1(n17401), .A2(n14350), .B1(n17398), .B2(n16826), .ZN(
        n9468) );
  OAI22_X1 U3844 ( .A1(n17466), .A2(n15543), .B1(n17463), .B2(n16826), .ZN(
        n9473) );
  OAI22_X1 U3845 ( .A1(n17492), .A2(n14813), .B1(n17489), .B2(n16826), .ZN(
        n9475) );
  OAI22_X1 U3846 ( .A1(n17505), .A2(n15630), .B1(n17502), .B2(n16826), .ZN(
        n9476) );
  OAI22_X1 U3847 ( .A1(n17065), .A2(n15175), .B1(n17062), .B2(n16829), .ZN(
        n9513) );
  OAI22_X1 U3848 ( .A1(n17091), .A2(n15488), .B1(n17088), .B2(n16830), .ZN(
        n9515) );
  OAI22_X1 U3849 ( .A1(n17104), .A2(n11867), .B1(n17101), .B2(n16830), .ZN(
        n9516) );
  OAI22_X1 U3850 ( .A1(n17258), .A2(n14824), .B1(n17255), .B2(n16831), .ZN(
        n9529) );
  OAI22_X1 U3851 ( .A1(n17284), .A2(n14413), .B1(n17281), .B2(n16831), .ZN(
        n9531) );
  OAI22_X1 U3852 ( .A1(n17297), .A2(n14598), .B1(n17294), .B2(n16831), .ZN(
        n9532) );
  OAI22_X1 U3853 ( .A1(n17362), .A2(n15662), .B1(n17359), .B2(n16831), .ZN(
        n9537) );
  OAI22_X1 U3854 ( .A1(n17388), .A2(n14700), .B1(n17385), .B2(n16832), .ZN(
        n9539) );
  OAI22_X1 U3855 ( .A1(n17401), .A2(n14351), .B1(n17398), .B2(n16832), .ZN(
        n9540) );
  OAI22_X1 U3856 ( .A1(n17466), .A2(n15544), .B1(n17463), .B2(n16832), .ZN(
        n9545) );
  OAI22_X1 U3857 ( .A1(n17492), .A2(n14757), .B1(n17489), .B2(n16832), .ZN(
        n9547) );
  OAI22_X1 U3858 ( .A1(n17505), .A2(n15631), .B1(n17502), .B2(n16832), .ZN(
        n9548) );
  OAI22_X1 U3859 ( .A1(n17065), .A2(n15176), .B1(n17062), .B2(n16835), .ZN(
        n9585) );
  OAI22_X1 U3860 ( .A1(n17091), .A2(n15489), .B1(n17088), .B2(n16836), .ZN(
        n9587) );
  OAI22_X1 U3861 ( .A1(n17104), .A2(n11869), .B1(n17101), .B2(n16836), .ZN(
        n9588) );
  OAI22_X1 U3862 ( .A1(n17258), .A2(n14825), .B1(n17255), .B2(n16837), .ZN(
        n9601) );
  OAI22_X1 U3863 ( .A1(n17284), .A2(n14414), .B1(n17281), .B2(n16837), .ZN(
        n9603) );
  OAI22_X1 U3864 ( .A1(n17297), .A2(n14599), .B1(n17294), .B2(n16837), .ZN(
        n9604) );
  OAI22_X1 U3865 ( .A1(n17363), .A2(n15663), .B1(n17359), .B2(n16837), .ZN(
        n9609) );
  OAI22_X1 U3866 ( .A1(n17389), .A2(n14701), .B1(n17385), .B2(n16838), .ZN(
        n9611) );
  OAI22_X1 U3867 ( .A1(n17402), .A2(n14352), .B1(n17398), .B2(n16838), .ZN(
        n9612) );
  OAI22_X1 U3868 ( .A1(n17466), .A2(n15452), .B1(n17463), .B2(n16838), .ZN(
        n9617) );
  OAI22_X1 U3869 ( .A1(n17492), .A2(n14759), .B1(n17489), .B2(n16838), .ZN(
        n9619) );
  OAI22_X1 U3870 ( .A1(n17505), .A2(n15632), .B1(n17502), .B2(n16838), .ZN(
        n9620) );
  OAI22_X1 U3871 ( .A1(n17065), .A2(n15177), .B1(n17062), .B2(n16841), .ZN(
        n9657) );
  OAI22_X1 U3872 ( .A1(n17091), .A2(n15490), .B1(n17088), .B2(n16842), .ZN(
        n9659) );
  OAI22_X1 U3873 ( .A1(n17104), .A2(n11870), .B1(n17101), .B2(n16842), .ZN(
        n9660) );
  OAI22_X1 U3874 ( .A1(n17258), .A2(n14826), .B1(n17255), .B2(n16843), .ZN(
        n9673) );
  OAI22_X1 U3875 ( .A1(n17284), .A2(n14415), .B1(n17281), .B2(n16843), .ZN(
        n9675) );
  OAI22_X1 U3876 ( .A1(n17297), .A2(n14600), .B1(n17294), .B2(n16843), .ZN(
        n9676) );
  OAI22_X1 U3877 ( .A1(n17362), .A2(n15664), .B1(n17359), .B2(n16843), .ZN(
        n9681) );
  OAI22_X1 U3878 ( .A1(n17388), .A2(n14702), .B1(n17385), .B2(n16844), .ZN(
        n9683) );
  OAI22_X1 U3879 ( .A1(n17401), .A2(n14353), .B1(n17398), .B2(n16844), .ZN(
        n9684) );
  OAI22_X1 U3880 ( .A1(n17466), .A2(n15453), .B1(n17463), .B2(n16844), .ZN(
        n9689) );
  OAI22_X1 U3881 ( .A1(n17492), .A2(n14761), .B1(n17489), .B2(n16844), .ZN(
        n9691) );
  OAI22_X1 U3882 ( .A1(n17505), .A2(n15633), .B1(n17502), .B2(n16844), .ZN(
        n9692) );
  OAI22_X1 U3883 ( .A1(n17065), .A2(n15178), .B1(n17062), .B2(n16847), .ZN(
        n9729) );
  OAI22_X1 U3884 ( .A1(n17091), .A2(n15491), .B1(n17088), .B2(n16848), .ZN(
        n9731) );
  OAI22_X1 U3885 ( .A1(n17104), .A2(n11871), .B1(n17101), .B2(n16848), .ZN(
        n9732) );
  OAI22_X1 U3886 ( .A1(n17258), .A2(n14827), .B1(n17255), .B2(n16849), .ZN(
        n9745) );
  OAI22_X1 U3887 ( .A1(n17284), .A2(n14416), .B1(n17281), .B2(n16849), .ZN(
        n9747) );
  OAI22_X1 U3888 ( .A1(n17297), .A2(n14601), .B1(n17294), .B2(n16849), .ZN(
        n9748) );
  OAI22_X1 U3889 ( .A1(n17362), .A2(n15665), .B1(n17359), .B2(n16849), .ZN(
        n9753) );
  OAI22_X1 U3890 ( .A1(n17388), .A2(n14704), .B1(n17385), .B2(n16850), .ZN(
        n9755) );
  OAI22_X1 U3891 ( .A1(n17401), .A2(n14354), .B1(n17398), .B2(n16850), .ZN(
        n9756) );
  OAI22_X1 U3892 ( .A1(n17465), .A2(n15454), .B1(n17463), .B2(n16850), .ZN(
        n9761) );
  OAI22_X1 U3893 ( .A1(n17491), .A2(n14763), .B1(n17489), .B2(n16850), .ZN(
        n9763) );
  OAI22_X1 U3894 ( .A1(n17504), .A2(n15634), .B1(n17502), .B2(n16850), .ZN(
        n9764) );
  OAI22_X1 U3895 ( .A1(n17064), .A2(n15179), .B1(n17062), .B2(n16853), .ZN(
        n9801) );
  OAI22_X1 U3896 ( .A1(n17090), .A2(n15492), .B1(n17088), .B2(n16854), .ZN(
        n9803) );
  OAI22_X1 U3897 ( .A1(n17103), .A2(n11872), .B1(n17101), .B2(n16854), .ZN(
        n9804) );
  OAI22_X1 U3898 ( .A1(n17257), .A2(n14828), .B1(n17255), .B2(n16855), .ZN(
        n9817) );
  OAI22_X1 U3899 ( .A1(n17283), .A2(n14417), .B1(n17281), .B2(n16855), .ZN(
        n9819) );
  OAI22_X1 U3900 ( .A1(n17296), .A2(n14602), .B1(n17294), .B2(n16855), .ZN(
        n9820) );
  OAI22_X1 U3901 ( .A1(n17361), .A2(n15666), .B1(n17359), .B2(n16855), .ZN(
        n9825) );
  OAI22_X1 U3902 ( .A1(n17387), .A2(n14706), .B1(n17385), .B2(n16856), .ZN(
        n9827) );
  OAI22_X1 U3903 ( .A1(n17400), .A2(n14355), .B1(n17398), .B2(n16856), .ZN(
        n9828) );
  OAI22_X1 U3904 ( .A1(n17465), .A2(n15455), .B1(n17463), .B2(n16856), .ZN(
        n9833) );
  OAI22_X1 U3905 ( .A1(n17491), .A2(n14765), .B1(n17489), .B2(n16856), .ZN(
        n9835) );
  OAI22_X1 U3906 ( .A1(n17504), .A2(n15635), .B1(n17502), .B2(n16856), .ZN(
        n9836) );
  OAI22_X1 U3907 ( .A1(n17064), .A2(n15180), .B1(n17062), .B2(n16859), .ZN(
        n9873) );
  OAI22_X1 U3908 ( .A1(n17090), .A2(n15493), .B1(n17088), .B2(n16860), .ZN(
        n9875) );
  OAI22_X1 U3909 ( .A1(n17103), .A2(n11873), .B1(n17101), .B2(n16860), .ZN(
        n9876) );
  OAI22_X1 U3910 ( .A1(n17257), .A2(n14829), .B1(n17255), .B2(n16861), .ZN(
        n9889) );
  OAI22_X1 U3911 ( .A1(n17283), .A2(n14418), .B1(n17281), .B2(n16861), .ZN(
        n9891) );
  OAI22_X1 U3912 ( .A1(n17296), .A2(n14603), .B1(n17294), .B2(n16861), .ZN(
        n9892) );
  OAI22_X1 U3913 ( .A1(n17361), .A2(n15667), .B1(n17359), .B2(n16861), .ZN(
        n9897) );
  OAI22_X1 U3914 ( .A1(n17387), .A2(n14708), .B1(n17385), .B2(n16862), .ZN(
        n9899) );
  OAI22_X1 U3915 ( .A1(n17400), .A2(n14356), .B1(n17398), .B2(n16862), .ZN(
        n9900) );
  OAI22_X1 U3916 ( .A1(n17465), .A2(n15456), .B1(n17463), .B2(n16862), .ZN(
        n9905) );
  OAI22_X1 U3917 ( .A1(n17491), .A2(n14767), .B1(n17489), .B2(n16862), .ZN(
        n9907) );
  OAI22_X1 U3918 ( .A1(n17504), .A2(n15636), .B1(n17502), .B2(n16862), .ZN(
        n9908) );
  OAI22_X1 U3919 ( .A1(n17122), .A2(n12315), .B1(n17115), .B2(n16727), .ZN(
        n8293) );
  OAI22_X1 U3920 ( .A1(n17315), .A2(n15704), .B1(n17308), .B2(n16728), .ZN(
        n8309) );
  OAI22_X1 U3921 ( .A1(n17419), .A2(n15215), .B1(n17412), .B2(n16729), .ZN(
        n8317) );
  OAI22_X1 U3922 ( .A1(n17122), .A2(n12316), .B1(n17115), .B2(n16734), .ZN(
        n8365) );
  OAI22_X1 U3923 ( .A1(n17315), .A2(n15705), .B1(n17308), .B2(n16735), .ZN(
        n8381) );
  OAI22_X1 U3924 ( .A1(n17419), .A2(n15216), .B1(n17412), .B2(n16736), .ZN(
        n8389) );
  OAI22_X1 U3925 ( .A1(n17121), .A2(n12317), .B1(n17115), .B2(n16740), .ZN(
        n8437) );
  OAI22_X1 U3926 ( .A1(n17314), .A2(n15706), .B1(n17308), .B2(n16741), .ZN(
        n8453) );
  OAI22_X1 U3927 ( .A1(n17418), .A2(n15217), .B1(n17412), .B2(n16742), .ZN(
        n8461) );
  OAI22_X1 U3928 ( .A1(n17121), .A2(n12318), .B1(n17115), .B2(n16746), .ZN(
        n8509) );
  OAI22_X1 U3929 ( .A1(n17314), .A2(n15707), .B1(n17308), .B2(n16747), .ZN(
        n8525) );
  OAI22_X1 U3930 ( .A1(n17418), .A2(n15218), .B1(n17412), .B2(n16748), .ZN(
        n8533) );
  OAI22_X1 U3931 ( .A1(n17121), .A2(n12319), .B1(n17115), .B2(n16752), .ZN(
        n8581) );
  OAI22_X1 U3932 ( .A1(n17314), .A2(n15708), .B1(n17308), .B2(n16753), .ZN(
        n8597) );
  OAI22_X1 U3933 ( .A1(n17418), .A2(n15219), .B1(n17412), .B2(n16754), .ZN(
        n8605) );
  OAI22_X1 U3934 ( .A1(n17121), .A2(n12320), .B1(n17115), .B2(n16758), .ZN(
        n8653) );
  OAI22_X1 U3935 ( .A1(n17314), .A2(n15709), .B1(n17308), .B2(n16759), .ZN(
        n8669) );
  OAI22_X1 U3936 ( .A1(n17418), .A2(n15220), .B1(n17412), .B2(n16760), .ZN(
        n8677) );
  OAI22_X1 U3937 ( .A1(n17120), .A2(n12321), .B1(n17115), .B2(n16764), .ZN(
        n8725) );
  OAI22_X1 U3938 ( .A1(n17313), .A2(n15710), .B1(n17308), .B2(n16765), .ZN(
        n8741) );
  OAI22_X1 U3939 ( .A1(n17417), .A2(n15221), .B1(n17412), .B2(n16766), .ZN(
        n8749) );
  OAI22_X1 U3940 ( .A1(n17120), .A2(n12322), .B1(n17115), .B2(n16770), .ZN(
        n8797) );
  OAI22_X1 U3941 ( .A1(n17313), .A2(n15711), .B1(n17308), .B2(n16771), .ZN(
        n8813) );
  OAI22_X1 U3942 ( .A1(n17417), .A2(n15222), .B1(n17412), .B2(n16772), .ZN(
        n8821) );
  OAI22_X1 U3943 ( .A1(n17120), .A2(n12323), .B1(n17115), .B2(n16776), .ZN(
        n8869) );
  OAI22_X1 U3944 ( .A1(n17313), .A2(n15712), .B1(n17308), .B2(n16777), .ZN(
        n8885) );
  OAI22_X1 U3945 ( .A1(n17417), .A2(n15223), .B1(n17412), .B2(n16778), .ZN(
        n8893) );
  OAI22_X1 U3946 ( .A1(n17119), .A2(n12324), .B1(n17115), .B2(n16782), .ZN(
        n8941) );
  OAI22_X1 U3947 ( .A1(n17312), .A2(n15713), .B1(n17308), .B2(n16783), .ZN(
        n8957) );
  OAI22_X1 U3948 ( .A1(n17416), .A2(n15224), .B1(n17412), .B2(n16784), .ZN(
        n8965) );
  OAI22_X1 U3949 ( .A1(n17119), .A2(n12325), .B1(n17115), .B2(n16788), .ZN(
        n9013) );
  OAI22_X1 U3950 ( .A1(n17312), .A2(n15714), .B1(n17308), .B2(n16789), .ZN(
        n9029) );
  OAI22_X1 U3951 ( .A1(n17416), .A2(n15225), .B1(n17412), .B2(n16790), .ZN(
        n9037) );
  OAI22_X1 U3952 ( .A1(n17119), .A2(n12326), .B1(n17114), .B2(n16794), .ZN(
        n9085) );
  OAI22_X1 U3953 ( .A1(n17312), .A2(n15715), .B1(n17307), .B2(n16795), .ZN(
        n9101) );
  OAI22_X1 U3954 ( .A1(n17416), .A2(n15226), .B1(n17411), .B2(n16796), .ZN(
        n9109) );
  OAI22_X1 U3955 ( .A1(n17119), .A2(n12327), .B1(n17114), .B2(n16800), .ZN(
        n9157) );
  OAI22_X1 U3956 ( .A1(n17312), .A2(n15716), .B1(n17307), .B2(n16801), .ZN(
        n9173) );
  OAI22_X1 U3957 ( .A1(n17416), .A2(n15227), .B1(n17411), .B2(n16802), .ZN(
        n9181) );
  OAI22_X1 U3958 ( .A1(n17118), .A2(n12328), .B1(n17114), .B2(n16806), .ZN(
        n9229) );
  OAI22_X1 U3959 ( .A1(n17311), .A2(n15717), .B1(n17307), .B2(n16807), .ZN(
        n9245) );
  OAI22_X1 U3960 ( .A1(n17415), .A2(n15228), .B1(n17411), .B2(n16808), .ZN(
        n9253) );
  OAI22_X1 U3961 ( .A1(n17118), .A2(n12329), .B1(n17114), .B2(n16812), .ZN(
        n9301) );
  OAI22_X1 U3962 ( .A1(n17311), .A2(n15718), .B1(n17307), .B2(n16813), .ZN(
        n9317) );
  OAI22_X1 U3963 ( .A1(n17415), .A2(n15229), .B1(n17411), .B2(n16814), .ZN(
        n9325) );
  OAI22_X1 U3964 ( .A1(n17118), .A2(n12330), .B1(n17114), .B2(n16818), .ZN(
        n9373) );
  OAI22_X1 U3965 ( .A1(n17311), .A2(n15719), .B1(n17307), .B2(n16819), .ZN(
        n9389) );
  OAI22_X1 U3966 ( .A1(n17415), .A2(n15230), .B1(n17411), .B2(n16820), .ZN(
        n9397) );
  OAI22_X1 U3967 ( .A1(n17118), .A2(n12331), .B1(n17114), .B2(n16824), .ZN(
        n9445) );
  OAI22_X1 U3968 ( .A1(n17311), .A2(n15720), .B1(n17307), .B2(n16825), .ZN(
        n9461) );
  OAI22_X1 U3969 ( .A1(n17414), .A2(n15231), .B1(n17411), .B2(n16826), .ZN(
        n9469) );
  OAI22_X1 U3970 ( .A1(n17117), .A2(n12332), .B1(n17114), .B2(n16830), .ZN(
        n9517) );
  OAI22_X1 U3971 ( .A1(n17310), .A2(n15692), .B1(n17307), .B2(n16831), .ZN(
        n9533) );
  OAI22_X1 U3972 ( .A1(n17414), .A2(n15232), .B1(n17411), .B2(n16832), .ZN(
        n9541) );
  OAI22_X1 U3973 ( .A1(n17117), .A2(n12333), .B1(n17114), .B2(n16836), .ZN(
        n9589) );
  OAI22_X1 U3974 ( .A1(n17310), .A2(n15693), .B1(n17307), .B2(n16837), .ZN(
        n9605) );
  OAI22_X1 U3975 ( .A1(n17415), .A2(n15233), .B1(n17411), .B2(n16838), .ZN(
        n9613) );
  OAI22_X1 U3976 ( .A1(n17117), .A2(n12334), .B1(n17114), .B2(n16842), .ZN(
        n9661) );
  OAI22_X1 U3977 ( .A1(n17310), .A2(n15694), .B1(n17307), .B2(n16843), .ZN(
        n9677) );
  OAI22_X1 U3978 ( .A1(n17414), .A2(n15234), .B1(n17411), .B2(n16844), .ZN(
        n9685) );
  OAI22_X1 U3979 ( .A1(n17117), .A2(n12335), .B1(n17114), .B2(n16848), .ZN(
        n9733) );
  OAI22_X1 U3980 ( .A1(n17310), .A2(n15695), .B1(n17307), .B2(n16849), .ZN(
        n9749) );
  OAI22_X1 U3981 ( .A1(n17414), .A2(n15235), .B1(n17411), .B2(n16850), .ZN(
        n9757) );
  OAI22_X1 U3982 ( .A1(n17116), .A2(n12336), .B1(n17114), .B2(n16854), .ZN(
        n9805) );
  OAI22_X1 U3983 ( .A1(n17309), .A2(n15696), .B1(n17307), .B2(n16855), .ZN(
        n9821) );
  OAI22_X1 U3984 ( .A1(n17413), .A2(n15236), .B1(n17411), .B2(n16856), .ZN(
        n9829) );
  OAI22_X1 U3985 ( .A1(n17116), .A2(n12337), .B1(n17114), .B2(n16860), .ZN(
        n9877) );
  OAI22_X1 U3986 ( .A1(n17309), .A2(n15697), .B1(n17307), .B2(n16861), .ZN(
        n9893) );
  OAI22_X1 U3987 ( .A1(n17413), .A2(n15237), .B1(n17411), .B2(n16862), .ZN(
        n9901) );
  OAI22_X1 U3988 ( .A1(n17120), .A2(n12339), .B1(n17115), .B2(n17515), .ZN(
        n9949) );
  OAI22_X1 U3989 ( .A1(n17313), .A2(n15698), .B1(n17308), .B2(n17516), .ZN(
        n9965) );
  OAI22_X1 U3990 ( .A1(n17417), .A2(n15238), .B1(n17412), .B2(n17517), .ZN(
        n9973) );
  INV_X1 U3991 ( .A(N9926), .ZN(n14174) );
  OAI22_X1 U3992 ( .A1(n16885), .A2(n18031), .B1(n14855), .B2(n4462), .ZN(
        n10001) );
  OAI22_X1 U3993 ( .A1(n16895), .A2(n18031), .B1(n15272), .B2(n4459), .ZN(
        n10002) );
  OAI22_X1 U3994 ( .A1(n16918), .A2(n18031), .B1(n14065), .B2(n4451), .ZN(
        n10004) );
  OAI22_X1 U3995 ( .A1(n16953), .A2(n18031), .B1(n11670), .B2(n4438), .ZN(
        n10007) );
  OAI22_X1 U3996 ( .A1(n16964), .A2(n18031), .B1(n14631), .B2(n4435), .ZN(
        n10008) );
  OAI22_X1 U3997 ( .A1(n16974), .A2(n18031), .B1(n15275), .B2(n16966), .ZN(
        n10009) );
  OAI22_X1 U3998 ( .A1(n16984), .A2(n18031), .B1(n14854), .B2(n4429), .ZN(
        n10010) );
  OAI22_X1 U3999 ( .A1(n17007), .A2(n18030), .B1(n14069), .B2(n16999), .ZN(
        n10012) );
  OAI22_X1 U4000 ( .A1(n17145), .A2(n18030), .B1(n14628), .B2(n4382), .ZN(
        n10023) );
  OAI22_X1 U4001 ( .A1(n17168), .A2(n18029), .B1(n14857), .B2(n4376), .ZN(
        n10025) );
  OAI22_X1 U4002 ( .A1(n17179), .A2(n18029), .B1(n11904), .B2(n4373), .ZN(
        n10026) );
  OAI22_X1 U4003 ( .A1(n17190), .A2(n18029), .B1(n12197), .B2(n4370), .ZN(
        n10027) );
  OAI22_X1 U4004 ( .A1(n17200), .A2(n18029), .B1(n14054), .B2(n4367), .ZN(
        n10028) );
  INV_X1 U4005 ( .A(N9922), .ZN(n14173) );
  INV_X1 U4006 ( .A(n14178), .ZN(n14003) );
  OAI22_X1 U4007 ( .A1(n17944), .A2(n14886), .B1(n17947), .B2(n17513), .ZN(
        n9923) );
  OAI22_X1 U4008 ( .A1(n17965), .A2(n15269), .B1(n17968), .B2(n17513), .ZN(
        n9924) );
  OAI22_X1 U4009 ( .A1(n17836), .A2(n14483), .B1(n17840), .B2(n17512), .ZN(
        n9918) );
  OAI22_X1 U4010 ( .A1(n17902), .A2(n14644), .B1(n17905), .B2(n17512), .ZN(
        n9921) );
  OAI22_X1 U4011 ( .A1(n17946), .A2(n14912), .B1(n17959), .B2(n16448), .ZN(
        n7917) );
  OAI22_X1 U4012 ( .A1(n17967), .A2(n15244), .B1(n17980), .B2(n16448), .ZN(
        n7918) );
  OAI22_X1 U4013 ( .A1(n17925), .A2(n15435), .B1(n17938), .B2(n16725), .ZN(
        n8266) );
  OAI22_X1 U4014 ( .A1(n17946), .A2(n14913), .B1(n17958), .B2(n16725), .ZN(
        n8267) );
  OAI22_X1 U4015 ( .A1(n17967), .A2(n15246), .B1(n17979), .B2(n16725), .ZN(
        n8268) );
  OAI22_X1 U4016 ( .A1(n17925), .A2(n15436), .B1(n17938), .B2(n16732), .ZN(
        n8338) );
  OAI22_X1 U4017 ( .A1(n17946), .A2(n14914), .B1(n17959), .B2(n16732), .ZN(
        n8339) );
  OAI22_X1 U4018 ( .A1(n17967), .A2(n15247), .B1(n17980), .B2(n16732), .ZN(
        n8340) );
  OAI22_X1 U4019 ( .A1(n17925), .A2(n15437), .B1(n17937), .B2(n16738), .ZN(
        n8410) );
  OAI22_X1 U4020 ( .A1(n17946), .A2(n14915), .B1(n17957), .B2(n16738), .ZN(
        n8411) );
  OAI22_X1 U4021 ( .A1(n17967), .A2(n15248), .B1(n17978), .B2(n16738), .ZN(
        n8412) );
  OAI22_X1 U4022 ( .A1(n17925), .A2(n15438), .B1(n17937), .B2(n16744), .ZN(
        n8482) );
  OAI22_X1 U4023 ( .A1(n17946), .A2(n14916), .B1(n17958), .B2(n16744), .ZN(
        n8483) );
  OAI22_X1 U4024 ( .A1(n17967), .A2(n15249), .B1(n17979), .B2(n16744), .ZN(
        n8484) );
  OAI22_X1 U4025 ( .A1(n17924), .A2(n15439), .B1(n17936), .B2(n16750), .ZN(
        n8554) );
  OAI22_X1 U4026 ( .A1(n17945), .A2(n14917), .B1(n17956), .B2(n16750), .ZN(
        n8555) );
  OAI22_X1 U4027 ( .A1(n17966), .A2(n15250), .B1(n17977), .B2(n16750), .ZN(
        n8556) );
  OAI22_X1 U4028 ( .A1(n17924), .A2(n15440), .B1(n17936), .B2(n16756), .ZN(
        n8626) );
  OAI22_X1 U4029 ( .A1(n17945), .A2(n14918), .B1(n17957), .B2(n16756), .ZN(
        n8627) );
  OAI22_X1 U4030 ( .A1(n17966), .A2(n15251), .B1(n17978), .B2(n16756), .ZN(
        n8628) );
  OAI22_X1 U4031 ( .A1(n17924), .A2(n15441), .B1(n17935), .B2(n16762), .ZN(
        n8698) );
  OAI22_X1 U4032 ( .A1(n17945), .A2(n14919), .B1(n17955), .B2(n16762), .ZN(
        n8699) );
  OAI22_X1 U4033 ( .A1(n17966), .A2(n15252), .B1(n17976), .B2(n16762), .ZN(
        n8700) );
  OAI22_X1 U4034 ( .A1(n17924), .A2(n15442), .B1(n17935), .B2(n16768), .ZN(
        n8770) );
  OAI22_X1 U4035 ( .A1(n17945), .A2(n14920), .B1(n17956), .B2(n16768), .ZN(
        n8771) );
  OAI22_X1 U4036 ( .A1(n17966), .A2(n15253), .B1(n17977), .B2(n16768), .ZN(
        n8772) );
  OAI22_X1 U4037 ( .A1(n17924), .A2(n15443), .B1(n17934), .B2(n16774), .ZN(
        n8842) );
  OAI22_X1 U4038 ( .A1(n17945), .A2(n14921), .B1(n17955), .B2(n16774), .ZN(
        n8843) );
  OAI22_X1 U4039 ( .A1(n17966), .A2(n15254), .B1(n17976), .B2(n16774), .ZN(
        n8844) );
  OAI22_X1 U4040 ( .A1(n17924), .A2(n15444), .B1(n17934), .B2(n16780), .ZN(
        n8914) );
  OAI22_X1 U4041 ( .A1(n17945), .A2(n14922), .B1(n17954), .B2(n16780), .ZN(
        n8915) );
  OAI22_X1 U4042 ( .A1(n17966), .A2(n15255), .B1(n17975), .B2(n16780), .ZN(
        n8916) );
  OAI22_X1 U4043 ( .A1(n17924), .A2(n15445), .B1(n17933), .B2(n16786), .ZN(
        n8986) );
  OAI22_X1 U4044 ( .A1(n17945), .A2(n14923), .B1(n17954), .B2(n16786), .ZN(
        n8987) );
  OAI22_X1 U4045 ( .A1(n17966), .A2(n15256), .B1(n17975), .B2(n16786), .ZN(
        n8988) );
  OAI22_X1 U4046 ( .A1(n17924), .A2(n15446), .B1(n17933), .B2(n16792), .ZN(
        n9058) );
  OAI22_X1 U4047 ( .A1(n17945), .A2(n14924), .B1(n17953), .B2(n16792), .ZN(
        n9059) );
  OAI22_X1 U4048 ( .A1(n17966), .A2(n15257), .B1(n17974), .B2(n16792), .ZN(
        n9060) );
  OAI22_X1 U4049 ( .A1(n17924), .A2(n15447), .B1(n17932), .B2(n16798), .ZN(
        n9130) );
  OAI22_X1 U4050 ( .A1(n17945), .A2(n14925), .B1(n17953), .B2(n16798), .ZN(
        n9131) );
  OAI22_X1 U4051 ( .A1(n17966), .A2(n15258), .B1(n17974), .B2(n16798), .ZN(
        n9132) );
  OAI22_X1 U4052 ( .A1(n17924), .A2(n15448), .B1(n17932), .B2(n16804), .ZN(
        n9202) );
  OAI22_X1 U4053 ( .A1(n17945), .A2(n14926), .B1(n17952), .B2(n16804), .ZN(
        n9203) );
  OAI22_X1 U4054 ( .A1(n17966), .A2(n15259), .B1(n17973), .B2(n16804), .ZN(
        n9204) );
  OAI22_X1 U4055 ( .A1(n17924), .A2(n15449), .B1(n17931), .B2(n16810), .ZN(
        n9274) );
  OAI22_X1 U4056 ( .A1(n17945), .A2(n14927), .B1(n17952), .B2(n16810), .ZN(
        n9275) );
  OAI22_X1 U4057 ( .A1(n17966), .A2(n15260), .B1(n17973), .B2(n16810), .ZN(
        n9276) );
  OAI22_X1 U4058 ( .A1(n17924), .A2(n15450), .B1(n17931), .B2(n16816), .ZN(
        n9346) );
  OAI22_X1 U4059 ( .A1(n17945), .A2(n14928), .B1(n17951), .B2(n16816), .ZN(
        n9347) );
  OAI22_X1 U4060 ( .A1(n17966), .A2(n15261), .B1(n17972), .B2(n16816), .ZN(
        n9348) );
  OAI22_X1 U4061 ( .A1(n17924), .A2(n15451), .B1(n17930), .B2(n16822), .ZN(
        n9418) );
  OAI22_X1 U4062 ( .A1(n17945), .A2(n14929), .B1(n17951), .B2(n16822), .ZN(
        n9419) );
  OAI22_X1 U4063 ( .A1(n17966), .A2(n15262), .B1(n17972), .B2(n16822), .ZN(
        n9420) );
  OAI22_X1 U4064 ( .A1(n17923), .A2(n15518), .B1(n17930), .B2(n16828), .ZN(
        n9490) );
  OAI22_X1 U4065 ( .A1(n17944), .A2(n14930), .B1(n17950), .B2(n16828), .ZN(
        n9491) );
  OAI22_X1 U4066 ( .A1(n17965), .A2(n15263), .B1(n17971), .B2(n16828), .ZN(
        n9492) );
  OAI22_X1 U4067 ( .A1(n17923), .A2(n15519), .B1(n17929), .B2(n16834), .ZN(
        n9562) );
  OAI22_X1 U4068 ( .A1(n17944), .A2(n14876), .B1(n17950), .B2(n16834), .ZN(
        n9563) );
  OAI22_X1 U4069 ( .A1(n17965), .A2(n15264), .B1(n17971), .B2(n16834), .ZN(
        n9564) );
  OAI22_X1 U4070 ( .A1(n17923), .A2(n15520), .B1(n17929), .B2(n16840), .ZN(
        n9634) );
  OAI22_X1 U4071 ( .A1(n17944), .A2(n14878), .B1(n17949), .B2(n16840), .ZN(
        n9635) );
  OAI22_X1 U4072 ( .A1(n17965), .A2(n15265), .B1(n17970), .B2(n16840), .ZN(
        n9636) );
  OAI22_X1 U4073 ( .A1(n17923), .A2(n15428), .B1(n17928), .B2(n16846), .ZN(
        n9706) );
  OAI22_X1 U4074 ( .A1(n17944), .A2(n14880), .B1(n17949), .B2(n16846), .ZN(
        n9707) );
  OAI22_X1 U4075 ( .A1(n17965), .A2(n15266), .B1(n17970), .B2(n16846), .ZN(
        n9708) );
  OAI22_X1 U4076 ( .A1(n17923), .A2(n15429), .B1(n17928), .B2(n16852), .ZN(
        n9778) );
  OAI22_X1 U4077 ( .A1(n17944), .A2(n14882), .B1(n17948), .B2(n16852), .ZN(
        n9779) );
  OAI22_X1 U4078 ( .A1(n17965), .A2(n15267), .B1(n17969), .B2(n16852), .ZN(
        n9780) );
  OAI22_X1 U4079 ( .A1(n17923), .A2(n15430), .B1(n17927), .B2(n16858), .ZN(
        n9850) );
  OAI22_X1 U4080 ( .A1(n17944), .A2(n14884), .B1(n17948), .B2(n16858), .ZN(
        n9851) );
  OAI22_X1 U4081 ( .A1(n17965), .A2(n15268), .B1(n17969), .B2(n16858), .ZN(
        n9852) );
  OAI22_X1 U4082 ( .A1(n17923), .A2(n15431), .B1(n17927), .B2(n17513), .ZN(
        n9922) );
  OAI22_X1 U4083 ( .A1(n17904), .A2(n14645), .B1(n17917), .B2(n16442), .ZN(
        n7841) );
  OAI22_X1 U4084 ( .A1(n17838), .A2(n14509), .B1(n17851), .B2(n16725), .ZN(
        n8262) );
  OAI22_X1 U4085 ( .A1(n17860), .A2(n15126), .B1(n17873), .B2(n16725), .ZN(
        n8263) );
  OAI22_X1 U4086 ( .A1(n17882), .A2(n15637), .B1(n17895), .B2(n16725), .ZN(
        n8264) );
  OAI22_X1 U4087 ( .A1(n17904), .A2(n14646), .B1(n17916), .B2(n16725), .ZN(
        n8265) );
  OAI22_X1 U4088 ( .A1(n17860), .A2(n15127), .B1(n17873), .B2(n16731), .ZN(
        n8335) );
  OAI22_X1 U4089 ( .A1(n17882), .A2(n15638), .B1(n17895), .B2(n16731), .ZN(
        n8336) );
  OAI22_X1 U4090 ( .A1(n17904), .A2(n14647), .B1(n17917), .B2(n16731), .ZN(
        n8337) );
  OAI22_X1 U4091 ( .A1(n17838), .A2(n14511), .B1(n17848), .B2(n16737), .ZN(
        n8406) );
  OAI22_X1 U4092 ( .A1(n17860), .A2(n15128), .B1(n17872), .B2(n16737), .ZN(
        n8407) );
  OAI22_X1 U4093 ( .A1(n17882), .A2(n15639), .B1(n17894), .B2(n16737), .ZN(
        n8408) );
  OAI22_X1 U4094 ( .A1(n17904), .A2(n14648), .B1(n17915), .B2(n16737), .ZN(
        n8409) );
  OAI22_X1 U4095 ( .A1(n17838), .A2(n14512), .B1(n17851), .B2(n16743), .ZN(
        n8478) );
  OAI22_X1 U4096 ( .A1(n17860), .A2(n15129), .B1(n17872), .B2(n16743), .ZN(
        n8479) );
  OAI22_X1 U4097 ( .A1(n17882), .A2(n15640), .B1(n17894), .B2(n16743), .ZN(
        n8480) );
  OAI22_X1 U4098 ( .A1(n17904), .A2(n14649), .B1(n17916), .B2(n16743), .ZN(
        n8481) );
  OAI22_X1 U4099 ( .A1(n17837), .A2(n14513), .B1(n17850), .B2(n16749), .ZN(
        n8550) );
  OAI22_X1 U4100 ( .A1(n17859), .A2(n15130), .B1(n17871), .B2(n16749), .ZN(
        n8551) );
  OAI22_X1 U4101 ( .A1(n17881), .A2(n15641), .B1(n17893), .B2(n16749), .ZN(
        n8552) );
  OAI22_X1 U4102 ( .A1(n17903), .A2(n14650), .B1(n17914), .B2(n16749), .ZN(
        n8553) );
  OAI22_X1 U4103 ( .A1(n17837), .A2(n14514), .B1(n17850), .B2(n16755), .ZN(
        n8622) );
  OAI22_X1 U4104 ( .A1(n17859), .A2(n15131), .B1(n17871), .B2(n16755), .ZN(
        n8623) );
  OAI22_X1 U4105 ( .A1(n17881), .A2(n15642), .B1(n17893), .B2(n16755), .ZN(
        n8624) );
  OAI22_X1 U4106 ( .A1(n17903), .A2(n14651), .B1(n17915), .B2(n16755), .ZN(
        n8625) );
  OAI22_X1 U4107 ( .A1(n17837), .A2(n14515), .B1(n17849), .B2(n16761), .ZN(
        n8694) );
  OAI22_X1 U4108 ( .A1(n17859), .A2(n15132), .B1(n17870), .B2(n16761), .ZN(
        n8695) );
  OAI22_X1 U4109 ( .A1(n17881), .A2(n15643), .B1(n17892), .B2(n16761), .ZN(
        n8696) );
  OAI22_X1 U4110 ( .A1(n17903), .A2(n14652), .B1(n17913), .B2(n16761), .ZN(
        n8697) );
  OAI22_X1 U4111 ( .A1(n17837), .A2(n14516), .B1(n17849), .B2(n16767), .ZN(
        n8766) );
  OAI22_X1 U4112 ( .A1(n17859), .A2(n15133), .B1(n17870), .B2(n16767), .ZN(
        n8767) );
  OAI22_X1 U4113 ( .A1(n17881), .A2(n15644), .B1(n17892), .B2(n16767), .ZN(
        n8768) );
  OAI22_X1 U4114 ( .A1(n17903), .A2(n14653), .B1(n17914), .B2(n16767), .ZN(
        n8769) );
  OAI22_X1 U4115 ( .A1(n17837), .A2(n14517), .B1(n17847), .B2(n16773), .ZN(
        n8838) );
  OAI22_X1 U4116 ( .A1(n17859), .A2(n15134), .B1(n17869), .B2(n16773), .ZN(
        n8839) );
  OAI22_X1 U4117 ( .A1(n17881), .A2(n15645), .B1(n17891), .B2(n16773), .ZN(
        n8840) );
  OAI22_X1 U4118 ( .A1(n17903), .A2(n14654), .B1(n17913), .B2(n16773), .ZN(
        n8841) );
  OAI22_X1 U4119 ( .A1(n17837), .A2(n14518), .B1(n17848), .B2(n16779), .ZN(
        n8910) );
  OAI22_X1 U4120 ( .A1(n17859), .A2(n15135), .B1(n17869), .B2(n16779), .ZN(
        n8911) );
  OAI22_X1 U4121 ( .A1(n17881), .A2(n15646), .B1(n17891), .B2(n16779), .ZN(
        n8912) );
  OAI22_X1 U4122 ( .A1(n17903), .A2(n14655), .B1(n17912), .B2(n16779), .ZN(
        n8913) );
  OAI22_X1 U4123 ( .A1(n17837), .A2(n14519), .B1(n17847), .B2(n16785), .ZN(
        n8982) );
  OAI22_X1 U4124 ( .A1(n17859), .A2(n15136), .B1(n17868), .B2(n16785), .ZN(
        n8983) );
  OAI22_X1 U4125 ( .A1(n17881), .A2(n15647), .B1(n17890), .B2(n16785), .ZN(
        n8984) );
  OAI22_X1 U4126 ( .A1(n17903), .A2(n14656), .B1(n17912), .B2(n16785), .ZN(
        n8985) );
  OAI22_X1 U4127 ( .A1(n17837), .A2(n14520), .B1(n17846), .B2(n16791), .ZN(
        n9054) );
  OAI22_X1 U4128 ( .A1(n17859), .A2(n15137), .B1(n17868), .B2(n16791), .ZN(
        n9055) );
  OAI22_X1 U4129 ( .A1(n17881), .A2(n15648), .B1(n17890), .B2(n16791), .ZN(
        n9056) );
  OAI22_X1 U4130 ( .A1(n17903), .A2(n14657), .B1(n17911), .B2(n16791), .ZN(
        n9057) );
  OAI22_X1 U4131 ( .A1(n17837), .A2(n14521), .B1(n17846), .B2(n16797), .ZN(
        n9126) );
  OAI22_X1 U4132 ( .A1(n17859), .A2(n15138), .B1(n17867), .B2(n16797), .ZN(
        n9127) );
  OAI22_X1 U4133 ( .A1(n17881), .A2(n15649), .B1(n17889), .B2(n16797), .ZN(
        n9128) );
  OAI22_X1 U4134 ( .A1(n17903), .A2(n14658), .B1(n17911), .B2(n16797), .ZN(
        n9129) );
  OAI22_X1 U4135 ( .A1(n17837), .A2(n14522), .B1(n17845), .B2(n16803), .ZN(
        n9198) );
  OAI22_X1 U4136 ( .A1(n17859), .A2(n15139), .B1(n17867), .B2(n16803), .ZN(
        n9199) );
  OAI22_X1 U4137 ( .A1(n17881), .A2(n15650), .B1(n17889), .B2(n16803), .ZN(
        n9200) );
  OAI22_X1 U4138 ( .A1(n17903), .A2(n14659), .B1(n17910), .B2(n16803), .ZN(
        n9201) );
  OAI22_X1 U4139 ( .A1(n17837), .A2(n14523), .B1(n17845), .B2(n16809), .ZN(
        n9270) );
  OAI22_X1 U4140 ( .A1(n17859), .A2(n15140), .B1(n17866), .B2(n16809), .ZN(
        n9271) );
  OAI22_X1 U4141 ( .A1(n17881), .A2(n15651), .B1(n17888), .B2(n16809), .ZN(
        n9272) );
  OAI22_X1 U4142 ( .A1(n17903), .A2(n14660), .B1(n17910), .B2(n16809), .ZN(
        n9273) );
  OAI22_X1 U4143 ( .A1(n17837), .A2(n14524), .B1(n17844), .B2(n16815), .ZN(
        n9342) );
  OAI22_X1 U4144 ( .A1(n17859), .A2(n15141), .B1(n17866), .B2(n16815), .ZN(
        n9343) );
  OAI22_X1 U4145 ( .A1(n17881), .A2(n15652), .B1(n17888), .B2(n16815), .ZN(
        n9344) );
  OAI22_X1 U4146 ( .A1(n17903), .A2(n14661), .B1(n17909), .B2(n16815), .ZN(
        n9345) );
  OAI22_X1 U4147 ( .A1(n17837), .A2(n14525), .B1(n17844), .B2(n16821), .ZN(
        n9414) );
  OAI22_X1 U4148 ( .A1(n17859), .A2(n15142), .B1(n17865), .B2(n16821), .ZN(
        n9415) );
  OAI22_X1 U4149 ( .A1(n17881), .A2(n15653), .B1(n17887), .B2(n16821), .ZN(
        n9416) );
  OAI22_X1 U4150 ( .A1(n17903), .A2(n14662), .B1(n17909), .B2(n16821), .ZN(
        n9417) );
  OAI22_X1 U4151 ( .A1(n17836), .A2(n14526), .B1(n17843), .B2(n16827), .ZN(
        n9486) );
  OAI22_X1 U4152 ( .A1(n17858), .A2(n15143), .B1(n17865), .B2(n16827), .ZN(
        n9487) );
  OAI22_X1 U4153 ( .A1(n17880), .A2(n15654), .B1(n17887), .B2(n16827), .ZN(
        n9488) );
  OAI22_X1 U4154 ( .A1(n17902), .A2(n14663), .B1(n17908), .B2(n16827), .ZN(
        n9489) );
  OAI22_X1 U4155 ( .A1(n17836), .A2(n14478), .B1(n17843), .B2(n16833), .ZN(
        n9558) );
  OAI22_X1 U4156 ( .A1(n17858), .A2(n15117), .B1(n17864), .B2(n16833), .ZN(
        n9559) );
  OAI22_X1 U4157 ( .A1(n17880), .A2(n15655), .B1(n17886), .B2(n16833), .ZN(
        n9560) );
  OAI22_X1 U4158 ( .A1(n17902), .A2(n14664), .B1(n17908), .B2(n16833), .ZN(
        n9561) );
  OAI22_X1 U4159 ( .A1(n17836), .A2(n14479), .B1(n17842), .B2(n16839), .ZN(
        n9630) );
  OAI22_X1 U4160 ( .A1(n17858), .A2(n15118), .B1(n17864), .B2(n16839), .ZN(
        n9631) );
  OAI22_X1 U4161 ( .A1(n17880), .A2(n15656), .B1(n17886), .B2(n16839), .ZN(
        n9632) );
  OAI22_X1 U4162 ( .A1(n17902), .A2(n14665), .B1(n17907), .B2(n16839), .ZN(
        n9633) );
  OAI22_X1 U4163 ( .A1(n17836), .A2(n14480), .B1(n17842), .B2(n16845), .ZN(
        n9702) );
  OAI22_X1 U4164 ( .A1(n17858), .A2(n15119), .B1(n17863), .B2(n16845), .ZN(
        n9703) );
  OAI22_X1 U4165 ( .A1(n17880), .A2(n15657), .B1(n17885), .B2(n16845), .ZN(
        n9704) );
  OAI22_X1 U4166 ( .A1(n17902), .A2(n14666), .B1(n17907), .B2(n16845), .ZN(
        n9705) );
  OAI22_X1 U4167 ( .A1(n17836), .A2(n14481), .B1(n17841), .B2(n16851), .ZN(
        n9774) );
  OAI22_X1 U4168 ( .A1(n17858), .A2(n15120), .B1(n17863), .B2(n16851), .ZN(
        n9775) );
  OAI22_X1 U4169 ( .A1(n17880), .A2(n15658), .B1(n17885), .B2(n16851), .ZN(
        n9776) );
  OAI22_X1 U4170 ( .A1(n17902), .A2(n14667), .B1(n17906), .B2(n16851), .ZN(
        n9777) );
  OAI22_X1 U4171 ( .A1(n17836), .A2(n14482), .B1(n17841), .B2(n16857), .ZN(
        n9846) );
  OAI22_X1 U4172 ( .A1(n17858), .A2(n15121), .B1(n17862), .B2(n16857), .ZN(
        n9847) );
  OAI22_X1 U4173 ( .A1(n17880), .A2(n15659), .B1(n17884), .B2(n16857), .ZN(
        n9848) );
  OAI22_X1 U4174 ( .A1(n17902), .A2(n14668), .B1(n17906), .B2(n16857), .ZN(
        n9849) );
  OAI22_X1 U4175 ( .A1(n17858), .A2(n15122), .B1(n17862), .B2(n17512), .ZN(
        n9919) );
  OAI22_X1 U4176 ( .A1(n17880), .A2(n15660), .B1(n17884), .B2(n17512), .ZN(
        n9920) );
  OAI22_X1 U4177 ( .A1(n17944), .A2(n14910), .B1(n17960), .B2(n16436), .ZN(
        n7767) );
  OAI22_X1 U4178 ( .A1(n17967), .A2(n15243), .B1(n17981), .B2(n16442), .ZN(
        n7842) );
  OAI22_X1 U4179 ( .A1(n17925), .A2(n15434), .B1(n17939), .B2(n16448), .ZN(
        n7916) );
  OAI22_X1 U4180 ( .A1(n17858), .A2(n15123), .B1(n17874), .B2(n16436), .ZN(
        n7765) );
  OAI22_X1 U4181 ( .A1(n17902), .A2(n14669), .B1(n17918), .B2(n16436), .ZN(
        n7766) );
  OAI22_X1 U4182 ( .A1(n17882), .A2(n15661), .B1(n17896), .B2(n16442), .ZN(
        n7840) );
  OAI22_X1 U4183 ( .A1(n17838), .A2(n14510), .B1(n17852), .B2(n16731), .ZN(
        n8334) );
  OAI22_X1 U4184 ( .A1(n16692), .A2(n18027), .B1(n16693), .B2(n14860), .ZN(
        n8107) );
  OAI22_X1 U4185 ( .A1(n16692), .A2(n16702), .B1(n16693), .B2(n14051), .ZN(
        n8109) );
  OAI22_X1 U4186 ( .A1(n17577), .A2(n18027), .B1(n17578), .B2(n14052), .ZN(
        n9985) );
  OAI22_X1 U4187 ( .A1(n18003), .A2(n18026), .B1(n18005), .B2(n12048), .ZN(
        n9998) );
  OAI22_X1 U4188 ( .A1(n18016), .A2(n18026), .B1(n18018), .B2(n14534), .ZN(
        n9999) );
  OAI22_X1 U4189 ( .A1(n16934), .A2(n18031), .B1(n14279), .B2(n16936), .ZN(
        n10006) );
  OAI22_X1 U4190 ( .A1(n17017), .A2(n18030), .B1(n14871), .B2(n4420), .ZN(
        n10013) );
  OAI22_X1 U4191 ( .A1(n17036), .A2(n18030), .B1(n14869), .B2(n17038), .ZN(
        n10015) );
  OAI22_X1 U4192 ( .A1(n17049), .A2(n18030), .B1(n14056), .B2(n17051), .ZN(
        n10016) );
  OAI22_X1 U4193 ( .A1(n17577), .A2(n16701), .B1(n17578), .B2(n14856), .ZN(
        n10057) );
  OAI22_X1 U4194 ( .A1(n17281), .A2(n18029), .B1(n14057), .B2(n17283), .ZN(
        n10035) );
  OAI22_X1 U4195 ( .A1(n17294), .A2(n18028), .B1(n14299), .B2(n17296), .ZN(
        n10036) );
  OAI22_X1 U4196 ( .A1(n17346), .A2(n18028), .B1(n14870), .B2(n17348), .ZN(
        n10040) );
  OAI22_X1 U4197 ( .A1(n17372), .A2(n18028), .B1(n14060), .B2(n17374), .ZN(
        n10042) );
  OAI22_X1 U4198 ( .A1(n17398), .A2(n18028), .B1(n14055), .B2(n17400), .ZN(
        n10044) );
  OAI22_X1 U4199 ( .A1(n18004), .A2(n16702), .B1(n18005), .B2(n12049), .ZN(
        n10070) );
  OAI22_X1 U4200 ( .A1(n18017), .A2(n16702), .B1(n18018), .B2(n14535), .ZN(
        n10071) );
  OAI22_X1 U4201 ( .A1(n16877), .A2(n14938), .B1(n16884), .B2(n16436), .ZN(
        n7770) );
  OAI22_X1 U4202 ( .A1(n16920), .A2(n15552), .B1(n16927), .B2(n16436), .ZN(
        n7772) );
  OAI22_X1 U4203 ( .A1(n16945), .A2(n11951), .B1(n16952), .B2(n16437), .ZN(
        n7773) );
  OAI22_X1 U4204 ( .A1(n16966), .A2(n15466), .B1(n16973), .B2(n16437), .ZN(
        n7774) );
  OAI22_X1 U4205 ( .A1(n17009), .A2(n15073), .B1(n17016), .B2(n16437), .ZN(
        n7776) );
  OAI22_X1 U4206 ( .A1(n17137), .A2(n14678), .B1(n17144), .B2(n16437), .ZN(
        n7781) );
  OAI22_X1 U4207 ( .A1(n17160), .A2(n15004), .B1(n17167), .B2(n16437), .ZN(
        n7782) );
  OAI22_X1 U4208 ( .A1(n17182), .A2(n12356), .B1(n17189), .B2(n16437), .ZN(
        n7783) );
  OAI22_X1 U4209 ( .A1(n17202), .A2(n15181), .B1(n17209), .B2(n16437), .ZN(
        n7784) );
  OAI22_X1 U4210 ( .A1(n16877), .A2(n14939), .B1(n16884), .B2(n16442), .ZN(
        n7845) );
  OAI22_X1 U4211 ( .A1(n16910), .A2(n14485), .B1(n16917), .B2(n16442), .ZN(
        n7846) );
  OAI22_X1 U4212 ( .A1(n16920), .A2(n15553), .B1(n16927), .B2(n16442), .ZN(
        n7847) );
  OAI22_X1 U4213 ( .A1(n16956), .A2(n14774), .B1(n16963), .B2(n16443), .ZN(
        n7848) );
  OAI22_X1 U4214 ( .A1(n16966), .A2(n15467), .B1(n16973), .B2(n16443), .ZN(
        n7849) );
  OAI22_X1 U4215 ( .A1(n16999), .A2(n14429), .B1(n17006), .B2(n16443), .ZN(
        n7850) );
  OAI22_X1 U4216 ( .A1(n17009), .A2(n15075), .B1(n17016), .B2(n16443), .ZN(
        n7851) );
  OAI22_X1 U4217 ( .A1(n17160), .A2(n15005), .B1(n17167), .B2(n16443), .ZN(
        n7857) );
  OAI22_X1 U4218 ( .A1(n17192), .A2(n14301), .B1(n17199), .B2(n16443), .ZN(
        n7858) );
  OAI22_X1 U4219 ( .A1(n17202), .A2(n15182), .B1(n17209), .B2(n16443), .ZN(
        n7859) );
  OAI22_X1 U4220 ( .A1(n16887), .A2(n15401), .B1(n16894), .B2(n16448), .ZN(
        n7920) );
  OAI22_X1 U4221 ( .A1(n16910), .A2(n14486), .B1(n16917), .B2(n16448), .ZN(
        n7922) );
  OAI22_X1 U4222 ( .A1(n16920), .A2(n15554), .B1(n16927), .B2(n16448), .ZN(
        n7923) );
  OAI22_X1 U4223 ( .A1(n16976), .A2(n14890), .B1(n16983), .B2(n16449), .ZN(
        n7924) );
  OAI22_X1 U4224 ( .A1(n16999), .A2(n14431), .B1(n17006), .B2(n16449), .ZN(
        n7926) );
  OAI22_X1 U4225 ( .A1(n17009), .A2(n15077), .B1(n17016), .B2(n16449), .ZN(
        n7927) );
  OAI22_X1 U4226 ( .A1(n17171), .A2(n12020), .B1(n17178), .B2(n16449), .ZN(
        n7932) );
  OAI22_X1 U4227 ( .A1(n17182), .A2(n12360), .B1(n17189), .B2(n16449), .ZN(
        n7933) );
  OAI22_X1 U4228 ( .A1(n17192), .A2(n14302), .B1(n17199), .B2(n16449), .ZN(
        n7934) );
  OAI22_X1 U4229 ( .A1(n17202), .A2(n15183), .B1(n17209), .B2(n16449), .ZN(
        n7935) );
  OAI22_X1 U4230 ( .A1(n16877), .A2(n14941), .B1(n16884), .B2(n16456), .ZN(
        n7993) );
  OAI22_X1 U4231 ( .A1(n16887), .A2(n15402), .B1(n16894), .B2(n16457), .ZN(
        n7994) );
  OAI22_X1 U4232 ( .A1(n16910), .A2(n14487), .B1(n16917), .B2(n16457), .ZN(
        n7996) );
  OAI22_X1 U4233 ( .A1(n16920), .A2(n15555), .B1(n16927), .B2(n16457), .ZN(
        n7997) );
  OAI22_X1 U4234 ( .A1(n16944), .A2(n11997), .B1(n16952), .B2(n16709), .ZN(
        n8119) );
  OAI22_X1 U4235 ( .A1(n16956), .A2(n14779), .B1(n16963), .B2(n16709), .ZN(
        n8120) );
  OAI22_X1 U4236 ( .A1(n16966), .A2(n15469), .B1(n16973), .B2(n16709), .ZN(
        n8121) );
  OAI22_X1 U4237 ( .A1(n16976), .A2(n14891), .B1(n16983), .B2(n16710), .ZN(
        n8122) );
  OAI22_X1 U4238 ( .A1(n16999), .A2(n14433), .B1(n17006), .B2(n16710), .ZN(
        n8124) );
  OAI22_X1 U4239 ( .A1(n17009), .A2(n15079), .B1(n17016), .B2(n16710), .ZN(
        n8125) );
  OAI22_X1 U4240 ( .A1(n17137), .A2(n14681), .B1(n17144), .B2(n16718), .ZN(
        n8199) );
  OAI22_X1 U4241 ( .A1(n17160), .A2(n15007), .B1(n17167), .B2(n16718), .ZN(
        n8201) );
  OAI22_X1 U4242 ( .A1(n17170), .A2(n12021), .B1(n17178), .B2(n16719), .ZN(
        n8202) );
  OAI22_X1 U4243 ( .A1(n17182), .A2(n12364), .B1(n17189), .B2(n16719), .ZN(
        n8203) );
  OAI22_X1 U4244 ( .A1(n17192), .A2(n14303), .B1(n17199), .B2(n16719), .ZN(
        n8204) );
  OAI22_X1 U4245 ( .A1(n17202), .A2(n15184), .B1(n17209), .B2(n16719), .ZN(
        n8205) );
  OAI22_X1 U4246 ( .A1(n17062), .A2(n18030), .B1(n14872), .B2(n17064), .ZN(
        n10017) );
  OAI22_X1 U4247 ( .A1(n17210), .A2(n18029), .B1(n14873), .B2(n4362), .ZN(
        n10029) );
  OAI22_X1 U4248 ( .A1(n17411), .A2(n18028), .B1(n14874), .B2(n17413), .ZN(
        n10045) );
  OAI22_X1 U4249 ( .A1(n16877), .A2(n14942), .B1(n16884), .B2(n16725), .ZN(
        n8273) );
  OAI22_X1 U4250 ( .A1(n16887), .A2(n15403), .B1(n16894), .B2(n16726), .ZN(
        n8274) );
  OAI22_X1 U4251 ( .A1(n16910), .A2(n14488), .B1(n16917), .B2(n16726), .ZN(
        n8276) );
  OAI22_X1 U4252 ( .A1(n4448), .A2(n15556), .B1(n16926), .B2(n16726), .ZN(
        n8277) );
  OAI22_X1 U4253 ( .A1(n16945), .A2(n11998), .B1(n16952), .B2(n16726), .ZN(
        n8279) );
  OAI22_X1 U4254 ( .A1(n16956), .A2(n14782), .B1(n16963), .B2(n16726), .ZN(
        n8280) );
  OAI22_X1 U4255 ( .A1(n4432), .A2(n15470), .B1(n16973), .B2(n16726), .ZN(
        n8281) );
  OAI22_X1 U4256 ( .A1(n16976), .A2(n14892), .B1(n16983), .B2(n16726), .ZN(
        n8282) );
  OAI22_X1 U4257 ( .A1(n4423), .A2(n14436), .B1(n17006), .B2(n16726), .ZN(
        n8284) );
  OAI22_X1 U4258 ( .A1(n17009), .A2(n15082), .B1(n17015), .B2(n16726), .ZN(
        n8285) );
  OAI22_X1 U4259 ( .A1(n17137), .A2(n14682), .B1(n17144), .B2(n16727), .ZN(
        n8295) );
  OAI22_X1 U4260 ( .A1(n17160), .A2(n15008), .B1(n17167), .B2(n16727), .ZN(
        n8297) );
  OAI22_X1 U4261 ( .A1(n17171), .A2(n12022), .B1(n17178), .B2(n16728), .ZN(
        n8298) );
  OAI22_X1 U4262 ( .A1(n17182), .A2(n12366), .B1(n17189), .B2(n16728), .ZN(
        n8299) );
  OAI22_X1 U4263 ( .A1(n17192), .A2(n14304), .B1(n17199), .B2(n16728), .ZN(
        n8300) );
  OAI22_X1 U4264 ( .A1(n17202), .A2(n15185), .B1(n17208), .B2(n16728), .ZN(
        n8301) );
  OAI22_X1 U4265 ( .A1(n16877), .A2(n14943), .B1(n16883), .B2(n16732), .ZN(
        n8345) );
  OAI22_X1 U4266 ( .A1(n16887), .A2(n15404), .B1(n16894), .B2(n16732), .ZN(
        n8346) );
  OAI22_X1 U4267 ( .A1(n16910), .A2(n14489), .B1(n16916), .B2(n16732), .ZN(
        n8348) );
  OAI22_X1 U4268 ( .A1(n4448), .A2(n15557), .B1(n16926), .B2(n16732), .ZN(
        n8349) );
  OAI22_X1 U4269 ( .A1(n16945), .A2(n11999), .B1(n16952), .B2(n16733), .ZN(
        n8351) );
  OAI22_X1 U4270 ( .A1(n16956), .A2(n14784), .B1(n16963), .B2(n16733), .ZN(
        n8352) );
  OAI22_X1 U4271 ( .A1(n4432), .A2(n15471), .B1(n16972), .B2(n16733), .ZN(
        n8353) );
  OAI22_X1 U4272 ( .A1(n16976), .A2(n14893), .B1(n16983), .B2(n16733), .ZN(
        n8354) );
  OAI22_X1 U4273 ( .A1(n4423), .A2(n14438), .B1(n17005), .B2(n16733), .ZN(
        n8356) );
  OAI22_X1 U4274 ( .A1(n17009), .A2(n15084), .B1(n17015), .B2(n16733), .ZN(
        n8357) );
  OAI22_X1 U4275 ( .A1(n17137), .A2(n14683), .B1(n17144), .B2(n16734), .ZN(
        n8367) );
  OAI22_X1 U4276 ( .A1(n17160), .A2(n15009), .B1(n17166), .B2(n16734), .ZN(
        n8369) );
  OAI22_X1 U4277 ( .A1(n17171), .A2(n12023), .B1(n17178), .B2(n16734), .ZN(
        n8370) );
  OAI22_X1 U4278 ( .A1(n17182), .A2(n12368), .B1(n17188), .B2(n16734), .ZN(
        n8371) );
  OAI22_X1 U4279 ( .A1(n17192), .A2(n14305), .B1(n17198), .B2(n16734), .ZN(
        n8372) );
  OAI22_X1 U4280 ( .A1(n17202), .A2(n15186), .B1(n17208), .B2(n16734), .ZN(
        n8373) );
  OAI22_X1 U4281 ( .A1(n16877), .A2(n14944), .B1(n16883), .B2(n16738), .ZN(
        n8417) );
  OAI22_X1 U4282 ( .A1(n16887), .A2(n15405), .B1(n16893), .B2(n16738), .ZN(
        n8418) );
  OAI22_X1 U4283 ( .A1(n16910), .A2(n14490), .B1(n16916), .B2(n16738), .ZN(
        n8420) );
  OAI22_X1 U4284 ( .A1(n4448), .A2(n15558), .B1(n16926), .B2(n16738), .ZN(
        n8421) );
  OAI22_X1 U4285 ( .A1(n16945), .A2(n12000), .B1(n16951), .B2(n16739), .ZN(
        n8423) );
  OAI22_X1 U4286 ( .A1(n16956), .A2(n14786), .B1(n16962), .B2(n16739), .ZN(
        n8424) );
  OAI22_X1 U4287 ( .A1(n4432), .A2(n15472), .B1(n16972), .B2(n16739), .ZN(
        n8425) );
  OAI22_X1 U4288 ( .A1(n16976), .A2(n14894), .B1(n16982), .B2(n16739), .ZN(
        n8426) );
  OAI22_X1 U4289 ( .A1(n4423), .A2(n14440), .B1(n17005), .B2(n16739), .ZN(
        n8428) );
  OAI22_X1 U4290 ( .A1(n17009), .A2(n15086), .B1(n17015), .B2(n16739), .ZN(
        n8429) );
  OAI22_X1 U4291 ( .A1(n17137), .A2(n14684), .B1(n17143), .B2(n16740), .ZN(
        n8439) );
  OAI22_X1 U4292 ( .A1(n17160), .A2(n15010), .B1(n17166), .B2(n16740), .ZN(
        n8441) );
  OAI22_X1 U4293 ( .A1(n17171), .A2(n12024), .B1(n17177), .B2(n16740), .ZN(
        n8442) );
  OAI22_X1 U4294 ( .A1(n17182), .A2(n12407), .B1(n17188), .B2(n16740), .ZN(
        n8443) );
  OAI22_X1 U4295 ( .A1(n17192), .A2(n14306), .B1(n17198), .B2(n16740), .ZN(
        n8444) );
  OAI22_X1 U4296 ( .A1(n17202), .A2(n15187), .B1(n17208), .B2(n16740), .ZN(
        n8445) );
  OAI22_X1 U4297 ( .A1(n16877), .A2(n14945), .B1(n16883), .B2(n16744), .ZN(
        n8489) );
  OAI22_X1 U4298 ( .A1(n16887), .A2(n15406), .B1(n16893), .B2(n16744), .ZN(
        n8490) );
  OAI22_X1 U4299 ( .A1(n16910), .A2(n14491), .B1(n16916), .B2(n16744), .ZN(
        n8492) );
  OAI22_X1 U4300 ( .A1(n4448), .A2(n15559), .B1(n16926), .B2(n16744), .ZN(
        n8493) );
  OAI22_X1 U4301 ( .A1(n16945), .A2(n12001), .B1(n16951), .B2(n16745), .ZN(
        n8495) );
  OAI22_X1 U4302 ( .A1(n16956), .A2(n14788), .B1(n16962), .B2(n16745), .ZN(
        n8496) );
  OAI22_X1 U4303 ( .A1(n4432), .A2(n15473), .B1(n16972), .B2(n16745), .ZN(
        n8497) );
  OAI22_X1 U4304 ( .A1(n16976), .A2(n14895), .B1(n16982), .B2(n16745), .ZN(
        n8498) );
  OAI22_X1 U4305 ( .A1(n4423), .A2(n14442), .B1(n17005), .B2(n16745), .ZN(
        n8500) );
  OAI22_X1 U4306 ( .A1(n17009), .A2(n15088), .B1(n17015), .B2(n16745), .ZN(
        n8501) );
  OAI22_X1 U4307 ( .A1(n17137), .A2(n14685), .B1(n17143), .B2(n16746), .ZN(
        n8511) );
  OAI22_X1 U4308 ( .A1(n17160), .A2(n15011), .B1(n17166), .B2(n16746), .ZN(
        n8513) );
  OAI22_X1 U4309 ( .A1(n17171), .A2(n12025), .B1(n17177), .B2(n16746), .ZN(
        n8514) );
  OAI22_X1 U4310 ( .A1(n17182), .A2(n12409), .B1(n17188), .B2(n16746), .ZN(
        n8515) );
  OAI22_X1 U4311 ( .A1(n17192), .A2(n14307), .B1(n17198), .B2(n16746), .ZN(
        n8516) );
  OAI22_X1 U4312 ( .A1(n17202), .A2(n15188), .B1(n17208), .B2(n16746), .ZN(
        n8517) );
  OAI22_X1 U4313 ( .A1(n16877), .A2(n14946), .B1(n16883), .B2(n16750), .ZN(
        n8561) );
  OAI22_X1 U4314 ( .A1(n16887), .A2(n15407), .B1(n16893), .B2(n16750), .ZN(
        n8562) );
  OAI22_X1 U4315 ( .A1(n16910), .A2(n14492), .B1(n16916), .B2(n16750), .ZN(
        n8564) );
  OAI22_X1 U4316 ( .A1(n4448), .A2(n15560), .B1(n16925), .B2(n16750), .ZN(
        n8565) );
  OAI22_X1 U4317 ( .A1(n16945), .A2(n12002), .B1(n16951), .B2(n16751), .ZN(
        n8567) );
  OAI22_X1 U4318 ( .A1(n16956), .A2(n14790), .B1(n16962), .B2(n16751), .ZN(
        n8568) );
  OAI22_X1 U4319 ( .A1(n4432), .A2(n15474), .B1(n16972), .B2(n16751), .ZN(
        n8569) );
  OAI22_X1 U4320 ( .A1(n16976), .A2(n14896), .B1(n16982), .B2(n16751), .ZN(
        n8570) );
  OAI22_X1 U4321 ( .A1(n4423), .A2(n14444), .B1(n17005), .B2(n16751), .ZN(
        n8572) );
  OAI22_X1 U4322 ( .A1(n17009), .A2(n15090), .B1(n17014), .B2(n16751), .ZN(
        n8573) );
  OAI22_X1 U4323 ( .A1(n17137), .A2(n14686), .B1(n17143), .B2(n16752), .ZN(
        n8583) );
  OAI22_X1 U4324 ( .A1(n17160), .A2(n15012), .B1(n17166), .B2(n16752), .ZN(
        n8585) );
  OAI22_X1 U4325 ( .A1(n17171), .A2(n12026), .B1(n17177), .B2(n16752), .ZN(
        n8586) );
  OAI22_X1 U4326 ( .A1(n17182), .A2(n12411), .B1(n17188), .B2(n16752), .ZN(
        n8587) );
  OAI22_X1 U4327 ( .A1(n17192), .A2(n14308), .B1(n17198), .B2(n16752), .ZN(
        n8588) );
  OAI22_X1 U4328 ( .A1(n17202), .A2(n15189), .B1(n17207), .B2(n16752), .ZN(
        n8589) );
  OAI22_X1 U4329 ( .A1(n16877), .A2(n14947), .B1(n16882), .B2(n16756), .ZN(
        n8633) );
  OAI22_X1 U4330 ( .A1(n16887), .A2(n15408), .B1(n16893), .B2(n16756), .ZN(
        n8634) );
  OAI22_X1 U4331 ( .A1(n16910), .A2(n14493), .B1(n16915), .B2(n16756), .ZN(
        n8636) );
  OAI22_X1 U4332 ( .A1(n4448), .A2(n15561), .B1(n16925), .B2(n16756), .ZN(
        n8637) );
  OAI22_X1 U4333 ( .A1(n16945), .A2(n12003), .B1(n16951), .B2(n16757), .ZN(
        n8639) );
  OAI22_X1 U4334 ( .A1(n16956), .A2(n14792), .B1(n16962), .B2(n16757), .ZN(
        n8640) );
  OAI22_X1 U4335 ( .A1(n4432), .A2(n15475), .B1(n16971), .B2(n16757), .ZN(
        n8641) );
  OAI22_X1 U4336 ( .A1(n16976), .A2(n14897), .B1(n16982), .B2(n16757), .ZN(
        n8642) );
  OAI22_X1 U4337 ( .A1(n4423), .A2(n14446), .B1(n17004), .B2(n16757), .ZN(
        n8644) );
  OAI22_X1 U4338 ( .A1(n17009), .A2(n15092), .B1(n17014), .B2(n16757), .ZN(
        n8645) );
  OAI22_X1 U4339 ( .A1(n17137), .A2(n14687), .B1(n17143), .B2(n16758), .ZN(
        n8655) );
  OAI22_X1 U4340 ( .A1(n17160), .A2(n15013), .B1(n17165), .B2(n16758), .ZN(
        n8657) );
  OAI22_X1 U4341 ( .A1(n17171), .A2(n12027), .B1(n17177), .B2(n16758), .ZN(
        n8658) );
  OAI22_X1 U4342 ( .A1(n17182), .A2(n12600), .B1(n17187), .B2(n16758), .ZN(
        n8659) );
  OAI22_X1 U4343 ( .A1(n17192), .A2(n14309), .B1(n17197), .B2(n16758), .ZN(
        n8660) );
  OAI22_X1 U4344 ( .A1(n17202), .A2(n15190), .B1(n17207), .B2(n16758), .ZN(
        n8661) );
  OAI22_X1 U4345 ( .A1(n16877), .A2(n14948), .B1(n16882), .B2(n16762), .ZN(
        n8705) );
  OAI22_X1 U4346 ( .A1(n16887), .A2(n15409), .B1(n16892), .B2(n16762), .ZN(
        n8706) );
  OAI22_X1 U4347 ( .A1(n16910), .A2(n14494), .B1(n16915), .B2(n16762), .ZN(
        n8708) );
  OAI22_X1 U4348 ( .A1(n4448), .A2(n15562), .B1(n16925), .B2(n16762), .ZN(
        n8709) );
  OAI22_X1 U4349 ( .A1(n16945), .A2(n12004), .B1(n16950), .B2(n16763), .ZN(
        n8711) );
  OAI22_X1 U4350 ( .A1(n16956), .A2(n14794), .B1(n16961), .B2(n16763), .ZN(
        n8712) );
  OAI22_X1 U4351 ( .A1(n4432), .A2(n15476), .B1(n16971), .B2(n16763), .ZN(
        n8713) );
  OAI22_X1 U4352 ( .A1(n16976), .A2(n14898), .B1(n16981), .B2(n16763), .ZN(
        n8714) );
  OAI22_X1 U4353 ( .A1(n4423), .A2(n14448), .B1(n17004), .B2(n16763), .ZN(
        n8716) );
  OAI22_X1 U4354 ( .A1(n17009), .A2(n15094), .B1(n17014), .B2(n16763), .ZN(
        n8717) );
  OAI22_X1 U4355 ( .A1(n17137), .A2(n14688), .B1(n17142), .B2(n16764), .ZN(
        n8727) );
  OAI22_X1 U4356 ( .A1(n17160), .A2(n15014), .B1(n17165), .B2(n16764), .ZN(
        n8729) );
  OAI22_X1 U4357 ( .A1(n17171), .A2(n12028), .B1(n17176), .B2(n16764), .ZN(
        n8730) );
  OAI22_X1 U4358 ( .A1(n17182), .A2(n12652), .B1(n17187), .B2(n16764), .ZN(
        n8731) );
  OAI22_X1 U4359 ( .A1(n17192), .A2(n14310), .B1(n17197), .B2(n16764), .ZN(
        n8732) );
  OAI22_X1 U4360 ( .A1(n17202), .A2(n15191), .B1(n17207), .B2(n16764), .ZN(
        n8733) );
  OAI22_X1 U4361 ( .A1(n16877), .A2(n14949), .B1(n16882), .B2(n16768), .ZN(
        n8777) );
  OAI22_X1 U4362 ( .A1(n16887), .A2(n15410), .B1(n16892), .B2(n16768), .ZN(
        n8778) );
  OAI22_X1 U4363 ( .A1(n16910), .A2(n14495), .B1(n16915), .B2(n16768), .ZN(
        n8780) );
  OAI22_X1 U4364 ( .A1(n16920), .A2(n15563), .B1(n16924), .B2(n16768), .ZN(
        n8781) );
  OAI22_X1 U4365 ( .A1(n16945), .A2(n12005), .B1(n16950), .B2(n16769), .ZN(
        n8783) );
  OAI22_X1 U4366 ( .A1(n16956), .A2(n14796), .B1(n16961), .B2(n16769), .ZN(
        n8784) );
  OAI22_X1 U4367 ( .A1(n16966), .A2(n15477), .B1(n16971), .B2(n16769), .ZN(
        n8785) );
  OAI22_X1 U4368 ( .A1(n16976), .A2(n14899), .B1(n16981), .B2(n16769), .ZN(
        n8786) );
  OAI22_X1 U4369 ( .A1(n16999), .A2(n14450), .B1(n17004), .B2(n16769), .ZN(
        n8788) );
  OAI22_X1 U4370 ( .A1(n17009), .A2(n15096), .B1(n17013), .B2(n16769), .ZN(
        n8789) );
  OAI22_X1 U4371 ( .A1(n17137), .A2(n14689), .B1(n17142), .B2(n16770), .ZN(
        n8799) );
  OAI22_X1 U4372 ( .A1(n17160), .A2(n15015), .B1(n17165), .B2(n16770), .ZN(
        n8801) );
  OAI22_X1 U4373 ( .A1(n17171), .A2(n12030), .B1(n17176), .B2(n16770), .ZN(
        n8802) );
  OAI22_X1 U4374 ( .A1(n17182), .A2(n13996), .B1(n17187), .B2(n16770), .ZN(
        n8803) );
  OAI22_X1 U4375 ( .A1(n17192), .A2(n14311), .B1(n17197), .B2(n16770), .ZN(
        n8804) );
  OAI22_X1 U4376 ( .A1(n17202), .A2(n15192), .B1(n17206), .B2(n16770), .ZN(
        n8805) );
  OAI22_X1 U4377 ( .A1(n16877), .A2(n14950), .B1(n16881), .B2(n16774), .ZN(
        n8849) );
  OAI22_X1 U4378 ( .A1(n16887), .A2(n15411), .B1(n16892), .B2(n16774), .ZN(
        n8850) );
  OAI22_X1 U4379 ( .A1(n16910), .A2(n14496), .B1(n16914), .B2(n16774), .ZN(
        n8852) );
  OAI22_X1 U4380 ( .A1(n4448), .A2(n15564), .B1(n16924), .B2(n16774), .ZN(
        n8853) );
  OAI22_X1 U4381 ( .A1(n16945), .A2(n12006), .B1(n16950), .B2(n16775), .ZN(
        n8855) );
  OAI22_X1 U4382 ( .A1(n16956), .A2(n14798), .B1(n16961), .B2(n16775), .ZN(
        n8856) );
  OAI22_X1 U4383 ( .A1(n4432), .A2(n15478), .B1(n16970), .B2(n16775), .ZN(
        n8857) );
  OAI22_X1 U4384 ( .A1(n16976), .A2(n14900), .B1(n16981), .B2(n16775), .ZN(
        n8858) );
  OAI22_X1 U4385 ( .A1(n4423), .A2(n14452), .B1(n17003), .B2(n16775), .ZN(
        n8860) );
  OAI22_X1 U4386 ( .A1(n17009), .A2(n15098), .B1(n17013), .B2(n16775), .ZN(
        n8861) );
  OAI22_X1 U4387 ( .A1(n17137), .A2(n14690), .B1(n17142), .B2(n16776), .ZN(
        n8871) );
  OAI22_X1 U4388 ( .A1(n17160), .A2(n15016), .B1(n17164), .B2(n16776), .ZN(
        n8873) );
  OAI22_X1 U4389 ( .A1(n17171), .A2(n12031), .B1(n17176), .B2(n16776), .ZN(
        n8874) );
  OAI22_X1 U4390 ( .A1(n17182), .A2(n14008), .B1(n17186), .B2(n16776), .ZN(
        n8875) );
  OAI22_X1 U4391 ( .A1(n17192), .A2(n14312), .B1(n17196), .B2(n16776), .ZN(
        n8876) );
  OAI22_X1 U4392 ( .A1(n17202), .A2(n15193), .B1(n17206), .B2(n16776), .ZN(
        n8877) );
  OAI22_X1 U4393 ( .A1(n16877), .A2(n14951), .B1(n16881), .B2(n16780), .ZN(
        n8921) );
  OAI22_X1 U4394 ( .A1(n16887), .A2(n15412), .B1(n16891), .B2(n16780), .ZN(
        n8922) );
  OAI22_X1 U4395 ( .A1(n16910), .A2(n14497), .B1(n16914), .B2(n16780), .ZN(
        n8924) );
  OAI22_X1 U4396 ( .A1(n4448), .A2(n15565), .B1(n16924), .B2(n16780), .ZN(
        n8925) );
  OAI22_X1 U4397 ( .A1(n16945), .A2(n12007), .B1(n16949), .B2(n16781), .ZN(
        n8927) );
  OAI22_X1 U4398 ( .A1(n16956), .A2(n14800), .B1(n16960), .B2(n16781), .ZN(
        n8928) );
  OAI22_X1 U4399 ( .A1(n4432), .A2(n15479), .B1(n16970), .B2(n16781), .ZN(
        n8929) );
  OAI22_X1 U4400 ( .A1(n16976), .A2(n14901), .B1(n16980), .B2(n16781), .ZN(
        n8930) );
  OAI22_X1 U4401 ( .A1(n4423), .A2(n14454), .B1(n17003), .B2(n16781), .ZN(
        n8932) );
  OAI22_X1 U4402 ( .A1(n17009), .A2(n15100), .B1(n17013), .B2(n16781), .ZN(
        n8933) );
  OAI22_X1 U4403 ( .A1(n17137), .A2(n14691), .B1(n17141), .B2(n16782), .ZN(
        n8943) );
  OAI22_X1 U4404 ( .A1(n17160), .A2(n15017), .B1(n17164), .B2(n16782), .ZN(
        n8945) );
  OAI22_X1 U4405 ( .A1(n17171), .A2(n12032), .B1(n17175), .B2(n16782), .ZN(
        n8946) );
  OAI22_X1 U4406 ( .A1(n17182), .A2(n14015), .B1(n17186), .B2(n16782), .ZN(
        n8947) );
  OAI22_X1 U4407 ( .A1(n17192), .A2(n14313), .B1(n17196), .B2(n16782), .ZN(
        n8948) );
  OAI22_X1 U4408 ( .A1(n17202), .A2(n15194), .B1(n17206), .B2(n16782), .ZN(
        n8949) );
  OAI22_X1 U4409 ( .A1(n16877), .A2(n14952), .B1(n16881), .B2(n16786), .ZN(
        n8993) );
  OAI22_X1 U4410 ( .A1(n16887), .A2(n15413), .B1(n16891), .B2(n16786), .ZN(
        n8994) );
  OAI22_X1 U4411 ( .A1(n16910), .A2(n14498), .B1(n16914), .B2(n16786), .ZN(
        n8996) );
  OAI22_X1 U4412 ( .A1(n4448), .A2(n15566), .B1(n16924), .B2(n16786), .ZN(
        n8997) );
  OAI22_X1 U4413 ( .A1(n16945), .A2(n12008), .B1(n16949), .B2(n16787), .ZN(
        n8999) );
  OAI22_X1 U4414 ( .A1(n16956), .A2(n14802), .B1(n16960), .B2(n16787), .ZN(
        n9000) );
  OAI22_X1 U4415 ( .A1(n4432), .A2(n15480), .B1(n16970), .B2(n16787), .ZN(
        n9001) );
  OAI22_X1 U4416 ( .A1(n16976), .A2(n14902), .B1(n16980), .B2(n16787), .ZN(
        n9002) );
  OAI22_X1 U4417 ( .A1(n4423), .A2(n14456), .B1(n17003), .B2(n16787), .ZN(
        n9004) );
  OAI22_X1 U4418 ( .A1(n17009), .A2(n15102), .B1(n17013), .B2(n16787), .ZN(
        n9005) );
  OAI22_X1 U4419 ( .A1(n17137), .A2(n14692), .B1(n17141), .B2(n16788), .ZN(
        n9015) );
  OAI22_X1 U4420 ( .A1(n17160), .A2(n15018), .B1(n17164), .B2(n16788), .ZN(
        n9017) );
  OAI22_X1 U4421 ( .A1(n17171), .A2(n12033), .B1(n17175), .B2(n16788), .ZN(
        n9018) );
  OAI22_X1 U4422 ( .A1(n17182), .A2(n14035), .B1(n17186), .B2(n16788), .ZN(
        n9019) );
  OAI22_X1 U4423 ( .A1(n17192), .A2(n14314), .B1(n17196), .B2(n16788), .ZN(
        n9020) );
  OAI22_X1 U4424 ( .A1(n17202), .A2(n15195), .B1(n17206), .B2(n16788), .ZN(
        n9021) );
  OAI22_X1 U4425 ( .A1(n16877), .A2(n14953), .B1(n16881), .B2(n16792), .ZN(
        n9065) );
  OAI22_X1 U4426 ( .A1(n16887), .A2(n15414), .B1(n16891), .B2(n16792), .ZN(
        n9066) );
  OAI22_X1 U4427 ( .A1(n16910), .A2(n14499), .B1(n16914), .B2(n16792), .ZN(
        n9068) );
  OAI22_X1 U4428 ( .A1(n16920), .A2(n15567), .B1(n16923), .B2(n16792), .ZN(
        n9069) );
  OAI22_X1 U4429 ( .A1(n16945), .A2(n12009), .B1(n16949), .B2(n16793), .ZN(
        n9071) );
  OAI22_X1 U4430 ( .A1(n16956), .A2(n14804), .B1(n16960), .B2(n16793), .ZN(
        n9072) );
  OAI22_X1 U4431 ( .A1(n16966), .A2(n15481), .B1(n16970), .B2(n16793), .ZN(
        n9073) );
  OAI22_X1 U4432 ( .A1(n16976), .A2(n14903), .B1(n16980), .B2(n16793), .ZN(
        n9074) );
  OAI22_X1 U4433 ( .A1(n16999), .A2(n14458), .B1(n17003), .B2(n16793), .ZN(
        n9076) );
  OAI22_X1 U4434 ( .A1(n17009), .A2(n15104), .B1(n17012), .B2(n16793), .ZN(
        n9077) );
  OAI22_X1 U4435 ( .A1(n17137), .A2(n14693), .B1(n17141), .B2(n16794), .ZN(
        n9087) );
  OAI22_X1 U4436 ( .A1(n17160), .A2(n15019), .B1(n17164), .B2(n16794), .ZN(
        n9089) );
  OAI22_X1 U4437 ( .A1(n17171), .A2(n12034), .B1(n17175), .B2(n16794), .ZN(
        n9090) );
  OAI22_X1 U4438 ( .A1(n17182), .A2(n14037), .B1(n17186), .B2(n16794), .ZN(
        n9091) );
  OAI22_X1 U4439 ( .A1(n17192), .A2(n14315), .B1(n17196), .B2(n16794), .ZN(
        n9092) );
  OAI22_X1 U4440 ( .A1(n17202), .A2(n15196), .B1(n17205), .B2(n16794), .ZN(
        n9093) );
  OAI22_X1 U4441 ( .A1(n16877), .A2(n14954), .B1(n16880), .B2(n16798), .ZN(
        n9137) );
  OAI22_X1 U4442 ( .A1(n16887), .A2(n15415), .B1(n16891), .B2(n16798), .ZN(
        n9138) );
  OAI22_X1 U4443 ( .A1(n16910), .A2(n14500), .B1(n16913), .B2(n16798), .ZN(
        n9140) );
  OAI22_X1 U4444 ( .A1(n16920), .A2(n15568), .B1(n16923), .B2(n16798), .ZN(
        n9141) );
  OAI22_X1 U4445 ( .A1(n16945), .A2(n12010), .B1(n16949), .B2(n16799), .ZN(
        n9143) );
  OAI22_X1 U4446 ( .A1(n16956), .A2(n14806), .B1(n16960), .B2(n16799), .ZN(
        n9144) );
  OAI22_X1 U4447 ( .A1(n16966), .A2(n15482), .B1(n16969), .B2(n16799), .ZN(
        n9145) );
  OAI22_X1 U4448 ( .A1(n16976), .A2(n14904), .B1(n16980), .B2(n16799), .ZN(
        n9146) );
  OAI22_X1 U4449 ( .A1(n16999), .A2(n14460), .B1(n17002), .B2(n16799), .ZN(
        n9148) );
  OAI22_X1 U4450 ( .A1(n17009), .A2(n15106), .B1(n17012), .B2(n16799), .ZN(
        n9149) );
  OAI22_X1 U4451 ( .A1(n17137), .A2(n14694), .B1(n17141), .B2(n16800), .ZN(
        n9159) );
  OAI22_X1 U4452 ( .A1(n17160), .A2(n15020), .B1(n17163), .B2(n16800), .ZN(
        n9161) );
  OAI22_X1 U4453 ( .A1(n17171), .A2(n12035), .B1(n17175), .B2(n16800), .ZN(
        n9162) );
  OAI22_X1 U4454 ( .A1(n17182), .A2(n14039), .B1(n17185), .B2(n16800), .ZN(
        n9163) );
  OAI22_X1 U4455 ( .A1(n17192), .A2(n14316), .B1(n17195), .B2(n16800), .ZN(
        n9164) );
  OAI22_X1 U4456 ( .A1(n17202), .A2(n15197), .B1(n17205), .B2(n16800), .ZN(
        n9165) );
  OAI22_X1 U4457 ( .A1(n16877), .A2(n14955), .B1(n16880), .B2(n16804), .ZN(
        n9209) );
  OAI22_X1 U4458 ( .A1(n16887), .A2(n15416), .B1(n16890), .B2(n16804), .ZN(
        n9210) );
  OAI22_X1 U4459 ( .A1(n16910), .A2(n14501), .B1(n16913), .B2(n16804), .ZN(
        n9212) );
  OAI22_X1 U4460 ( .A1(n4448), .A2(n15569), .B1(n16923), .B2(n16804), .ZN(
        n9213) );
  OAI22_X1 U4461 ( .A1(n16945), .A2(n12011), .B1(n16948), .B2(n16805), .ZN(
        n9215) );
  OAI22_X1 U4462 ( .A1(n16956), .A2(n14808), .B1(n16959), .B2(n16805), .ZN(
        n9216) );
  OAI22_X1 U4463 ( .A1(n4432), .A2(n15483), .B1(n16969), .B2(n16805), .ZN(
        n9217) );
  OAI22_X1 U4464 ( .A1(n16976), .A2(n14905), .B1(n16979), .B2(n16805), .ZN(
        n9218) );
  OAI22_X1 U4465 ( .A1(n4423), .A2(n14462), .B1(n17002), .B2(n16805), .ZN(
        n9220) );
  OAI22_X1 U4466 ( .A1(n17009), .A2(n15108), .B1(n17012), .B2(n16805), .ZN(
        n9221) );
  OAI22_X1 U4467 ( .A1(n17137), .A2(n14695), .B1(n17140), .B2(n16806), .ZN(
        n9231) );
  OAI22_X1 U4468 ( .A1(n17160), .A2(n15021), .B1(n17163), .B2(n16806), .ZN(
        n9233) );
  OAI22_X1 U4469 ( .A1(n17171), .A2(n12036), .B1(n17174), .B2(n16806), .ZN(
        n9234) );
  OAI22_X1 U4470 ( .A1(n17182), .A2(n14041), .B1(n17185), .B2(n16806), .ZN(
        n9235) );
  OAI22_X1 U4471 ( .A1(n17192), .A2(n14317), .B1(n17195), .B2(n16806), .ZN(
        n9236) );
  OAI22_X1 U4472 ( .A1(n17202), .A2(n15198), .B1(n17205), .B2(n16806), .ZN(
        n9237) );
  OAI22_X1 U4473 ( .A1(n4462), .A2(n14956), .B1(n16880), .B2(n16810), .ZN(
        n9281) );
  OAI22_X1 U4474 ( .A1(n4459), .A2(n15417), .B1(n16890), .B2(n16810), .ZN(
        n9282) );
  OAI22_X1 U4475 ( .A1(n4451), .A2(n14502), .B1(n16913), .B2(n16810), .ZN(
        n9284) );
  OAI22_X1 U4476 ( .A1(n16920), .A2(n15570), .B1(n16923), .B2(n16810), .ZN(
        n9285) );
  OAI22_X1 U4477 ( .A1(n4438), .A2(n12012), .B1(n16948), .B2(n16811), .ZN(
        n9287) );
  OAI22_X1 U4478 ( .A1(n4435), .A2(n14810), .B1(n16959), .B2(n16811), .ZN(
        n9288) );
  OAI22_X1 U4479 ( .A1(n16966), .A2(n15484), .B1(n16969), .B2(n16811), .ZN(
        n9289) );
  OAI22_X1 U4480 ( .A1(n4429), .A2(n14906), .B1(n16979), .B2(n16811), .ZN(
        n9290) );
  OAI22_X1 U4481 ( .A1(n16999), .A2(n14464), .B1(n17002), .B2(n16811), .ZN(
        n9292) );
  OAI22_X1 U4482 ( .A1(n4420), .A2(n15110), .B1(n17012), .B2(n16811), .ZN(
        n9293) );
  OAI22_X1 U4483 ( .A1(n4382), .A2(n14696), .B1(n17140), .B2(n16812), .ZN(
        n9303) );
  OAI22_X1 U4484 ( .A1(n4376), .A2(n15022), .B1(n17163), .B2(n16812), .ZN(
        n9305) );
  OAI22_X1 U4485 ( .A1(n4373), .A2(n12037), .B1(n17174), .B2(n16812), .ZN(
        n9306) );
  OAI22_X1 U4486 ( .A1(n4370), .A2(n14043), .B1(n17185), .B2(n16812), .ZN(
        n9307) );
  OAI22_X1 U4487 ( .A1(n4367), .A2(n14318), .B1(n17195), .B2(n16812), .ZN(
        n9308) );
  OAI22_X1 U4488 ( .A1(n4362), .A2(n15199), .B1(n17205), .B2(n16812), .ZN(
        n9309) );
  OAI22_X1 U4489 ( .A1(n4462), .A2(n14957), .B1(n16880), .B2(n16816), .ZN(
        n9353) );
  OAI22_X1 U4490 ( .A1(n4459), .A2(n15418), .B1(n16890), .B2(n16816), .ZN(
        n9354) );
  OAI22_X1 U4491 ( .A1(n4451), .A2(n14503), .B1(n16913), .B2(n16816), .ZN(
        n9356) );
  OAI22_X1 U4492 ( .A1(n16920), .A2(n15571), .B1(n16922), .B2(n16816), .ZN(
        n9357) );
  OAI22_X1 U4493 ( .A1(n4438), .A2(n12013), .B1(n16948), .B2(n16817), .ZN(
        n9359) );
  OAI22_X1 U4494 ( .A1(n4435), .A2(n14812), .B1(n16959), .B2(n16817), .ZN(
        n9360) );
  OAI22_X1 U4495 ( .A1(n16966), .A2(n15485), .B1(n16969), .B2(n16817), .ZN(
        n9361) );
  OAI22_X1 U4496 ( .A1(n4429), .A2(n14907), .B1(n16979), .B2(n16817), .ZN(
        n9362) );
  OAI22_X1 U4497 ( .A1(n16999), .A2(n14466), .B1(n17002), .B2(n16817), .ZN(
        n9364) );
  OAI22_X1 U4498 ( .A1(n4420), .A2(n15112), .B1(n17011), .B2(n16817), .ZN(
        n9365) );
  OAI22_X1 U4499 ( .A1(n4382), .A2(n14697), .B1(n17140), .B2(n16818), .ZN(
        n9375) );
  OAI22_X1 U4500 ( .A1(n4376), .A2(n15023), .B1(n17163), .B2(n16818), .ZN(
        n9377) );
  OAI22_X1 U4501 ( .A1(n4373), .A2(n12038), .B1(n17174), .B2(n16818), .ZN(
        n9378) );
  OAI22_X1 U4502 ( .A1(n4370), .A2(n14045), .B1(n17185), .B2(n16818), .ZN(
        n9379) );
  OAI22_X1 U4503 ( .A1(n4367), .A2(n14319), .B1(n17195), .B2(n16818), .ZN(
        n9380) );
  OAI22_X1 U4504 ( .A1(n4362), .A2(n15200), .B1(n17204), .B2(n16818), .ZN(
        n9381) );
  OAI22_X1 U4505 ( .A1(n4462), .A2(n14958), .B1(n16879), .B2(n16822), .ZN(
        n9425) );
  OAI22_X1 U4506 ( .A1(n4459), .A2(n15419), .B1(n16890), .B2(n16822), .ZN(
        n9426) );
  OAI22_X1 U4507 ( .A1(n4451), .A2(n14504), .B1(n16912), .B2(n16822), .ZN(
        n9428) );
  OAI22_X1 U4508 ( .A1(n16920), .A2(n15572), .B1(n16922), .B2(n16822), .ZN(
        n9429) );
  OAI22_X1 U4509 ( .A1(n4438), .A2(n12014), .B1(n16948), .B2(n16823), .ZN(
        n9431) );
  OAI22_X1 U4510 ( .A1(n4435), .A2(n14814), .B1(n16959), .B2(n16823), .ZN(
        n9432) );
  OAI22_X1 U4511 ( .A1(n16966), .A2(n15486), .B1(n16968), .B2(n16823), .ZN(
        n9433) );
  OAI22_X1 U4512 ( .A1(n4429), .A2(n14908), .B1(n16979), .B2(n16823), .ZN(
        n9434) );
  OAI22_X1 U4513 ( .A1(n16999), .A2(n14468), .B1(n17001), .B2(n16823), .ZN(
        n9436) );
  OAI22_X1 U4514 ( .A1(n4420), .A2(n15114), .B1(n17011), .B2(n16823), .ZN(
        n9437) );
  OAI22_X1 U4515 ( .A1(n4382), .A2(n14698), .B1(n17140), .B2(n16824), .ZN(
        n9447) );
  OAI22_X1 U4516 ( .A1(n4376), .A2(n15024), .B1(n17162), .B2(n16824), .ZN(
        n9449) );
  OAI22_X1 U4517 ( .A1(n4373), .A2(n12039), .B1(n17174), .B2(n16824), .ZN(
        n9450) );
  OAI22_X1 U4518 ( .A1(n4370), .A2(n14047), .B1(n17184), .B2(n16824), .ZN(
        n9451) );
  OAI22_X1 U4519 ( .A1(n4367), .A2(n14320), .B1(n17194), .B2(n16824), .ZN(
        n9452) );
  OAI22_X1 U4520 ( .A1(n4362), .A2(n15201), .B1(n17204), .B2(n16824), .ZN(
        n9453) );
  OAI22_X1 U4521 ( .A1(n4462), .A2(n14959), .B1(n16879), .B2(n16828), .ZN(
        n9497) );
  OAI22_X1 U4522 ( .A1(n4459), .A2(n15420), .B1(n16889), .B2(n16828), .ZN(
        n9498) );
  OAI22_X1 U4523 ( .A1(n4451), .A2(n14505), .B1(n16912), .B2(n16828), .ZN(
        n9500) );
  OAI22_X1 U4524 ( .A1(n16920), .A2(n15573), .B1(n16922), .B2(n16828), .ZN(
        n9501) );
  OAI22_X1 U4525 ( .A1(n4438), .A2(n12015), .B1(n16947), .B2(n16829), .ZN(
        n9503) );
  OAI22_X1 U4526 ( .A1(n4435), .A2(n14758), .B1(n16958), .B2(n16829), .ZN(
        n9504) );
  OAI22_X1 U4527 ( .A1(n16966), .A2(n15459), .B1(n16968), .B2(n16829), .ZN(
        n9505) );
  OAI22_X1 U4528 ( .A1(n4429), .A2(n14909), .B1(n16978), .B2(n16829), .ZN(
        n9506) );
  OAI22_X1 U4529 ( .A1(n16999), .A2(n14470), .B1(n17001), .B2(n16829), .ZN(
        n9508) );
  OAI22_X1 U4530 ( .A1(n4420), .A2(n15116), .B1(n17011), .B2(n16829), .ZN(
        n9509) );
  OAI22_X1 U4531 ( .A1(n4382), .A2(n14671), .B1(n17139), .B2(n16830), .ZN(
        n9519) );
  OAI22_X1 U4532 ( .A1(n4376), .A2(n15025), .B1(n17162), .B2(n16830), .ZN(
        n9521) );
  OAI22_X1 U4533 ( .A1(n4373), .A2(n12040), .B1(n17173), .B2(n16830), .ZN(
        n9522) );
  OAI22_X1 U4534 ( .A1(n4370), .A2(n14049), .B1(n17184), .B2(n16830), .ZN(
        n9523) );
  OAI22_X1 U4535 ( .A1(n4367), .A2(n14321), .B1(n17194), .B2(n16830), .ZN(
        n9524) );
  OAI22_X1 U4536 ( .A1(n4362), .A2(n15202), .B1(n17204), .B2(n16830), .ZN(
        n9525) );
  OAI22_X1 U4537 ( .A1(n4462), .A2(n14931), .B1(n16879), .B2(n16834), .ZN(
        n9569) );
  OAI22_X1 U4538 ( .A1(n4459), .A2(n15421), .B1(n16889), .B2(n16834), .ZN(
        n9570) );
  OAI22_X1 U4539 ( .A1(n4451), .A2(n14471), .B1(n16912), .B2(n16834), .ZN(
        n9572) );
  OAI22_X1 U4540 ( .A1(n16920), .A2(n15545), .B1(n16922), .B2(n16834), .ZN(
        n9573) );
  OAI22_X1 U4541 ( .A1(n4438), .A2(n11907), .B1(n16947), .B2(n16835), .ZN(
        n9575) );
  OAI22_X1 U4542 ( .A1(n4435), .A2(n14760), .B1(n16958), .B2(n16835), .ZN(
        n9576) );
  OAI22_X1 U4543 ( .A1(n16966), .A2(n15460), .B1(n16968), .B2(n16835), .ZN(
        n9577) );
  OAI22_X1 U4544 ( .A1(n4429), .A2(n14875), .B1(n16978), .B2(n16835), .ZN(
        n9578) );
  OAI22_X1 U4545 ( .A1(n16999), .A2(n14527), .B1(n17001), .B2(n16835), .ZN(
        n9580) );
  OAI22_X1 U4546 ( .A1(n4420), .A2(n15144), .B1(n17011), .B2(n16835), .ZN(
        n9581) );
  OAI22_X1 U4547 ( .A1(n4382), .A2(n14672), .B1(n17139), .B2(n16836), .ZN(
        n9591) );
  OAI22_X1 U4548 ( .A1(n4376), .A2(n15026), .B1(n17162), .B2(n16836), .ZN(
        n9593) );
  OAI22_X1 U4549 ( .A1(n4373), .A2(n12041), .B1(n17173), .B2(n16836), .ZN(
        n9594) );
  OAI22_X1 U4550 ( .A1(n4370), .A2(n12349), .B1(n17184), .B2(n16836), .ZN(
        n9595) );
  OAI22_X1 U4551 ( .A1(n4367), .A2(n14322), .B1(n17194), .B2(n16836), .ZN(
        n9596) );
  OAI22_X1 U4552 ( .A1(n4362), .A2(n15203), .B1(n17204), .B2(n16836), .ZN(
        n9597) );
  OAI22_X1 U4553 ( .A1(n4462), .A2(n14932), .B1(n16878), .B2(n16840), .ZN(
        n9641) );
  OAI22_X1 U4554 ( .A1(n4459), .A2(n15422), .B1(n16889), .B2(n16840), .ZN(
        n9642) );
  OAI22_X1 U4555 ( .A1(n4451), .A2(n14472), .B1(n16912), .B2(n16840), .ZN(
        n9644) );
  OAI22_X1 U4556 ( .A1(n16920), .A2(n15546), .B1(n16921), .B2(n16840), .ZN(
        n9645) );
  OAI22_X1 U4557 ( .A1(n4438), .A2(n11945), .B1(n16947), .B2(n16841), .ZN(
        n9647) );
  OAI22_X1 U4558 ( .A1(n4435), .A2(n14762), .B1(n16958), .B2(n16841), .ZN(
        n9648) );
  OAI22_X1 U4559 ( .A1(n16966), .A2(n15461), .B1(n16967), .B2(n16841), .ZN(
        n9649) );
  OAI22_X1 U4560 ( .A1(n4429), .A2(n14877), .B1(n16978), .B2(n16841), .ZN(
        n9650) );
  OAI22_X1 U4561 ( .A1(n16999), .A2(n14528), .B1(n17001), .B2(n16841), .ZN(
        n9652) );
  OAI22_X1 U4562 ( .A1(n4420), .A2(n15145), .B1(n17010), .B2(n16841), .ZN(
        n9653) );
  OAI22_X1 U4563 ( .A1(n4382), .A2(n14673), .B1(n17139), .B2(n16842), .ZN(
        n9663) );
  OAI22_X1 U4564 ( .A1(n4376), .A2(n15027), .B1(n17161), .B2(n16842), .ZN(
        n9665) );
  OAI22_X1 U4565 ( .A1(n4373), .A2(n12042), .B1(n17173), .B2(n16842), .ZN(
        n9666) );
  OAI22_X1 U4566 ( .A1(n4370), .A2(n12350), .B1(n17184), .B2(n16842), .ZN(
        n9667) );
  OAI22_X1 U4567 ( .A1(n4367), .A2(n14323), .B1(n17194), .B2(n16842), .ZN(
        n9668) );
  OAI22_X1 U4568 ( .A1(n4362), .A2(n15204), .B1(n17203), .B2(n16842), .ZN(
        n9669) );
  OAI22_X1 U4569 ( .A1(n4462), .A2(n14933), .B1(n16878), .B2(n16846), .ZN(
        n9713) );
  OAI22_X1 U4570 ( .A1(n4459), .A2(n15423), .B1(n16889), .B2(n16846), .ZN(
        n9714) );
  OAI22_X1 U4571 ( .A1(n4451), .A2(n14473), .B1(n16911), .B2(n16846), .ZN(
        n9716) );
  OAI22_X1 U4572 ( .A1(n16920), .A2(n15547), .B1(n16921), .B2(n16846), .ZN(
        n9717) );
  OAI22_X1 U4573 ( .A1(n4438), .A2(n11946), .B1(n16947), .B2(n16847), .ZN(
        n9719) );
  OAI22_X1 U4574 ( .A1(n4435), .A2(n14764), .B1(n16958), .B2(n16847), .ZN(
        n9720) );
  OAI22_X1 U4575 ( .A1(n16966), .A2(n15462), .B1(n16967), .B2(n16847), .ZN(
        n9721) );
  OAI22_X1 U4576 ( .A1(n4429), .A2(n14879), .B1(n16978), .B2(n16847), .ZN(
        n9722) );
  OAI22_X1 U4577 ( .A1(n16999), .A2(n14529), .B1(n17000), .B2(n16847), .ZN(
        n9724) );
  OAI22_X1 U4578 ( .A1(n4420), .A2(n15146), .B1(n17010), .B2(n16847), .ZN(
        n9725) );
  OAI22_X1 U4579 ( .A1(n4382), .A2(n14674), .B1(n17139), .B2(n16848), .ZN(
        n9735) );
  OAI22_X1 U4580 ( .A1(n4376), .A2(n15028), .B1(n17161), .B2(n16848), .ZN(
        n9737) );
  OAI22_X1 U4581 ( .A1(n4373), .A2(n12043), .B1(n17173), .B2(n16848), .ZN(
        n9738) );
  OAI22_X1 U4582 ( .A1(n4370), .A2(n12351), .B1(n17183), .B2(n16848), .ZN(
        n9739) );
  OAI22_X1 U4583 ( .A1(n4367), .A2(n14324), .B1(n17193), .B2(n16848), .ZN(
        n9740) );
  OAI22_X1 U4584 ( .A1(n4362), .A2(n15205), .B1(n17203), .B2(n16848), .ZN(
        n9741) );
  OAI22_X1 U4585 ( .A1(n4462), .A2(n14934), .B1(n16879), .B2(n16852), .ZN(
        n9785) );
  OAI22_X1 U4586 ( .A1(n4459), .A2(n15424), .B1(n16888), .B2(n16852), .ZN(
        n9786) );
  OAI22_X1 U4587 ( .A1(n4451), .A2(n14474), .B1(n16911), .B2(n16852), .ZN(
        n9788) );
  OAI22_X1 U4588 ( .A1(n16920), .A2(n15548), .B1(n16921), .B2(n16852), .ZN(
        n9789) );
  OAI22_X1 U4589 ( .A1(n4438), .A2(n11947), .B1(n16946), .B2(n16853), .ZN(
        n9791) );
  OAI22_X1 U4590 ( .A1(n4435), .A2(n14766), .B1(n16957), .B2(n16853), .ZN(
        n9792) );
  OAI22_X1 U4591 ( .A1(n16966), .A2(n15463), .B1(n16968), .B2(n16853), .ZN(
        n9793) );
  OAI22_X1 U4592 ( .A1(n4429), .A2(n14881), .B1(n16977), .B2(n16853), .ZN(
        n9794) );
  OAI22_X1 U4593 ( .A1(n16999), .A2(n14530), .B1(n17000), .B2(n16853), .ZN(
        n9796) );
  OAI22_X1 U4594 ( .A1(n4420), .A2(n15147), .B1(n17010), .B2(n16853), .ZN(
        n9797) );
  OAI22_X1 U4595 ( .A1(n4382), .A2(n14675), .B1(n17138), .B2(n16854), .ZN(
        n9807) );
  OAI22_X1 U4596 ( .A1(n4376), .A2(n15029), .B1(n17162), .B2(n16854), .ZN(
        n9809) );
  OAI22_X1 U4597 ( .A1(n4373), .A2(n12044), .B1(n17172), .B2(n16854), .ZN(
        n9810) );
  OAI22_X1 U4598 ( .A1(n4370), .A2(n12352), .B1(n17183), .B2(n16854), .ZN(
        n9811) );
  OAI22_X1 U4599 ( .A1(n4367), .A2(n14325), .B1(n17193), .B2(n16854), .ZN(
        n9812) );
  OAI22_X1 U4600 ( .A1(n4362), .A2(n15206), .B1(n17203), .B2(n16854), .ZN(
        n9813) );
  OAI22_X1 U4601 ( .A1(n4462), .A2(n14935), .B1(n16878), .B2(n16858), .ZN(
        n9857) );
  OAI22_X1 U4602 ( .A1(n4459), .A2(n15425), .B1(n16888), .B2(n16858), .ZN(
        n9858) );
  OAI22_X1 U4603 ( .A1(n4451), .A2(n14475), .B1(n16911), .B2(n16858), .ZN(
        n9860) );
  OAI22_X1 U4604 ( .A1(n16920), .A2(n15549), .B1(n16921), .B2(n16858), .ZN(
        n9861) );
  OAI22_X1 U4605 ( .A1(n4438), .A2(n11948), .B1(n16946), .B2(n16859), .ZN(
        n9863) );
  OAI22_X1 U4606 ( .A1(n4435), .A2(n14768), .B1(n16957), .B2(n16859), .ZN(
        n9864) );
  OAI22_X1 U4607 ( .A1(n16966), .A2(n15464), .B1(n16967), .B2(n16859), .ZN(
        n9865) );
  OAI22_X1 U4608 ( .A1(n4429), .A2(n14883), .B1(n16977), .B2(n16859), .ZN(
        n9866) );
  OAI22_X1 U4609 ( .A1(n16999), .A2(n14531), .B1(n17000), .B2(n16859), .ZN(
        n9868) );
  OAI22_X1 U4610 ( .A1(n4420), .A2(n15148), .B1(n17010), .B2(n16859), .ZN(
        n9869) );
  OAI22_X1 U4611 ( .A1(n4382), .A2(n14676), .B1(n17138), .B2(n16860), .ZN(
        n9879) );
  OAI22_X1 U4612 ( .A1(n4376), .A2(n15030), .B1(n17161), .B2(n16860), .ZN(
        n9881) );
  OAI22_X1 U4613 ( .A1(n4373), .A2(n12045), .B1(n17172), .B2(n16860), .ZN(
        n9882) );
  OAI22_X1 U4614 ( .A1(n4370), .A2(n12353), .B1(n17183), .B2(n16860), .ZN(
        n9883) );
  OAI22_X1 U4615 ( .A1(n4367), .A2(n14326), .B1(n17193), .B2(n16860), .ZN(
        n9884) );
  OAI22_X1 U4616 ( .A1(n4362), .A2(n15207), .B1(n17203), .B2(n16860), .ZN(
        n9885) );
  OAI22_X1 U4617 ( .A1(n16877), .A2(n14936), .B1(n16882), .B2(n17513), .ZN(
        n9929) );
  OAI22_X1 U4618 ( .A1(n16887), .A2(n15426), .B1(n16892), .B2(n17513), .ZN(
        n9930) );
  OAI22_X1 U4619 ( .A1(n16910), .A2(n14476), .B1(n16915), .B2(n17513), .ZN(
        n9932) );
  OAI22_X1 U4620 ( .A1(n16920), .A2(n15550), .B1(n16925), .B2(n17513), .ZN(
        n9933) );
  OAI22_X1 U4621 ( .A1(n16945), .A2(n11949), .B1(n16950), .B2(n17514), .ZN(
        n9935) );
  OAI22_X1 U4622 ( .A1(n16956), .A2(n14770), .B1(n16961), .B2(n17514), .ZN(
        n9936) );
  OAI22_X1 U4623 ( .A1(n16966), .A2(n15465), .B1(n16971), .B2(n17514), .ZN(
        n9937) );
  OAI22_X1 U4624 ( .A1(n16976), .A2(n14885), .B1(n16981), .B2(n17514), .ZN(
        n9938) );
  OAI22_X1 U4625 ( .A1(n16999), .A2(n14532), .B1(n17004), .B2(n17514), .ZN(
        n9940) );
  OAI22_X1 U4626 ( .A1(n17009), .A2(n15149), .B1(n17014), .B2(n17514), .ZN(
        n9941) );
  OAI22_X1 U4627 ( .A1(n17137), .A2(n14677), .B1(n17142), .B2(n17515), .ZN(
        n9951) );
  OAI22_X1 U4628 ( .A1(n17160), .A2(n15031), .B1(n17165), .B2(n17515), .ZN(
        n9953) );
  OAI22_X1 U4629 ( .A1(n17171), .A2(n12046), .B1(n17176), .B2(n17515), .ZN(
        n9954) );
  OAI22_X1 U4630 ( .A1(n17182), .A2(n12354), .B1(n17187), .B2(n17515), .ZN(
        n9955) );
  OAI22_X1 U4631 ( .A1(n17192), .A2(n14327), .B1(n17197), .B2(n17515), .ZN(
        n9956) );
  OAI22_X1 U4632 ( .A1(n17202), .A2(n15208), .B1(n17207), .B2(n17515), .ZN(
        n9957) );
  OAI22_X1 U4633 ( .A1(n16928), .A2(n18031), .B1(n15277), .B2(n16920), .ZN(
        n10005) );
  OAI22_X1 U4634 ( .A1(n17023), .A2(n18030), .B1(n12160), .B2(n17025), .ZN(
        n10014) );
  OAI22_X1 U4635 ( .A1(n17075), .A2(n18030), .B1(n15278), .B2(n17077), .ZN(
        n10018) );
  OAI22_X1 U4636 ( .A1(n17088), .A2(n18030), .B1(n15276), .B2(n17090), .ZN(
        n10019) );
  OAI22_X1 U4637 ( .A1(n17101), .A2(n18030), .B1(n11498), .B2(n17103), .ZN(
        n10020) );
  OAI22_X1 U4638 ( .A1(n17114), .A2(n18030), .B1(n12163), .B2(n17116), .ZN(
        n10021) );
  OAI22_X1 U4639 ( .A1(n17127), .A2(n18030), .B1(n15282), .B2(n17129), .ZN(
        n10022) );
  OAI22_X1 U4640 ( .A1(n17229), .A2(n18029), .B1(n15273), .B2(n17231), .ZN(
        n10031) );
  OAI22_X1 U4641 ( .A1(n17242), .A2(n18029), .B1(n12161), .B2(n17244), .ZN(
        n10032) );
  OAI22_X1 U4642 ( .A1(n17255), .A2(n18029), .B1(n14822), .B2(n17257), .ZN(
        n10033) );
  OAI22_X1 U4643 ( .A1(n17307), .A2(n18028), .B1(n15281), .B2(n17309), .ZN(
        n10037) );
  OAI22_X1 U4644 ( .A1(n17320), .A2(n18028), .B1(n15270), .B2(n17322), .ZN(
        n10038) );
  OAI22_X1 U4645 ( .A1(n17333), .A2(n18028), .B1(n11541), .B2(n17335), .ZN(
        n10039) );
  OAI22_X1 U4646 ( .A1(n17359), .A2(n18028), .B1(n15280), .B2(n17361), .ZN(
        n10041) );
  OAI22_X1 U4647 ( .A1(n17385), .A2(n18028), .B1(n14629), .B2(n17387), .ZN(
        n10043) );
  OAI22_X1 U4648 ( .A1(n17424), .A2(n18028), .B1(n15271), .B2(n17426), .ZN(
        n10046) );
  OAI22_X1 U4649 ( .A1(n17437), .A2(n18028), .B1(n12196), .B2(n17439), .ZN(
        n10047) );
  OAI22_X1 U4650 ( .A1(n17451), .A2(n18027), .B1(n14632), .B2(n17452), .ZN(
        n10048) );
  OAI22_X1 U4651 ( .A1(n17463), .A2(n18027), .B1(n15274), .B2(n17465), .ZN(
        n10049) );
  OAI22_X1 U4652 ( .A1(n17476), .A2(n18027), .B1(n15283), .B2(n17478), .ZN(
        n10050) );
  OAI22_X1 U4653 ( .A1(n17489), .A2(n18027), .B1(n14630), .B2(n17491), .ZN(
        n10051) );
  OAI22_X1 U4654 ( .A1(n17502), .A2(n18027), .B1(n15279), .B2(n17504), .ZN(
        n10052) );
  OAI22_X1 U4655 ( .A1(n4462), .A2(n14937), .B1(n16885), .B2(n16706), .ZN(
        n10073) );
  OAI22_X1 U4656 ( .A1(n4459), .A2(n15427), .B1(n16895), .B2(n16706), .ZN(
        n10074) );
  OAI22_X1 U4657 ( .A1(n4451), .A2(n14477), .B1(n16918), .B2(n16706), .ZN(
        n10076) );
  OAI22_X1 U4658 ( .A1(n16920), .A2(n15551), .B1(n16928), .B2(n16706), .ZN(
        n10077) );
  OAI22_X1 U4659 ( .A1(n4438), .A2(n11950), .B1(n16953), .B2(n16706), .ZN(
        n10079) );
  OAI22_X1 U4660 ( .A1(n4435), .A2(n14816), .B1(n16964), .B2(n16706), .ZN(
        n10080) );
  OAI22_X1 U4661 ( .A1(n16966), .A2(n15487), .B1(n16974), .B2(n16706), .ZN(
        n10081) );
  OAI22_X1 U4662 ( .A1(n16976), .A2(n14887), .B1(n16984), .B2(n16706), .ZN(
        n10082) );
  OAI22_X1 U4663 ( .A1(n16999), .A2(n14533), .B1(n17007), .B2(n16705), .ZN(
        n10084) );
  OAI22_X1 U4664 ( .A1(n17009), .A2(n15150), .B1(n17017), .B2(n16705), .ZN(
        n10085) );
  OAI22_X1 U4665 ( .A1(n17137), .A2(n14699), .B1(n17145), .B2(n16705), .ZN(
        n10095) );
  OAI22_X1 U4666 ( .A1(n17160), .A2(n15032), .B1(n17168), .B2(n16704), .ZN(
        n10097) );
  OAI22_X1 U4667 ( .A1(n17170), .A2(n12047), .B1(n17179), .B2(n16704), .ZN(
        n10098) );
  OAI22_X1 U4668 ( .A1(n17182), .A2(n12355), .B1(n17190), .B2(n16704), .ZN(
        n10099) );
  OAI22_X1 U4669 ( .A1(n17192), .A2(n14328), .B1(n17200), .B2(n16704), .ZN(
        n10100) );
  OAI22_X1 U4670 ( .A1(n17202), .A2(n15209), .B1(n17210), .B2(n16704), .ZN(
        n10101) );
  INV_X1 U4671 ( .A(N46298), .ZN(n13978) );
  INV_X1 U4672 ( .A(N45784), .ZN(n12497) );
  NAND2_X1 U4673 ( .A1(n14091), .A2(n14149), .ZN(n4175) );
  NAND2_X1 U4674 ( .A1(n14091), .A2(n14150), .ZN(n4186) );
  NAND2_X1 U4675 ( .A1(n14140), .A2(n14196), .ZN(n14120) );
  NAND2_X1 U4676 ( .A1(n14128), .A2(n14196), .ZN(n14166) );
  NAND2_X1 U4677 ( .A1(n14146), .A2(n14196), .ZN(n14163) );
  NOR2_X1 U4678 ( .A1(n13973), .A2(n13974), .ZN(n12624) );
  NAND2_X1 U4679 ( .A1(n14137), .A2(n14020), .ZN(n14117) );
  NAND2_X1 U4680 ( .A1(n14202), .A2(n14020), .ZN(n14125) );
  NAND2_X1 U4681 ( .A1(n14138), .A2(n14020), .ZN(n14123) );
  NAND2_X1 U4682 ( .A1(n14143), .A2(n14020), .ZN(n14160) );
  NAND2_X1 U4683 ( .A1(n14150), .A2(n14151), .ZN(n4173) );
  NAND2_X1 U4684 ( .A1(n14149), .A2(n14151), .ZN(n4242) );
  NAND2_X1 U4685 ( .A1(datain[0]), .A2(n18039), .ZN(n12338) );
  NAND2_X1 U4686 ( .A1(datain[1]), .A2(n18039), .ZN(n12184) );
  NAND2_X1 U4687 ( .A1(datain[2]), .A2(n18039), .ZN(n12029) );
  NOR2_X1 U4688 ( .A1(n18050), .A2(n14006), .ZN(n4090) );
  OR2_X1 U4689 ( .A1(n14144), .A2(n14020), .ZN(n14124) );
  AND2_X1 U4690 ( .A1(n14143), .A2(N9925), .ZN(n14108) );
  NAND2_X1 U4691 ( .A1(n14130), .A2(n14146), .ZN(n14136) );
  INV_X1 U4692 ( .A(N46299), .ZN(n13979) );
  INV_X1 U4693 ( .A(N45785), .ZN(n12498) );
  INV_X1 U4694 ( .A(N276), .ZN(n14234) );
  AND2_X1 U4695 ( .A1(n14094), .A2(n14105), .ZN(n4123) );
  AND2_X1 U4696 ( .A1(n14104), .A2(n14105), .ZN(n4124) );
  AND2_X1 U4697 ( .A1(n14108), .A2(n14105), .ZN(n4130) );
  AND2_X1 U4698 ( .A1(n14107), .A2(n14105), .ZN(n4131) );
  INV_X1 U4699 ( .A(n14263), .ZN(n14262) );
  AND2_X1 U4700 ( .A1(n14194), .A2(n14178), .ZN(n14170) );
  INV_X1 U4701 ( .A(n14146), .ZN(n14172) );
  NAND2_X1 U4702 ( .A1(n13903), .A2(n13901), .ZN(n12522) );
  NAND2_X1 U4703 ( .A1(n12422), .A2(n12420), .ZN(n10519) );
  NAND2_X1 U4704 ( .A1(n13901), .A2(n13902), .ZN(n12523) );
  NAND2_X1 U4705 ( .A1(n12420), .A2(n12421), .ZN(n10520) );
  AND2_X1 U4706 ( .A1(n14091), .A2(n14152), .ZN(n4170) );
  AND2_X1 U4707 ( .A1(n14091), .A2(n14092), .ZN(n4107) );
  AND2_X1 U4708 ( .A1(N9921), .A2(n14209), .ZN(n14137) );
  AND2_X1 U4709 ( .A1(n14152), .A2(n14151), .ZN(n4171) );
  OAI21_X1 U4710 ( .B1(n18051), .B2(n14821), .A(n13997), .ZN(n10185) );
  AND2_X1 U4711 ( .A1(N9923), .A2(N9921), .ZN(n14143) );
  NAND2_X1 U4712 ( .A1(datain[4]), .A2(n18038), .ZN(n10425) );
  AND2_X1 U4713 ( .A1(n13904), .A2(n13985), .ZN(n12524) );
  AND2_X1 U4714 ( .A1(n13904), .A2(n13902), .ZN(n12525) );
  AND2_X1 U4715 ( .A1(n12423), .A2(n12421), .ZN(n10523) );
  AND2_X1 U4716 ( .A1(n12423), .A2(n12504), .ZN(n10522) );
  AND2_X1 U4717 ( .A1(n13903), .A2(n13904), .ZN(n12520) );
  AND2_X1 U4718 ( .A1(n13905), .A2(n13904), .ZN(n12634) );
  AND2_X1 U4719 ( .A1(n12422), .A2(n12423), .ZN(n10517) );
  AND2_X1 U4720 ( .A1(n12424), .A2(n12423), .ZN(n10663) );
  AND2_X1 U4721 ( .A1(n13901), .A2(n13985), .ZN(n12633) );
  AND2_X1 U4722 ( .A1(n12420), .A2(n12504), .ZN(n10662) );
  AND2_X1 U4723 ( .A1(n13905), .A2(n13901), .ZN(n12519) );
  AND2_X1 U4724 ( .A1(n12424), .A2(n12420), .ZN(n10516) );
  NAND2_X1 U4725 ( .A1(n12492), .A2(n12507), .ZN(n12500) );
  INV_X1 U4726 ( .A(n12493), .ZN(n12507) );
  BUF_X1 U4727 ( .A(reset), .Z(n18032) );
  NAND2_X1 U4728 ( .A1(n13973), .A2(n13988), .ZN(n13981) );
  INV_X1 U4729 ( .A(n13974), .ZN(n13988) );
  INV_X1 U4730 ( .A(N9923), .ZN(n14209) );
  INV_X1 U4731 ( .A(n14114), .ZN(n4150) );
  OAI22_X1 U4732 ( .A1(n14115), .A2(n14116), .B1(n14117), .B2(n14118), .ZN(
        n14114) );
  INV_X1 U4733 ( .A(N46300), .ZN(n13976) );
  INV_X1 U4734 ( .A(N45786), .ZN(n12495) );
  INV_X1 U4735 ( .A(N274), .ZN(n14259) );
  INV_X1 U4736 ( .A(N46301), .ZN(n13975) );
  INV_X1 U4737 ( .A(N45787), .ZN(n12494) );
  INV_X1 U4738 ( .A(N275), .ZN(n14257) );
  INV_X1 U4739 ( .A(n14119), .ZN(n4148) );
  OAI22_X1 U4740 ( .A1(n14120), .A2(n14115), .B1(n14121), .B2(n14117), .ZN(
        n14119) );
  INV_X1 U4741 ( .A(n14195), .ZN(n4222) );
  OAI22_X1 U4742 ( .A1(n14166), .A2(n14115), .B1(n14167), .B2(n14117), .ZN(
        n14195) );
  NAND2_X1 U4743 ( .A1(datain[5]), .A2(n18038), .ZN(n10315) );
  AND2_X1 U4744 ( .A1(n14147), .A2(n14820), .ZN(n14130) );
  INV_X1 U4745 ( .A(n14128), .ZN(n14100) );
  NAND2_X1 U4746 ( .A1(datain[3]), .A2(n18038), .ZN(n11868) );
  INV_X1 U4747 ( .A(N46303), .ZN(n13963) );
  INV_X1 U4748 ( .A(N45789), .ZN(n12482) );
  INV_X1 U4749 ( .A(\add_73/carry[5] ), .ZN(n14265) );
  INV_X1 U4750 ( .A(n14006), .ZN(n14233) );
  INV_X1 U4751 ( .A(n14247), .ZN(n14239) );
  INV_X1 U4752 ( .A(n14149), .ZN(n14186) );
  INV_X1 U4753 ( .A(n14150), .ZN(n14184) );
  INV_X1 U4754 ( .A(N45788), .ZN(n12499) );
  INV_X1 U4755 ( .A(N46302), .ZN(n13980) );
  NOR2_X1 U4756 ( .A1(N9908), .A2(n14022), .ZN(n14017) );
  NOR2_X1 U4757 ( .A1(n18050), .A2(datain[0]), .ZN(n12302) );
  NOR2_X1 U4758 ( .A1(n18050), .A2(datain[1]), .ZN(n12149) );
  NOR2_X1 U4759 ( .A1(n18050), .A2(datain[2]), .ZN(n11996) );
  INV_X1 U4760 ( .A(datain[4]), .ZN(n10400) );
  INV_X1 U4761 ( .A(datain[5]), .ZN(n10290) );
  INV_X1 U4762 ( .A(datain[6]), .ZN(n10285) );
  INV_X1 U4763 ( .A(datain[3]), .ZN(n11843) );
  AOI221_X1 U4764 ( .B1(\registers[56][1] ), .B2(n16517), .C1(
        \registers[60][1] ), .C2(n16514), .A(n12297), .ZN(n12296) );
  OAI222_X1 U4765 ( .A1(n16511), .A2(n14570), .B1(n16508), .B2(n12052), .C1(
        n16505), .C2(n15243), .ZN(n12297) );
  AOI221_X1 U4766 ( .B1(\registers[56][2] ), .B2(n16517), .C1(
        \registers[60][2] ), .C2(n16514), .A(n12144), .ZN(n12143) );
  OAI222_X1 U4767 ( .A1(n16511), .A2(n14571), .B1(n16508), .B2(n12053), .C1(
        n16505), .C2(n15244), .ZN(n12144) );
  AOI221_X1 U4768 ( .B1(\registers[56][3] ), .B2(n16517), .C1(
        \registers[60][3] ), .C2(n16514), .A(n11991), .ZN(n11990) );
  OAI222_X1 U4769 ( .A1(n16511), .A2(n14572), .B1(n16508), .B2(n12054), .C1(
        n16505), .C2(n15240), .ZN(n11991) );
  NOR2_X1 U4770 ( .A1(N9910), .A2(n10189), .ZN(n14140) );
  AOI221_X1 U4771 ( .B1(\registers[2][0] ), .B2(n16364), .C1(
        \registers[29][0] ), .C2(n16361), .A(n13942), .ZN(n13941) );
  OAI222_X1 U4772 ( .A1(n16358), .A2(n15004), .B1(n16355), .B2(n14300), .C1(
        n16352), .C2(n12018), .ZN(n13942) );
  AOI221_X1 U4773 ( .B1(\registers[56][0] ), .B2(n16265), .C1(
        \registers[60][0] ), .C2(n16262), .A(n13968), .ZN(n13967) );
  OAI222_X1 U4774 ( .A1(n16259), .A2(n14573), .B1(n16256), .B2(n12055), .C1(
        n16253), .C2(n15245), .ZN(n13968) );
  AOI221_X1 U4775 ( .B1(\registers[2][1] ), .B2(n16364), .C1(
        \registers[29][1] ), .C2(n16361), .A(n13877), .ZN(n13876) );
  OAI222_X1 U4776 ( .A1(n16358), .A2(n15005), .B1(n16355), .B2(n14301), .C1(
        n16352), .C2(n12019), .ZN(n13877) );
  AOI221_X1 U4777 ( .B1(\registers[56][1] ), .B2(n16265), .C1(
        \registers[60][1] ), .C2(n16262), .A(n13893), .ZN(n13892) );
  OAI222_X1 U4778 ( .A1(n16259), .A2(n14570), .B1(n16256), .B2(n12052), .C1(
        n16253), .C2(n15243), .ZN(n13893) );
  AOI221_X1 U4779 ( .B1(\registers[2][2] ), .B2(n16364), .C1(
        \registers[29][2] ), .C2(n16361), .A(n13835), .ZN(n13834) );
  OAI222_X1 U4780 ( .A1(n16358), .A2(n15006), .B1(n16355), .B2(n14302), .C1(
        n16352), .C2(n12020), .ZN(n13835) );
  AOI221_X1 U4781 ( .B1(\registers[56][2] ), .B2(n16265), .C1(
        \registers[60][2] ), .C2(n16262), .A(n13851), .ZN(n13850) );
  OAI222_X1 U4782 ( .A1(n16259), .A2(n14571), .B1(n16256), .B2(n12053), .C1(
        n16253), .C2(n15244), .ZN(n13851) );
  AOI221_X1 U4783 ( .B1(\registers[2][3] ), .B2(n16364), .C1(
        \registers[29][3] ), .C2(n16361), .A(n13793), .ZN(n13792) );
  OAI222_X1 U4784 ( .A1(n16358), .A2(n14989), .B1(n16355), .B2(n14282), .C1(
        n16352), .C2(n12016), .ZN(n13793) );
  AOI221_X1 U4785 ( .B1(\registers[56][3] ), .B2(n16265), .C1(
        \registers[60][3] ), .C2(n16262), .A(n13809), .ZN(n13808) );
  OAI222_X1 U4786 ( .A1(n16259), .A2(n14572), .B1(n16256), .B2(n12054), .C1(
        n16253), .C2(n15240), .ZN(n13809) );
  AOI221_X1 U4787 ( .B1(\registers[2][4] ), .B2(n16364), .C1(
        \registers[29][4] ), .C2(n16361), .A(n13751), .ZN(n13750) );
  OAI222_X1 U4788 ( .A1(n16358), .A2(n14990), .B1(n16355), .B2(n14283), .C1(
        n16352), .C2(n12017), .ZN(n13751) );
  AOI221_X1 U4789 ( .B1(\registers[56][4] ), .B2(n16265), .C1(
        \registers[60][4] ), .C2(n16262), .A(n13767), .ZN(n13766) );
  OAI222_X1 U4790 ( .A1(n16259), .A2(n14538), .B1(n16256), .B2(n12050), .C1(
        n16253), .C2(n15241), .ZN(n13767) );
  AOI221_X1 U4791 ( .B1(\registers[2][5] ), .B2(n16364), .C1(
        \registers[29][5] ), .C2(n16361), .A(n13709), .ZN(n13708) );
  OAI222_X1 U4792 ( .A1(n16358), .A2(n15007), .B1(n16355), .B2(n14303), .C1(
        n16352), .C2(n12021), .ZN(n13709) );
  AOI221_X1 U4793 ( .B1(\registers[56][5] ), .B2(n16265), .C1(
        \registers[60][5] ), .C2(n16262), .A(n13725), .ZN(n13724) );
  OAI222_X1 U4794 ( .A1(n16259), .A2(n14539), .B1(n16256), .B2(n12051), .C1(
        n16253), .C2(n15242), .ZN(n13725) );
  AOI221_X1 U4795 ( .B1(\registers[2][6] ), .B2(n16364), .C1(
        \registers[29][6] ), .C2(n16361), .A(n13667), .ZN(n13666) );
  OAI222_X1 U4796 ( .A1(n16358), .A2(n15008), .B1(n16355), .B2(n14304), .C1(
        n16352), .C2(n12022), .ZN(n13667) );
  AOI221_X1 U4797 ( .B1(\registers[56][6] ), .B2(n16265), .C1(
        \registers[60][6] ), .C2(n16262), .A(n13683), .ZN(n13682) );
  OAI222_X1 U4798 ( .A1(n16259), .A2(n14574), .B1(n16256), .B2(n12056), .C1(
        n16253), .C2(n15246), .ZN(n13683) );
  AOI221_X1 U4799 ( .B1(\registers[2][7] ), .B2(n16364), .C1(
        \registers[29][7] ), .C2(n16361), .A(n13625), .ZN(n13624) );
  OAI222_X1 U4800 ( .A1(n16358), .A2(n15009), .B1(n16355), .B2(n14305), .C1(
        n16352), .C2(n12023), .ZN(n13625) );
  AOI221_X1 U4801 ( .B1(\registers[56][7] ), .B2(n16265), .C1(
        \registers[60][7] ), .C2(n16262), .A(n13641), .ZN(n13640) );
  OAI222_X1 U4802 ( .A1(n16259), .A2(n14575), .B1(n16256), .B2(n12057), .C1(
        n16253), .C2(n15247), .ZN(n13641) );
  AOI221_X1 U4803 ( .B1(\registers[2][8] ), .B2(n16364), .C1(
        \registers[29][8] ), .C2(n16361), .A(n13583), .ZN(n13582) );
  OAI222_X1 U4804 ( .A1(n16358), .A2(n15010), .B1(n16355), .B2(n14306), .C1(
        n16352), .C2(n12024), .ZN(n13583) );
  AOI221_X1 U4805 ( .B1(\registers[56][8] ), .B2(n16265), .C1(
        \registers[60][8] ), .C2(n16262), .A(n13599), .ZN(n13598) );
  OAI222_X1 U4806 ( .A1(n16259), .A2(n14576), .B1(n16256), .B2(n12058), .C1(
        n16253), .C2(n15248), .ZN(n13599) );
  AOI221_X1 U4807 ( .B1(\registers[2][9] ), .B2(n16364), .C1(
        \registers[29][9] ), .C2(n16361), .A(n13541), .ZN(n13540) );
  OAI222_X1 U4808 ( .A1(n16358), .A2(n15011), .B1(n16355), .B2(n14307), .C1(
        n16352), .C2(n12025), .ZN(n13541) );
  AOI221_X1 U4809 ( .B1(\registers[56][9] ), .B2(n16265), .C1(
        \registers[60][9] ), .C2(n16262), .A(n13557), .ZN(n13556) );
  OAI222_X1 U4810 ( .A1(n16259), .A2(n14577), .B1(n16256), .B2(n12059), .C1(
        n16253), .C2(n15249), .ZN(n13557) );
  AOI221_X1 U4811 ( .B1(\registers[2][10] ), .B2(n16364), .C1(
        \registers[29][10] ), .C2(n16361), .A(n13499), .ZN(n13498) );
  OAI222_X1 U4812 ( .A1(n16358), .A2(n15012), .B1(n16355), .B2(n14308), .C1(
        n16352), .C2(n12026), .ZN(n13499) );
  AOI221_X1 U4813 ( .B1(\registers[56][10] ), .B2(n16265), .C1(
        \registers[60][10] ), .C2(n16262), .A(n13515), .ZN(n13514) );
  OAI222_X1 U4814 ( .A1(n16259), .A2(n14578), .B1(n16256), .B2(n12060), .C1(
        n16253), .C2(n15250), .ZN(n13515) );
  AOI221_X1 U4815 ( .B1(\registers[2][11] ), .B2(n16364), .C1(
        \registers[29][11] ), .C2(n16361), .A(n13457), .ZN(n13456) );
  OAI222_X1 U4816 ( .A1(n16358), .A2(n15013), .B1(n16355), .B2(n14309), .C1(
        n16352), .C2(n12027), .ZN(n13457) );
  AOI221_X1 U4817 ( .B1(\registers[56][11] ), .B2(n16265), .C1(
        \registers[60][11] ), .C2(n16262), .A(n13473), .ZN(n13472) );
  OAI222_X1 U4818 ( .A1(n16259), .A2(n14579), .B1(n16256), .B2(n12098), .C1(
        n16253), .C2(n15251), .ZN(n13473) );
  AOI221_X1 U4819 ( .B1(\registers[2][12] ), .B2(n16365), .C1(
        \registers[29][12] ), .C2(n16362), .A(n13415), .ZN(n13414) );
  OAI222_X1 U4820 ( .A1(n16359), .A2(n15014), .B1(n16356), .B2(n14310), .C1(
        n16353), .C2(n12028), .ZN(n13415) );
  AOI221_X1 U4821 ( .B1(\registers[56][12] ), .B2(n16266), .C1(
        \registers[60][12] ), .C2(n16263), .A(n13431), .ZN(n13430) );
  OAI222_X1 U4822 ( .A1(n16260), .A2(n14580), .B1(n16257), .B2(n12099), .C1(
        n16254), .C2(n15252), .ZN(n13431) );
  AOI221_X1 U4823 ( .B1(\registers[2][13] ), .B2(n16365), .C1(
        \registers[29][13] ), .C2(n16362), .A(n13373), .ZN(n13372) );
  OAI222_X1 U4824 ( .A1(n16359), .A2(n15015), .B1(n16356), .B2(n14311), .C1(
        n16353), .C2(n12030), .ZN(n13373) );
  AOI221_X1 U4825 ( .B1(\registers[56][13] ), .B2(n16266), .C1(
        \registers[60][13] ), .C2(n16263), .A(n13389), .ZN(n13388) );
  OAI222_X1 U4826 ( .A1(n16260), .A2(n14581), .B1(n16257), .B2(n12100), .C1(
        n16254), .C2(n15253), .ZN(n13389) );
  AOI221_X1 U4827 ( .B1(\registers[2][14] ), .B2(n16365), .C1(
        \registers[29][14] ), .C2(n16362), .A(n13331), .ZN(n13330) );
  OAI222_X1 U4828 ( .A1(n16359), .A2(n15016), .B1(n16356), .B2(n14312), .C1(
        n16353), .C2(n12031), .ZN(n13331) );
  AOI221_X1 U4829 ( .B1(\registers[56][14] ), .B2(n16266), .C1(
        \registers[60][14] ), .C2(n16263), .A(n13347), .ZN(n13346) );
  OAI222_X1 U4830 ( .A1(n16260), .A2(n14582), .B1(n16257), .B2(n12101), .C1(
        n16254), .C2(n15254), .ZN(n13347) );
  AOI221_X1 U4831 ( .B1(\registers[2][15] ), .B2(n16365), .C1(
        \registers[29][15] ), .C2(n16362), .A(n13289), .ZN(n13288) );
  OAI222_X1 U4832 ( .A1(n16359), .A2(n15017), .B1(n16356), .B2(n14313), .C1(
        n16353), .C2(n12032), .ZN(n13289) );
  AOI221_X1 U4833 ( .B1(\registers[56][15] ), .B2(n16266), .C1(
        \registers[60][15] ), .C2(n16263), .A(n13305), .ZN(n13304) );
  OAI222_X1 U4834 ( .A1(n16260), .A2(n14583), .B1(n16257), .B2(n12102), .C1(
        n16254), .C2(n15255), .ZN(n13305) );
  AOI221_X1 U4835 ( .B1(\registers[2][16] ), .B2(n16365), .C1(
        \registers[29][16] ), .C2(n16362), .A(n13247), .ZN(n13246) );
  OAI222_X1 U4836 ( .A1(n16359), .A2(n15018), .B1(n16356), .B2(n14314), .C1(
        n16353), .C2(n12033), .ZN(n13247) );
  AOI221_X1 U4837 ( .B1(\registers[56][16] ), .B2(n16266), .C1(
        \registers[60][16] ), .C2(n16263), .A(n13263), .ZN(n13262) );
  OAI222_X1 U4838 ( .A1(n16260), .A2(n14584), .B1(n16257), .B2(n12103), .C1(
        n16254), .C2(n15256), .ZN(n13263) );
  AOI221_X1 U4839 ( .B1(\registers[2][17] ), .B2(n16365), .C1(
        \registers[29][17] ), .C2(n16362), .A(n13205), .ZN(n13204) );
  OAI222_X1 U4840 ( .A1(n16359), .A2(n15019), .B1(n16356), .B2(n14315), .C1(
        n16353), .C2(n12034), .ZN(n13205) );
  AOI221_X1 U4841 ( .B1(\registers[56][17] ), .B2(n16266), .C1(
        \registers[60][17] ), .C2(n16263), .A(n13221), .ZN(n13220) );
  OAI222_X1 U4842 ( .A1(n16260), .A2(n14585), .B1(n16257), .B2(n12104), .C1(
        n16254), .C2(n15257), .ZN(n13221) );
  AOI221_X1 U4843 ( .B1(\registers[2][18] ), .B2(n16365), .C1(
        \registers[29][18] ), .C2(n16362), .A(n13163), .ZN(n13162) );
  OAI222_X1 U4844 ( .A1(n16359), .A2(n15020), .B1(n16356), .B2(n14316), .C1(
        n16353), .C2(n12035), .ZN(n13163) );
  AOI221_X1 U4845 ( .B1(\registers[56][18] ), .B2(n16266), .C1(
        \registers[60][18] ), .C2(n16263), .A(n13179), .ZN(n13178) );
  OAI222_X1 U4846 ( .A1(n16260), .A2(n14586), .B1(n16257), .B2(n12105), .C1(
        n16254), .C2(n15258), .ZN(n13179) );
  AOI221_X1 U4847 ( .B1(\registers[2][19] ), .B2(n16365), .C1(
        \registers[29][19] ), .C2(n16362), .A(n13121), .ZN(n13120) );
  OAI222_X1 U4848 ( .A1(n16359), .A2(n15021), .B1(n16356), .B2(n14317), .C1(
        n16353), .C2(n12036), .ZN(n13121) );
  AOI221_X1 U4849 ( .B1(\registers[56][19] ), .B2(n16266), .C1(
        \registers[60][19] ), .C2(n16263), .A(n13137), .ZN(n13136) );
  OAI222_X1 U4850 ( .A1(n16260), .A2(n14587), .B1(n16257), .B2(n12148), .C1(
        n16254), .C2(n15259), .ZN(n13137) );
  AOI221_X1 U4851 ( .B1(\registers[2][20] ), .B2(n16365), .C1(
        \registers[29][20] ), .C2(n16362), .A(n13079), .ZN(n13078) );
  OAI222_X1 U4852 ( .A1(n16359), .A2(n15022), .B1(n16356), .B2(n14318), .C1(
        n16353), .C2(n12037), .ZN(n13079) );
  AOI221_X1 U4853 ( .B1(\registers[56][20] ), .B2(n16266), .C1(
        \registers[60][20] ), .C2(n16263), .A(n13095), .ZN(n13094) );
  OAI222_X1 U4854 ( .A1(n16260), .A2(n14588), .B1(n16257), .B2(n12150), .C1(
        n16254), .C2(n15260), .ZN(n13095) );
  AOI221_X1 U4855 ( .B1(\registers[2][21] ), .B2(n16365), .C1(
        \registers[29][21] ), .C2(n16362), .A(n13037), .ZN(n13036) );
  OAI222_X1 U4856 ( .A1(n16359), .A2(n15023), .B1(n16356), .B2(n14319), .C1(
        n16353), .C2(n12038), .ZN(n13037) );
  AOI221_X1 U4857 ( .B1(\registers[56][21] ), .B2(n16266), .C1(
        \registers[60][21] ), .C2(n16263), .A(n13053), .ZN(n13052) );
  OAI222_X1 U4858 ( .A1(n16260), .A2(n14589), .B1(n16257), .B2(n12151), .C1(
        n16254), .C2(n15261), .ZN(n13053) );
  AOI221_X1 U4859 ( .B1(\registers[2][22] ), .B2(n16365), .C1(
        \registers[29][22] ), .C2(n16362), .A(n12995), .ZN(n12994) );
  OAI222_X1 U4860 ( .A1(n16359), .A2(n15024), .B1(n16356), .B2(n14320), .C1(
        n16353), .C2(n12039), .ZN(n12995) );
  AOI221_X1 U4861 ( .B1(\registers[56][22] ), .B2(n16266), .C1(
        \registers[60][22] ), .C2(n16263), .A(n13011), .ZN(n13010) );
  OAI222_X1 U4862 ( .A1(n16260), .A2(n14590), .B1(n16257), .B2(n12152), .C1(
        n16254), .C2(n15262), .ZN(n13011) );
  AOI221_X1 U4863 ( .B1(\registers[2][23] ), .B2(n16365), .C1(
        \registers[29][23] ), .C2(n16362), .A(n12953), .ZN(n12952) );
  OAI222_X1 U4864 ( .A1(n16359), .A2(n15025), .B1(n16356), .B2(n14321), .C1(
        n16353), .C2(n12040), .ZN(n12953) );
  AOI221_X1 U4865 ( .B1(\registers[56][23] ), .B2(n16266), .C1(
        \registers[60][23] ), .C2(n16263), .A(n12969), .ZN(n12968) );
  OAI222_X1 U4866 ( .A1(n16260), .A2(n14591), .B1(n16257), .B2(n12153), .C1(
        n16254), .C2(n15263), .ZN(n12969) );
  AOI221_X1 U4867 ( .B1(\registers[2][24] ), .B2(n16366), .C1(
        \registers[29][24] ), .C2(n16363), .A(n12911), .ZN(n12910) );
  OAI222_X1 U4868 ( .A1(n16360), .A2(n15026), .B1(n16357), .B2(n14322), .C1(
        n16354), .C2(n12041), .ZN(n12911) );
  AOI221_X1 U4869 ( .B1(\registers[12][24] ), .B2(n16411), .C1(
        \registers[17][24] ), .C2(n16408), .A(n12903), .ZN(n12902) );
  OAI22_X1 U4870 ( .A1(n16405), .A2(n15065), .B1(n16402), .B2(n14419), .ZN(
        n12903) );
  AOI221_X1 U4871 ( .B1(\registers[56][24] ), .B2(n16267), .C1(
        \registers[60][24] ), .C2(n16264), .A(n12927), .ZN(n12926) );
  OAI222_X1 U4872 ( .A1(n16261), .A2(n14592), .B1(n16258), .B2(n12154), .C1(
        n16255), .C2(n15264), .ZN(n12927) );
  AOI221_X1 U4873 ( .B1(\registers[2][25] ), .B2(n16366), .C1(
        \registers[29][25] ), .C2(n16363), .A(n12869), .ZN(n12868) );
  OAI222_X1 U4874 ( .A1(n16360), .A2(n15027), .B1(n16357), .B2(n14323), .C1(
        n16354), .C2(n12042), .ZN(n12869) );
  AOI221_X1 U4875 ( .B1(\registers[12][25] ), .B2(n16411), .C1(
        \registers[17][25] ), .C2(n16408), .A(n12861), .ZN(n12860) );
  OAI22_X1 U4876 ( .A1(n16405), .A2(n15066), .B1(n16402), .B2(n14420), .ZN(
        n12861) );
  AOI221_X1 U4877 ( .B1(\registers[56][25] ), .B2(n16267), .C1(
        \registers[60][25] ), .C2(n16264), .A(n12885), .ZN(n12884) );
  OAI222_X1 U4878 ( .A1(n16261), .A2(n14593), .B1(n16258), .B2(n12155), .C1(
        n16255), .C2(n15265), .ZN(n12885) );
  AOI221_X1 U4879 ( .B1(\registers[2][26] ), .B2(n16366), .C1(
        \registers[29][26] ), .C2(n16363), .A(n12827), .ZN(n12826) );
  OAI222_X1 U4880 ( .A1(n16360), .A2(n15028), .B1(n16357), .B2(n14324), .C1(
        n16354), .C2(n12043), .ZN(n12827) );
  AOI221_X1 U4881 ( .B1(\registers[12][26] ), .B2(n16411), .C1(
        \registers[17][26] ), .C2(n16408), .A(n12819), .ZN(n12818) );
  OAI22_X1 U4882 ( .A1(n16405), .A2(n15067), .B1(n16402), .B2(n14421), .ZN(
        n12819) );
  AOI221_X1 U4883 ( .B1(\registers[56][26] ), .B2(n16267), .C1(
        \registers[60][26] ), .C2(n16264), .A(n12843), .ZN(n12842) );
  OAI222_X1 U4884 ( .A1(n16261), .A2(n14594), .B1(n16258), .B2(n12156), .C1(
        n16255), .C2(n15266), .ZN(n12843) );
  AOI221_X1 U4885 ( .B1(\registers[2][27] ), .B2(n16366), .C1(
        \registers[29][27] ), .C2(n16363), .A(n12785), .ZN(n12784) );
  OAI222_X1 U4886 ( .A1(n16360), .A2(n15029), .B1(n16357), .B2(n14325), .C1(
        n16354), .C2(n12044), .ZN(n12785) );
  AOI221_X1 U4887 ( .B1(\registers[12][27] ), .B2(n16411), .C1(
        \registers[17][27] ), .C2(n16408), .A(n12777), .ZN(n12776) );
  OAI22_X1 U4888 ( .A1(n16405), .A2(n15068), .B1(n16402), .B2(n14422), .ZN(
        n12777) );
  AOI221_X1 U4889 ( .B1(\registers[56][27] ), .B2(n16267), .C1(
        \registers[60][27] ), .C2(n16264), .A(n12801), .ZN(n12800) );
  OAI222_X1 U4890 ( .A1(n16261), .A2(n14595), .B1(n16258), .B2(n12157), .C1(
        n16255), .C2(n15267), .ZN(n12801) );
  AOI221_X1 U4891 ( .B1(\registers[2][28] ), .B2(n16366), .C1(
        \registers[29][28] ), .C2(n16363), .A(n12743), .ZN(n12742) );
  OAI222_X1 U4892 ( .A1(n16360), .A2(n15030), .B1(n16357), .B2(n14326), .C1(
        n16354), .C2(n12045), .ZN(n12743) );
  AOI221_X1 U4893 ( .B1(\registers[12][28] ), .B2(n16411), .C1(
        \registers[17][28] ), .C2(n16408), .A(n12735), .ZN(n12734) );
  OAI22_X1 U4894 ( .A1(n16405), .A2(n15069), .B1(n16402), .B2(n14423), .ZN(
        n12735) );
  AOI221_X1 U4895 ( .B1(\registers[56][28] ), .B2(n16267), .C1(
        \registers[60][28] ), .C2(n16264), .A(n12759), .ZN(n12758) );
  OAI222_X1 U4896 ( .A1(n16261), .A2(n14596), .B1(n16258), .B2(n12158), .C1(
        n16255), .C2(n15268), .ZN(n12759) );
  AOI221_X1 U4897 ( .B1(\registers[2][29] ), .B2(n16366), .C1(
        \registers[29][29] ), .C2(n16363), .A(n12701), .ZN(n12700) );
  OAI222_X1 U4898 ( .A1(n16360), .A2(n15031), .B1(n16357), .B2(n14327), .C1(
        n16354), .C2(n12046), .ZN(n12701) );
  AOI221_X1 U4899 ( .B1(\registers[12][29] ), .B2(n16411), .C1(
        \registers[17][29] ), .C2(n16408), .A(n12693), .ZN(n12692) );
  OAI22_X1 U4900 ( .A1(n16405), .A2(n15070), .B1(n16402), .B2(n14424), .ZN(
        n12693) );
  AOI221_X1 U4901 ( .B1(\registers[56][29] ), .B2(n16267), .C1(
        \registers[60][29] ), .C2(n16264), .A(n12717), .ZN(n12716) );
  OAI222_X1 U4902 ( .A1(n16261), .A2(n14597), .B1(n16258), .B2(n12159), .C1(
        n16255), .C2(n15269), .ZN(n12717) );
  AOI221_X1 U4903 ( .B1(\registers[2][30] ), .B2(n16366), .C1(
        \registers[29][30] ), .C2(n16363), .A(n12658), .ZN(n12657) );
  OAI222_X1 U4904 ( .A1(n16360), .A2(n14857), .B1(n16357), .B2(n14054), .C1(
        n16354), .C2(n11904), .ZN(n12658) );
  AOI221_X1 U4905 ( .B1(\registers[12][30] ), .B2(n16411), .C1(
        \registers[17][30] ), .C2(n16408), .A(n12649), .ZN(n12648) );
  OAI22_X1 U4906 ( .A1(n16405), .A2(n14870), .B1(n16402), .B2(n14060), .ZN(
        n12649) );
  AOI221_X1 U4907 ( .B1(\registers[56][30] ), .B2(n16267), .C1(
        \registers[60][30] ), .C2(n16264), .A(n12675), .ZN(n12674) );
  OAI222_X1 U4908 ( .A1(n16261), .A2(n14534), .B1(n16258), .B2(n12048), .C1(
        n16255), .C2(n15033), .ZN(n12675) );
  AOI221_X1 U4909 ( .B1(\registers[2][31] ), .B2(n16366), .C1(
        \registers[29][31] ), .C2(n16363), .A(n12563), .ZN(n12560) );
  OAI222_X1 U4910 ( .A1(n16360), .A2(n15032), .B1(n16357), .B2(n14328), .C1(
        n16354), .C2(n12047), .ZN(n12563) );
  AOI221_X1 U4911 ( .B1(\registers[12][31] ), .B2(n16411), .C1(
        \registers[17][31] ), .C2(n16408), .A(n12539), .ZN(n12536) );
  OAI22_X1 U4912 ( .A1(n16405), .A2(n15071), .B1(n16402), .B2(n14425), .ZN(
        n12539) );
  AOI221_X1 U4913 ( .B1(\registers[56][31] ), .B2(n16267), .C1(
        \registers[60][31] ), .C2(n16264), .A(n12614), .ZN(n12611) );
  OAI222_X1 U4914 ( .A1(n16261), .A2(n14535), .B1(n16258), .B2(n12049), .C1(
        n16255), .C2(n15034), .ZN(n12614) );
  AOI221_X1 U4915 ( .B1(\registers[2][0] ), .B2(n16616), .C1(
        \registers[29][0] ), .C2(n16613), .A(n12461), .ZN(n12460) );
  OAI222_X1 U4916 ( .A1(n16610), .A2(n15004), .B1(n16607), .B2(n14300), .C1(
        n16604), .C2(n12018), .ZN(n12461) );
  AOI221_X1 U4917 ( .B1(\registers[56][0] ), .B2(n16517), .C1(
        \registers[60][0] ), .C2(n16514), .A(n12487), .ZN(n12486) );
  OAI222_X1 U4918 ( .A1(n16511), .A2(n14573), .B1(n16508), .B2(n12055), .C1(
        n16505), .C2(n15245), .ZN(n12487) );
  AOI221_X1 U4919 ( .B1(\registers[2][1] ), .B2(n16616), .C1(
        \registers[29][1] ), .C2(n16613), .A(n12281), .ZN(n12280) );
  OAI222_X1 U4920 ( .A1(n16610), .A2(n15005), .B1(n16607), .B2(n14301), .C1(
        n16604), .C2(n12019), .ZN(n12281) );
  AOI221_X1 U4921 ( .B1(\registers[2][2] ), .B2(n16616), .C1(
        \registers[29][2] ), .C2(n16613), .A(n12128), .ZN(n12127) );
  OAI222_X1 U4922 ( .A1(n16610), .A2(n15006), .B1(n16607), .B2(n14302), .C1(
        n16604), .C2(n12020), .ZN(n12128) );
  AOI221_X1 U4923 ( .B1(\registers[2][3] ), .B2(n16616), .C1(
        \registers[29][3] ), .C2(n16613), .A(n11975), .ZN(n11974) );
  OAI222_X1 U4924 ( .A1(n16610), .A2(n14989), .B1(n16607), .B2(n14282), .C1(
        n16604), .C2(n12016), .ZN(n11975) );
  AOI221_X1 U4925 ( .B1(\registers[2][4] ), .B2(n16616), .C1(
        \registers[29][4] ), .C2(n16613), .A(n11822), .ZN(n11821) );
  OAI222_X1 U4926 ( .A1(n16610), .A2(n14990), .B1(n16607), .B2(n14283), .C1(
        n16604), .C2(n12017), .ZN(n11822) );
  AOI221_X1 U4927 ( .B1(\registers[56][4] ), .B2(n16517), .C1(
        \registers[60][4] ), .C2(n16514), .A(n11838), .ZN(n11837) );
  OAI222_X1 U4928 ( .A1(n16511), .A2(n14538), .B1(n16508), .B2(n12050), .C1(
        n16505), .C2(n15241), .ZN(n11838) );
  AOI221_X1 U4929 ( .B1(\registers[2][5] ), .B2(n16616), .C1(
        \registers[29][5] ), .C2(n16613), .A(n11779), .ZN(n11778) );
  OAI222_X1 U4930 ( .A1(n16610), .A2(n15007), .B1(n16607), .B2(n14303), .C1(
        n16604), .C2(n12021), .ZN(n11779) );
  AOI221_X1 U4931 ( .B1(\registers[56][5] ), .B2(n16517), .C1(
        \registers[60][5] ), .C2(n16514), .A(n11795), .ZN(n11794) );
  OAI222_X1 U4932 ( .A1(n16511), .A2(n14539), .B1(n16508), .B2(n12051), .C1(
        n16505), .C2(n15242), .ZN(n11795) );
  AOI221_X1 U4933 ( .B1(\registers[2][6] ), .B2(n16616), .C1(
        \registers[29][6] ), .C2(n16613), .A(n11736), .ZN(n11735) );
  OAI222_X1 U4934 ( .A1(n16610), .A2(n15008), .B1(n16607), .B2(n14304), .C1(
        n16604), .C2(n12022), .ZN(n11736) );
  AOI221_X1 U4935 ( .B1(\registers[56][6] ), .B2(n16517), .C1(
        \registers[60][6] ), .C2(n16514), .A(n11752), .ZN(n11751) );
  OAI222_X1 U4936 ( .A1(n16511), .A2(n14574), .B1(n16508), .B2(n12056), .C1(
        n16505), .C2(n15246), .ZN(n11752) );
  AOI221_X1 U4937 ( .B1(\registers[2][7] ), .B2(n16616), .C1(
        \registers[29][7] ), .C2(n16613), .A(n11693), .ZN(n11692) );
  OAI222_X1 U4938 ( .A1(n16610), .A2(n15009), .B1(n16607), .B2(n14305), .C1(
        n16604), .C2(n12023), .ZN(n11693) );
  AOI221_X1 U4939 ( .B1(\registers[56][7] ), .B2(n16517), .C1(
        \registers[60][7] ), .C2(n16514), .A(n11709), .ZN(n11708) );
  OAI222_X1 U4940 ( .A1(n16511), .A2(n14575), .B1(n16508), .B2(n12057), .C1(
        n16505), .C2(n15247), .ZN(n11709) );
  AOI221_X1 U4941 ( .B1(\registers[2][8] ), .B2(n16616), .C1(
        \registers[29][8] ), .C2(n16613), .A(n11650), .ZN(n11649) );
  OAI222_X1 U4942 ( .A1(n16610), .A2(n15010), .B1(n16607), .B2(n14306), .C1(
        n16604), .C2(n12024), .ZN(n11650) );
  AOI221_X1 U4943 ( .B1(\registers[56][8] ), .B2(n16517), .C1(
        \registers[60][8] ), .C2(n16514), .A(n11666), .ZN(n11665) );
  OAI222_X1 U4944 ( .A1(n16511), .A2(n14576), .B1(n16508), .B2(n12058), .C1(
        n16505), .C2(n15248), .ZN(n11666) );
  AOI221_X1 U4945 ( .B1(\registers[2][9] ), .B2(n16616), .C1(
        \registers[29][9] ), .C2(n16613), .A(n11607), .ZN(n11606) );
  OAI222_X1 U4946 ( .A1(n16610), .A2(n15011), .B1(n16607), .B2(n14307), .C1(
        n16604), .C2(n12025), .ZN(n11607) );
  AOI221_X1 U4947 ( .B1(\registers[56][9] ), .B2(n16517), .C1(
        \registers[60][9] ), .C2(n16514), .A(n11623), .ZN(n11622) );
  OAI222_X1 U4948 ( .A1(n16511), .A2(n14577), .B1(n16508), .B2(n12059), .C1(
        n16505), .C2(n15249), .ZN(n11623) );
  AOI221_X1 U4949 ( .B1(\registers[2][10] ), .B2(n16616), .C1(
        \registers[29][10] ), .C2(n16613), .A(n11564), .ZN(n11563) );
  OAI222_X1 U4950 ( .A1(n16610), .A2(n15012), .B1(n16607), .B2(n14308), .C1(
        n16604), .C2(n12026), .ZN(n11564) );
  AOI221_X1 U4951 ( .B1(\registers[56][10] ), .B2(n16517), .C1(
        \registers[60][10] ), .C2(n16514), .A(n11580), .ZN(n11579) );
  OAI222_X1 U4952 ( .A1(n16511), .A2(n14578), .B1(n16508), .B2(n12060), .C1(
        n16505), .C2(n15250), .ZN(n11580) );
  AOI221_X1 U4953 ( .B1(\registers[2][11] ), .B2(n16616), .C1(
        \registers[29][11] ), .C2(n16613), .A(n11521), .ZN(n11520) );
  OAI222_X1 U4954 ( .A1(n16610), .A2(n15013), .B1(n16607), .B2(n14309), .C1(
        n16604), .C2(n12027), .ZN(n11521) );
  AOI221_X1 U4955 ( .B1(\registers[56][11] ), .B2(n16517), .C1(
        \registers[60][11] ), .C2(n16514), .A(n11537), .ZN(n11536) );
  OAI222_X1 U4956 ( .A1(n16511), .A2(n14579), .B1(n16508), .B2(n12098), .C1(
        n16505), .C2(n15251), .ZN(n11537) );
  AOI221_X1 U4957 ( .B1(\registers[2][12] ), .B2(n16617), .C1(
        \registers[29][12] ), .C2(n16614), .A(n11478), .ZN(n11477) );
  OAI222_X1 U4958 ( .A1(n16611), .A2(n15014), .B1(n16608), .B2(n14310), .C1(
        n16605), .C2(n12028), .ZN(n11478) );
  AOI221_X1 U4959 ( .B1(\registers[56][12] ), .B2(n16518), .C1(
        \registers[60][12] ), .C2(n16515), .A(n11494), .ZN(n11493) );
  OAI222_X1 U4960 ( .A1(n16512), .A2(n14580), .B1(n16509), .B2(n12099), .C1(
        n16506), .C2(n15252), .ZN(n11494) );
  AOI221_X1 U4961 ( .B1(\registers[2][13] ), .B2(n16617), .C1(
        \registers[29][13] ), .C2(n16614), .A(n11434), .ZN(n11433) );
  OAI222_X1 U4962 ( .A1(n16611), .A2(n15015), .B1(n16608), .B2(n14311), .C1(
        n16605), .C2(n12030), .ZN(n11434) );
  AOI221_X1 U4963 ( .B1(\registers[56][13] ), .B2(n16518), .C1(
        \registers[60][13] ), .C2(n16515), .A(n11450), .ZN(n11449) );
  OAI222_X1 U4964 ( .A1(n16512), .A2(n14581), .B1(n16509), .B2(n12100), .C1(
        n16506), .C2(n15253), .ZN(n11450) );
  AOI221_X1 U4965 ( .B1(\registers[2][14] ), .B2(n16617), .C1(
        \registers[29][14] ), .C2(n16614), .A(n11391), .ZN(n11390) );
  OAI222_X1 U4966 ( .A1(n16611), .A2(n15016), .B1(n16608), .B2(n14312), .C1(
        n16605), .C2(n12031), .ZN(n11391) );
  AOI221_X1 U4967 ( .B1(\registers[56][14] ), .B2(n16518), .C1(
        \registers[60][14] ), .C2(n16515), .A(n11407), .ZN(n11406) );
  OAI222_X1 U4968 ( .A1(n16512), .A2(n14582), .B1(n16509), .B2(n12101), .C1(
        n16506), .C2(n15254), .ZN(n11407) );
  AOI221_X1 U4969 ( .B1(\registers[2][15] ), .B2(n16617), .C1(
        \registers[29][15] ), .C2(n16614), .A(n11348), .ZN(n11347) );
  OAI222_X1 U4970 ( .A1(n16611), .A2(n15017), .B1(n16608), .B2(n14313), .C1(
        n16605), .C2(n12032), .ZN(n11348) );
  AOI221_X1 U4971 ( .B1(\registers[56][15] ), .B2(n16518), .C1(
        \registers[60][15] ), .C2(n16515), .A(n11364), .ZN(n11363) );
  OAI222_X1 U4972 ( .A1(n16512), .A2(n14583), .B1(n16509), .B2(n12102), .C1(
        n16506), .C2(n15255), .ZN(n11364) );
  AOI221_X1 U4973 ( .B1(\registers[2][16] ), .B2(n16617), .C1(
        \registers[29][16] ), .C2(n16614), .A(n11305), .ZN(n11304) );
  OAI222_X1 U4974 ( .A1(n16611), .A2(n15018), .B1(n16608), .B2(n14314), .C1(
        n16605), .C2(n12033), .ZN(n11305) );
  AOI221_X1 U4975 ( .B1(\registers[56][16] ), .B2(n16518), .C1(
        \registers[60][16] ), .C2(n16515), .A(n11321), .ZN(n11320) );
  OAI222_X1 U4976 ( .A1(n16512), .A2(n14584), .B1(n16509), .B2(n12103), .C1(
        n16506), .C2(n15256), .ZN(n11321) );
  AOI221_X1 U4977 ( .B1(\registers[2][17] ), .B2(n16617), .C1(
        \registers[29][17] ), .C2(n16614), .A(n11262), .ZN(n11261) );
  OAI222_X1 U4978 ( .A1(n16611), .A2(n15019), .B1(n16608), .B2(n14315), .C1(
        n16605), .C2(n12034), .ZN(n11262) );
  AOI221_X1 U4979 ( .B1(\registers[56][17] ), .B2(n16518), .C1(
        \registers[60][17] ), .C2(n16515), .A(n11278), .ZN(n11277) );
  OAI222_X1 U4980 ( .A1(n16512), .A2(n14585), .B1(n16509), .B2(n12104), .C1(
        n16506), .C2(n15257), .ZN(n11278) );
  AOI221_X1 U4981 ( .B1(\registers[2][18] ), .B2(n16617), .C1(
        \registers[29][18] ), .C2(n16614), .A(n11219), .ZN(n11218) );
  OAI222_X1 U4982 ( .A1(n16611), .A2(n15020), .B1(n16608), .B2(n14316), .C1(
        n16605), .C2(n12035), .ZN(n11219) );
  AOI221_X1 U4983 ( .B1(\registers[56][18] ), .B2(n16518), .C1(
        \registers[60][18] ), .C2(n16515), .A(n11235), .ZN(n11234) );
  OAI222_X1 U4984 ( .A1(n16512), .A2(n14586), .B1(n16509), .B2(n12105), .C1(
        n16506), .C2(n15258), .ZN(n11235) );
  AOI221_X1 U4985 ( .B1(\registers[2][19] ), .B2(n16617), .C1(
        \registers[29][19] ), .C2(n16614), .A(n11176), .ZN(n11175) );
  OAI222_X1 U4986 ( .A1(n16611), .A2(n15021), .B1(n16608), .B2(n14317), .C1(
        n16605), .C2(n12036), .ZN(n11176) );
  AOI221_X1 U4987 ( .B1(\registers[56][19] ), .B2(n16518), .C1(
        \registers[60][19] ), .C2(n16515), .A(n11192), .ZN(n11191) );
  OAI222_X1 U4988 ( .A1(n16512), .A2(n14587), .B1(n16509), .B2(n12148), .C1(
        n16506), .C2(n15259), .ZN(n11192) );
  AOI221_X1 U4989 ( .B1(\registers[2][20] ), .B2(n16617), .C1(
        \registers[29][20] ), .C2(n16614), .A(n11133), .ZN(n11132) );
  OAI222_X1 U4990 ( .A1(n16611), .A2(n15022), .B1(n16608), .B2(n14318), .C1(
        n16605), .C2(n12037), .ZN(n11133) );
  AOI221_X1 U4991 ( .B1(\registers[56][20] ), .B2(n16518), .C1(
        \registers[60][20] ), .C2(n16515), .A(n11149), .ZN(n11148) );
  OAI222_X1 U4992 ( .A1(n16512), .A2(n14588), .B1(n16509), .B2(n12150), .C1(
        n16506), .C2(n15260), .ZN(n11149) );
  AOI221_X1 U4993 ( .B1(\registers[2][21] ), .B2(n16617), .C1(
        \registers[29][21] ), .C2(n16614), .A(n11090), .ZN(n11089) );
  OAI222_X1 U4994 ( .A1(n16611), .A2(n15023), .B1(n16608), .B2(n14319), .C1(
        n16605), .C2(n12038), .ZN(n11090) );
  AOI221_X1 U4995 ( .B1(\registers[56][21] ), .B2(n16518), .C1(
        \registers[60][21] ), .C2(n16515), .A(n11106), .ZN(n11105) );
  OAI222_X1 U4996 ( .A1(n16512), .A2(n14589), .B1(n16509), .B2(n12151), .C1(
        n16506), .C2(n15261), .ZN(n11106) );
  AOI221_X1 U4997 ( .B1(\registers[2][22] ), .B2(n16617), .C1(
        \registers[29][22] ), .C2(n16614), .A(n11047), .ZN(n11046) );
  OAI222_X1 U4998 ( .A1(n16611), .A2(n15024), .B1(n16608), .B2(n14320), .C1(
        n16605), .C2(n12039), .ZN(n11047) );
  AOI221_X1 U4999 ( .B1(\registers[56][22] ), .B2(n16518), .C1(
        \registers[60][22] ), .C2(n16515), .A(n11063), .ZN(n11062) );
  OAI222_X1 U5000 ( .A1(n16512), .A2(n14590), .B1(n16509), .B2(n12152), .C1(
        n16506), .C2(n15262), .ZN(n11063) );
  AOI221_X1 U5001 ( .B1(\registers[2][23] ), .B2(n16617), .C1(
        \registers[29][23] ), .C2(n16614), .A(n11004), .ZN(n11003) );
  OAI222_X1 U5002 ( .A1(n16611), .A2(n15025), .B1(n16608), .B2(n14321), .C1(
        n16605), .C2(n12040), .ZN(n11004) );
  AOI221_X1 U5003 ( .B1(\registers[56][23] ), .B2(n16518), .C1(
        \registers[60][23] ), .C2(n16515), .A(n11020), .ZN(n11019) );
  OAI222_X1 U5004 ( .A1(n16512), .A2(n14591), .B1(n16509), .B2(n12153), .C1(
        n16506), .C2(n15263), .ZN(n11020) );
  AOI221_X1 U5005 ( .B1(\registers[2][24] ), .B2(n16618), .C1(
        \registers[29][24] ), .C2(n16615), .A(n10961), .ZN(n10960) );
  OAI222_X1 U5006 ( .A1(n16612), .A2(n15026), .B1(n16609), .B2(n14322), .C1(
        n16606), .C2(n12041), .ZN(n10961) );
  AOI221_X1 U5007 ( .B1(\registers[12][24] ), .B2(n16663), .C1(
        \registers[15][24] ), .C2(n16660), .A(n10953), .ZN(n10952) );
  OAI22_X1 U5008 ( .A1(n16657), .A2(n15065), .B1(n16654), .B2(n14419), .ZN(
        n10953) );
  AOI221_X1 U5009 ( .B1(net227344), .B2(n16567), .C1(\registers[44][24] ), 
        .C2(n16564), .A(n10969), .ZN(n10968) );
  OAI22_X1 U5010 ( .A1(n16561), .A2(n15144), .B1(n16558), .B2(n14527), .ZN(
        n10969) );
  AOI221_X1 U5011 ( .B1(\registers[56][24] ), .B2(n16519), .C1(
        \registers[60][24] ), .C2(n16516), .A(n10977), .ZN(n10976) );
  OAI222_X1 U5012 ( .A1(n16513), .A2(n14592), .B1(n16510), .B2(n12154), .C1(
        n16507), .C2(n15264), .ZN(n10977) );
  AOI221_X1 U5013 ( .B1(\registers[2][25] ), .B2(n16618), .C1(
        \registers[29][25] ), .C2(n16615), .A(n10918), .ZN(n10917) );
  OAI222_X1 U5014 ( .A1(n16612), .A2(n15027), .B1(n16609), .B2(n14323), .C1(
        n16606), .C2(n12042), .ZN(n10918) );
  AOI221_X1 U5015 ( .B1(\registers[12][25] ), .B2(n16663), .C1(
        \registers[15][25] ), .C2(n16660), .A(n10910), .ZN(n10909) );
  OAI22_X1 U5016 ( .A1(n16657), .A2(n15066), .B1(n16654), .B2(n14420), .ZN(
        n10910) );
  AOI221_X1 U5017 ( .B1(net227362), .B2(n16567), .C1(\registers[44][25] ), 
        .C2(n16564), .A(n10926), .ZN(n10925) );
  OAI22_X1 U5018 ( .A1(n16561), .A2(n15145), .B1(n16558), .B2(n14528), .ZN(
        n10926) );
  AOI221_X1 U5019 ( .B1(\registers[56][25] ), .B2(n16519), .C1(
        \registers[60][25] ), .C2(n16516), .A(n10934), .ZN(n10933) );
  OAI222_X1 U5020 ( .A1(n16513), .A2(n14593), .B1(n16510), .B2(n12155), .C1(
        n16507), .C2(n15265), .ZN(n10934) );
  AOI221_X1 U5021 ( .B1(\registers[2][26] ), .B2(n16618), .C1(
        \registers[29][26] ), .C2(n16615), .A(n10875), .ZN(n10874) );
  OAI222_X1 U5022 ( .A1(n16612), .A2(n15028), .B1(n16609), .B2(n14324), .C1(
        n16606), .C2(n12043), .ZN(n10875) );
  AOI221_X1 U5023 ( .B1(\registers[12][26] ), .B2(n16663), .C1(
        \registers[15][26] ), .C2(n16660), .A(n10867), .ZN(n10866) );
  OAI22_X1 U5024 ( .A1(n16657), .A2(n15067), .B1(n16654), .B2(n14421), .ZN(
        n10867) );
  AOI221_X1 U5025 ( .B1(net227380), .B2(n16567), .C1(\registers[44][26] ), 
        .C2(n16564), .A(n10883), .ZN(n10882) );
  OAI22_X1 U5026 ( .A1(n16561), .A2(n15146), .B1(n16558), .B2(n14529), .ZN(
        n10883) );
  AOI221_X1 U5027 ( .B1(\registers[56][26] ), .B2(n16519), .C1(
        \registers[60][26] ), .C2(n16516), .A(n10891), .ZN(n10890) );
  OAI222_X1 U5028 ( .A1(n16513), .A2(n14594), .B1(n16510), .B2(n12156), .C1(
        n16507), .C2(n15266), .ZN(n10891) );
  AOI221_X1 U5029 ( .B1(\registers[2][27] ), .B2(n16618), .C1(
        \registers[29][27] ), .C2(n16615), .A(n10832), .ZN(n10831) );
  OAI222_X1 U5030 ( .A1(n16612), .A2(n15029), .B1(n16609), .B2(n14325), .C1(
        n16606), .C2(n12044), .ZN(n10832) );
  AOI221_X1 U5031 ( .B1(\registers[12][27] ), .B2(n16663), .C1(
        \registers[15][27] ), .C2(n16660), .A(n10824), .ZN(n10823) );
  OAI22_X1 U5032 ( .A1(n16657), .A2(n15068), .B1(n16654), .B2(n14422), .ZN(
        n10824) );
  AOI221_X1 U5033 ( .B1(net227398), .B2(n16567), .C1(\registers[44][27] ), 
        .C2(n16564), .A(n10840), .ZN(n10839) );
  OAI22_X1 U5034 ( .A1(n16561), .A2(n15147), .B1(n16558), .B2(n14530), .ZN(
        n10840) );
  AOI221_X1 U5035 ( .B1(\registers[56][27] ), .B2(n16519), .C1(
        \registers[60][27] ), .C2(n16516), .A(n10848), .ZN(n10847) );
  OAI222_X1 U5036 ( .A1(n16513), .A2(n14595), .B1(n16510), .B2(n12157), .C1(
        n16507), .C2(n15267), .ZN(n10848) );
  AOI221_X1 U5037 ( .B1(\registers[2][28] ), .B2(n16618), .C1(
        \registers[29][28] ), .C2(n16615), .A(n10789), .ZN(n10788) );
  OAI222_X1 U5038 ( .A1(n16612), .A2(n15030), .B1(n16609), .B2(n14326), .C1(
        n16606), .C2(n12045), .ZN(n10789) );
  AOI221_X1 U5039 ( .B1(\registers[12][28] ), .B2(n16663), .C1(
        \registers[15][28] ), .C2(n16660), .A(n10781), .ZN(n10780) );
  OAI22_X1 U5040 ( .A1(n16657), .A2(n15069), .B1(n16654), .B2(n14423), .ZN(
        n10781) );
  AOI221_X1 U5041 ( .B1(net227416), .B2(n16567), .C1(\registers[44][28] ), 
        .C2(n16564), .A(n10797), .ZN(n10796) );
  OAI22_X1 U5042 ( .A1(n16561), .A2(n15148), .B1(n16558), .B2(n14531), .ZN(
        n10797) );
  AOI221_X1 U5043 ( .B1(\registers[56][28] ), .B2(n16519), .C1(
        \registers[60][28] ), .C2(n16516), .A(n10805), .ZN(n10804) );
  OAI222_X1 U5044 ( .A1(n16513), .A2(n14596), .B1(n16510), .B2(n12158), .C1(
        n16507), .C2(n15268), .ZN(n10805) );
  AOI221_X1 U5045 ( .B1(\registers[2][29] ), .B2(n16618), .C1(
        \registers[29][29] ), .C2(n16615), .A(n10746), .ZN(n10745) );
  OAI222_X1 U5046 ( .A1(n16612), .A2(n15031), .B1(n16609), .B2(n14327), .C1(
        n16606), .C2(n12046), .ZN(n10746) );
  AOI221_X1 U5047 ( .B1(\registers[12][29] ), .B2(n16663), .C1(
        \registers[15][29] ), .C2(n16660), .A(n10738), .ZN(n10737) );
  OAI22_X1 U5048 ( .A1(n16657), .A2(n15070), .B1(n16654), .B2(n14424), .ZN(
        n10738) );
  AOI221_X1 U5049 ( .B1(net227434), .B2(n16567), .C1(\registers[44][29] ), 
        .C2(n16564), .A(n10754), .ZN(n10753) );
  OAI22_X1 U5050 ( .A1(n16561), .A2(n15149), .B1(n16558), .B2(n14532), .ZN(
        n10754) );
  AOI221_X1 U5051 ( .B1(\registers[56][29] ), .B2(n16519), .C1(
        \registers[60][29] ), .C2(n16516), .A(n10762), .ZN(n10761) );
  OAI222_X1 U5052 ( .A1(n16513), .A2(n14597), .B1(n16510), .B2(n12159), .C1(
        n16507), .C2(n15269), .ZN(n10762) );
  AOI221_X1 U5053 ( .B1(\registers[2][30] ), .B2(n16618), .C1(
        \registers[29][30] ), .C2(n16615), .A(n10691), .ZN(n10690) );
  OAI222_X1 U5054 ( .A1(n16612), .A2(n14857), .B1(n16609), .B2(n14054), .C1(
        n16606), .C2(n11904), .ZN(n10691) );
  AOI221_X1 U5055 ( .B1(\registers[12][30] ), .B2(n16663), .C1(
        \registers[15][30] ), .C2(n16660), .A(n10679), .ZN(n10678) );
  OAI22_X1 U5056 ( .A1(n16657), .A2(n14870), .B1(n16654), .B2(n14060), .ZN(
        n10679) );
  AOI221_X1 U5057 ( .B1(net227452), .B2(n16567), .C1(\registers[44][30] ), 
        .C2(n16564), .A(n10704), .ZN(n10703) );
  OAI22_X1 U5058 ( .A1(n16561), .A2(n14871), .B1(n16558), .B2(n14069), .ZN(
        n10704) );
  AOI221_X1 U5059 ( .B1(\registers[56][30] ), .B2(n16519), .C1(
        \registers[60][30] ), .C2(n16516), .A(n10717), .ZN(n10716) );
  OAI222_X1 U5060 ( .A1(n16513), .A2(n14534), .B1(n16510), .B2(n12048), .C1(
        n16507), .C2(n15033), .ZN(n10717) );
  AOI221_X1 U5061 ( .B1(\registers[2][31] ), .B2(n16618), .C1(
        \registers[29][31] ), .C2(n16615), .A(n10568), .ZN(n10565) );
  OAI222_X1 U5062 ( .A1(n16612), .A2(n15032), .B1(n16609), .B2(n14328), .C1(
        n16606), .C2(n12047), .ZN(n10568) );
  AOI221_X1 U5063 ( .B1(\registers[12][31] ), .B2(n16663), .C1(
        \registers[15][31] ), .C2(n16660), .A(n10537), .ZN(n10534) );
  OAI22_X1 U5064 ( .A1(n16657), .A2(n15071), .B1(n16654), .B2(n14425), .ZN(
        n10537) );
  AOI221_X1 U5065 ( .B1(net227470), .B2(n16567), .C1(\registers[44][31] ), 
        .C2(n16564), .A(n10602), .ZN(n10599) );
  OAI22_X1 U5066 ( .A1(n16561), .A2(n15150), .B1(n16558), .B2(n14533), .ZN(
        n10602) );
  AOI221_X1 U5067 ( .B1(\registers[56][31] ), .B2(n16519), .C1(
        \registers[60][31] ), .C2(n16516), .A(n10634), .ZN(n10631) );
  OAI222_X1 U5068 ( .A1(n16513), .A2(n14535), .B1(n16510), .B2(n12049), .C1(
        n16507), .C2(n15034), .ZN(n10634) );
  AOI221_X1 U5069 ( .B1(\registers[37][23] ), .B2(n17819), .C1(
        \registers[0][23] ), .C2(n17816), .A(n5281), .ZN(n5280) );
  OAI22_X1 U5070 ( .A1(n17813), .A2(n15662), .B1(n17810), .B2(n14700), .ZN(
        n5281) );
  AOI221_X1 U5071 ( .B1(\registers[37][24] ), .B2(n17819), .C1(
        \registers[0][24] ), .C2(n17816), .A(n5116), .ZN(n5115) );
  OAI22_X1 U5072 ( .A1(n17813), .A2(n15663), .B1(n17810), .B2(n14701), .ZN(
        n5116) );
  AOI221_X1 U5073 ( .B1(\registers[37][25] ), .B2(n17819), .C1(
        \registers[0][25] ), .C2(n17816), .A(n5002), .ZN(n5001) );
  OAI22_X1 U5074 ( .A1(n17813), .A2(n15664), .B1(n17810), .B2(n14702), .ZN(
        n5002) );
  AOI221_X1 U5075 ( .B1(\registers[56][26] ), .B2(n17675), .C1(
        \registers[55][26] ), .C2(n17672), .A(n4910), .ZN(n4909) );
  OAI22_X1 U5076 ( .A1(n17669), .A2(n15428), .B1(n17666), .B2(n14703), .ZN(
        n4910) );
  AOI221_X1 U5077 ( .B1(\registers[37][26] ), .B2(n17819), .C1(
        \registers[0][26] ), .C2(n17816), .A(n4880), .ZN(n4879) );
  OAI22_X1 U5078 ( .A1(n17813), .A2(n15665), .B1(n17810), .B2(n14704), .ZN(
        n4880) );
  AOI221_X1 U5079 ( .B1(\registers[56][27] ), .B2(n17675), .C1(
        \registers[55][27] ), .C2(n17672), .A(n4779), .ZN(n4778) );
  OAI22_X1 U5080 ( .A1(n17669), .A2(n15429), .B1(n17666), .B2(n14705), .ZN(
        n4779) );
  AOI221_X1 U5081 ( .B1(\registers[37][27] ), .B2(n17819), .C1(
        \registers[0][27] ), .C2(n17816), .A(n4751), .ZN(n4750) );
  OAI22_X1 U5082 ( .A1(n17813), .A2(n15666), .B1(n17810), .B2(n14706), .ZN(
        n4751) );
  AOI221_X1 U5083 ( .B1(\registers[56][28] ), .B2(n17675), .C1(
        \registers[55][28] ), .C2(n17672), .A(n4650), .ZN(n4649) );
  OAI22_X1 U5084 ( .A1(n17669), .A2(n15430), .B1(n17666), .B2(n14707), .ZN(
        n4650) );
  AOI221_X1 U5085 ( .B1(\registers[37][28] ), .B2(n17819), .C1(
        \registers[0][28] ), .C2(n17816), .A(n4622), .ZN(n4621) );
  OAI22_X1 U5086 ( .A1(n17813), .A2(n15667), .B1(n17810), .B2(n14708), .ZN(
        n4622) );
  AOI221_X1 U5087 ( .B1(\registers[56][29] ), .B2(n17675), .C1(
        \registers[55][29] ), .C2(n17672), .A(n4521), .ZN(n4520) );
  OAI22_X1 U5088 ( .A1(n17669), .A2(n15431), .B1(n17666), .B2(n14709), .ZN(
        n4521) );
  AOI221_X1 U5089 ( .B1(\registers[37][29] ), .B2(n17819), .C1(
        \registers[0][29] ), .C2(n17816), .A(n4489), .ZN(n4488) );
  OAI22_X1 U5090 ( .A1(n17813), .A2(n15668), .B1(n17810), .B2(n14710), .ZN(
        n4489) );
  AOI221_X1 U5091 ( .B1(\registers[37][30] ), .B2(n17819), .C1(
        \registers[0][30] ), .C2(n17816), .A(n4109), .ZN(n4106) );
  OAI22_X1 U5092 ( .A1(n17813), .A2(n15280), .B1(n17810), .B2(n14629), .ZN(
        n4109) );
  AOI221_X1 U5093 ( .B1(\registers[12][0] ), .B2(n16409), .C1(
        \registers[17][0] ), .C2(n16406), .A(n13916), .ZN(n13915) );
  OAI22_X1 U5094 ( .A1(n16403), .A2(n15072), .B1(n16400), .B2(n14426), .ZN(
        n13916) );
  AOI221_X1 U5095 ( .B1(net226850), .B2(n16313), .C1(\registers[44][0] ), .C2(
        n16310), .A(n13952), .ZN(n13951) );
  OAI22_X1 U5096 ( .A1(n16307), .A2(n15073), .B1(n16304), .B2(n14427), .ZN(
        n13952) );
  AOI221_X1 U5097 ( .B1(\registers[12][1] ), .B2(n16409), .C1(
        \registers[17][1] ), .C2(n16406), .A(n13869), .ZN(n13868) );
  OAI22_X1 U5098 ( .A1(n16403), .A2(n15074), .B1(n16400), .B2(n14428), .ZN(
        n13869) );
  AOI221_X1 U5099 ( .B1(net226870), .B2(n16313), .C1(\registers[44][1] ), .C2(
        n16310), .A(n13885), .ZN(n13884) );
  OAI22_X1 U5100 ( .A1(n16307), .A2(n15075), .B1(n16304), .B2(n14429), .ZN(
        n13885) );
  AOI221_X1 U5101 ( .B1(\registers[12][2] ), .B2(n16409), .C1(
        \registers[17][2] ), .C2(n16406), .A(n13827), .ZN(n13826) );
  OAI22_X1 U5102 ( .A1(n16403), .A2(n15076), .B1(n16400), .B2(n14430), .ZN(
        n13827) );
  AOI221_X1 U5103 ( .B1(net226883), .B2(n16313), .C1(\registers[44][2] ), .C2(
        n16310), .A(n13843), .ZN(n13842) );
  OAI22_X1 U5104 ( .A1(n16307), .A2(n15077), .B1(n16304), .B2(n14431), .ZN(
        n13843) );
  AOI221_X1 U5105 ( .B1(\registers[12][3] ), .B2(n16409), .C1(
        \registers[17][3] ), .C2(n16406), .A(n13785), .ZN(n13784) );
  OAI22_X1 U5106 ( .A1(n16403), .A2(n14994), .B1(n16400), .B2(n14291), .ZN(
        n13785) );
  AOI221_X1 U5107 ( .B1(net226903), .B2(n16313), .C1(\registers[44][3] ), .C2(
        n16310), .A(n13801), .ZN(n13800) );
  OAI22_X1 U5108 ( .A1(n16307), .A2(n14995), .B1(n16304), .B2(n14292), .ZN(
        n13801) );
  AOI221_X1 U5109 ( .B1(\registers[12][4] ), .B2(n16409), .C1(
        \registers[17][4] ), .C2(n16406), .A(n13743), .ZN(n13742) );
  OAI22_X1 U5110 ( .A1(n16403), .A2(n15078), .B1(n16400), .B2(n14432), .ZN(
        n13743) );
  AOI221_X1 U5111 ( .B1(net226976), .B2(n16313), .C1(\registers[44][4] ), .C2(
        n16310), .A(n13759), .ZN(n13758) );
  OAI22_X1 U5112 ( .A1(n16307), .A2(n15079), .B1(n16304), .B2(n14433), .ZN(
        n13759) );
  AOI221_X1 U5113 ( .B1(\registers[12][5] ), .B2(n16409), .C1(
        \registers[17][5] ), .C2(n16406), .A(n13701), .ZN(n13700) );
  OAI22_X1 U5114 ( .A1(n16403), .A2(n15080), .B1(n16400), .B2(n14434), .ZN(
        n13701) );
  AOI221_X1 U5115 ( .B1(net226996), .B2(n16313), .C1(\registers[44][5] ), .C2(
        n16310), .A(n13717), .ZN(n13716) );
  OAI22_X1 U5116 ( .A1(n16307), .A2(n14996), .B1(n16304), .B2(n14293), .ZN(
        n13717) );
  AOI221_X1 U5117 ( .B1(\registers[12][6] ), .B2(n16409), .C1(
        \registers[17][6] ), .C2(n16406), .A(n13659), .ZN(n13658) );
  OAI22_X1 U5118 ( .A1(n16403), .A2(n15081), .B1(n16400), .B2(n14435), .ZN(
        n13659) );
  AOI221_X1 U5119 ( .B1(net227020), .B2(n16313), .C1(\registers[44][6] ), .C2(
        n16310), .A(n13675), .ZN(n13674) );
  OAI22_X1 U5120 ( .A1(n16307), .A2(n15082), .B1(n16304), .B2(n14436), .ZN(
        n13675) );
  AOI221_X1 U5121 ( .B1(\registers[12][7] ), .B2(n16409), .C1(
        \registers[17][7] ), .C2(n16406), .A(n13617), .ZN(n13616) );
  OAI22_X1 U5122 ( .A1(n16403), .A2(n15083), .B1(n16400), .B2(n14437), .ZN(
        n13617) );
  AOI221_X1 U5123 ( .B1(net227038), .B2(n16313), .C1(\registers[44][7] ), .C2(
        n16310), .A(n13633), .ZN(n13632) );
  OAI22_X1 U5124 ( .A1(n16307), .A2(n15084), .B1(n16304), .B2(n14438), .ZN(
        n13633) );
  AOI221_X1 U5125 ( .B1(\registers[12][8] ), .B2(n16409), .C1(
        \registers[17][8] ), .C2(n16406), .A(n13575), .ZN(n13574) );
  OAI22_X1 U5126 ( .A1(n16403), .A2(n15085), .B1(n16400), .B2(n14439), .ZN(
        n13575) );
  AOI221_X1 U5127 ( .B1(net227056), .B2(n16313), .C1(\registers[44][8] ), .C2(
        n16310), .A(n13591), .ZN(n13590) );
  OAI22_X1 U5128 ( .A1(n16307), .A2(n15086), .B1(n16304), .B2(n14440), .ZN(
        n13591) );
  AOI221_X1 U5129 ( .B1(\registers[12][9] ), .B2(n16409), .C1(
        \registers[17][9] ), .C2(n16406), .A(n13533), .ZN(n13532) );
  OAI22_X1 U5130 ( .A1(n16403), .A2(n15087), .B1(n16400), .B2(n14441), .ZN(
        n13533) );
  AOI221_X1 U5131 ( .B1(net227074), .B2(n16313), .C1(\registers[44][9] ), .C2(
        n16310), .A(n13549), .ZN(n13548) );
  OAI22_X1 U5132 ( .A1(n16307), .A2(n15088), .B1(n16304), .B2(n14442), .ZN(
        n13549) );
  AOI221_X1 U5133 ( .B1(\registers[12][10] ), .B2(n16409), .C1(
        \registers[17][10] ), .C2(n16406), .A(n13491), .ZN(n13490) );
  OAI22_X1 U5134 ( .A1(n16403), .A2(n15089), .B1(n16400), .B2(n14443), .ZN(
        n13491) );
  AOI221_X1 U5135 ( .B1(net227092), .B2(n16313), .C1(\registers[44][10] ), 
        .C2(n16310), .A(n13507), .ZN(n13506) );
  OAI22_X1 U5136 ( .A1(n16307), .A2(n15090), .B1(n16304), .B2(n14444), .ZN(
        n13507) );
  AOI221_X1 U5137 ( .B1(\registers[12][11] ), .B2(n16409), .C1(
        \registers[17][11] ), .C2(n16406), .A(n13449), .ZN(n13448) );
  OAI22_X1 U5138 ( .A1(n16403), .A2(n15091), .B1(n16400), .B2(n14445), .ZN(
        n13449) );
  AOI221_X1 U5139 ( .B1(net227110), .B2(n16313), .C1(\registers[44][11] ), 
        .C2(n16310), .A(n13465), .ZN(n13464) );
  OAI22_X1 U5140 ( .A1(n16307), .A2(n15092), .B1(n16304), .B2(n14446), .ZN(
        n13465) );
  AOI221_X1 U5141 ( .B1(\registers[12][12] ), .B2(n16410), .C1(
        \registers[17][12] ), .C2(n16407), .A(n13407), .ZN(n13406) );
  OAI22_X1 U5142 ( .A1(n16404), .A2(n15093), .B1(n16401), .B2(n14447), .ZN(
        n13407) );
  AOI221_X1 U5143 ( .B1(net227128), .B2(n16314), .C1(\registers[44][12] ), 
        .C2(n16311), .A(n13423), .ZN(n13422) );
  OAI22_X1 U5144 ( .A1(n16308), .A2(n15094), .B1(n16305), .B2(n14448), .ZN(
        n13423) );
  AOI221_X1 U5145 ( .B1(\registers[12][13] ), .B2(n16410), .C1(
        \registers[17][13] ), .C2(n16407), .A(n13365), .ZN(n13364) );
  OAI22_X1 U5146 ( .A1(n16404), .A2(n15095), .B1(n16401), .B2(n14449), .ZN(
        n13365) );
  AOI221_X1 U5147 ( .B1(net227146), .B2(n16314), .C1(\registers[44][13] ), 
        .C2(n16311), .A(n13381), .ZN(n13380) );
  OAI22_X1 U5148 ( .A1(n16308), .A2(n15096), .B1(n16305), .B2(n14450), .ZN(
        n13381) );
  AOI221_X1 U5149 ( .B1(\registers[12][14] ), .B2(n16410), .C1(
        \registers[17][14] ), .C2(n16407), .A(n13323), .ZN(n13322) );
  OAI22_X1 U5150 ( .A1(n16404), .A2(n15097), .B1(n16401), .B2(n14451), .ZN(
        n13323) );
  AOI221_X1 U5151 ( .B1(net227164), .B2(n16314), .C1(\registers[44][14] ), 
        .C2(n16311), .A(n13339), .ZN(n13338) );
  OAI22_X1 U5152 ( .A1(n16308), .A2(n15098), .B1(n16305), .B2(n14452), .ZN(
        n13339) );
  AOI221_X1 U5153 ( .B1(\registers[12][15] ), .B2(n16410), .C1(
        \registers[17][15] ), .C2(n16407), .A(n13281), .ZN(n13280) );
  OAI22_X1 U5154 ( .A1(n16404), .A2(n15099), .B1(n16401), .B2(n14453), .ZN(
        n13281) );
  AOI221_X1 U5155 ( .B1(net227182), .B2(n16314), .C1(\registers[44][15] ), 
        .C2(n16311), .A(n13297), .ZN(n13296) );
  OAI22_X1 U5156 ( .A1(n16308), .A2(n15100), .B1(n16305), .B2(n14454), .ZN(
        n13297) );
  AOI221_X1 U5157 ( .B1(\registers[12][16] ), .B2(n16410), .C1(
        \registers[17][16] ), .C2(n16407), .A(n13239), .ZN(n13238) );
  OAI22_X1 U5158 ( .A1(n16404), .A2(n15101), .B1(n16401), .B2(n14455), .ZN(
        n13239) );
  AOI221_X1 U5159 ( .B1(net227200), .B2(n16314), .C1(\registers[44][16] ), 
        .C2(n16311), .A(n13255), .ZN(n13254) );
  OAI22_X1 U5160 ( .A1(n16308), .A2(n15102), .B1(n16305), .B2(n14456), .ZN(
        n13255) );
  AOI221_X1 U5161 ( .B1(\registers[12][17] ), .B2(n16410), .C1(
        \registers[17][17] ), .C2(n16407), .A(n13197), .ZN(n13196) );
  OAI22_X1 U5162 ( .A1(n16404), .A2(n15103), .B1(n16401), .B2(n14457), .ZN(
        n13197) );
  AOI221_X1 U5163 ( .B1(net227218), .B2(n16314), .C1(\registers[44][17] ), 
        .C2(n16311), .A(n13213), .ZN(n13212) );
  OAI22_X1 U5164 ( .A1(n16308), .A2(n15104), .B1(n16305), .B2(n14458), .ZN(
        n13213) );
  AOI221_X1 U5165 ( .B1(\registers[12][18] ), .B2(n16410), .C1(
        \registers[17][18] ), .C2(n16407), .A(n13155), .ZN(n13154) );
  OAI22_X1 U5166 ( .A1(n16404), .A2(n15105), .B1(n16401), .B2(n14459), .ZN(
        n13155) );
  AOI221_X1 U5167 ( .B1(net227236), .B2(n16314), .C1(\registers[44][18] ), 
        .C2(n16311), .A(n13171), .ZN(n13170) );
  OAI22_X1 U5168 ( .A1(n16308), .A2(n15106), .B1(n16305), .B2(n14460), .ZN(
        n13171) );
  AOI221_X1 U5169 ( .B1(\registers[12][19] ), .B2(n16410), .C1(
        \registers[17][19] ), .C2(n16407), .A(n13113), .ZN(n13112) );
  OAI22_X1 U5170 ( .A1(n16404), .A2(n15107), .B1(n16401), .B2(n14461), .ZN(
        n13113) );
  AOI221_X1 U5171 ( .B1(net227254), .B2(n16314), .C1(\registers[44][19] ), 
        .C2(n16311), .A(n13129), .ZN(n13128) );
  OAI22_X1 U5172 ( .A1(n16308), .A2(n15108), .B1(n16305), .B2(n14462), .ZN(
        n13129) );
  AOI221_X1 U5173 ( .B1(\registers[12][20] ), .B2(n16410), .C1(
        \registers[17][20] ), .C2(n16407), .A(n13071), .ZN(n13070) );
  OAI22_X1 U5174 ( .A1(n16404), .A2(n15109), .B1(n16401), .B2(n14463), .ZN(
        n13071) );
  AOI221_X1 U5175 ( .B1(net227272), .B2(n16314), .C1(\registers[44][20] ), 
        .C2(n16311), .A(n13087), .ZN(n13086) );
  OAI22_X1 U5176 ( .A1(n16308), .A2(n15110), .B1(n16305), .B2(n14464), .ZN(
        n13087) );
  AOI221_X1 U5177 ( .B1(\registers[12][21] ), .B2(n16410), .C1(
        \registers[17][21] ), .C2(n16407), .A(n13029), .ZN(n13028) );
  OAI22_X1 U5178 ( .A1(n16404), .A2(n15111), .B1(n16401), .B2(n14465), .ZN(
        n13029) );
  AOI221_X1 U5179 ( .B1(net227290), .B2(n16314), .C1(\registers[44][21] ), 
        .C2(n16311), .A(n13045), .ZN(n13044) );
  OAI22_X1 U5180 ( .A1(n16308), .A2(n15112), .B1(n16305), .B2(n14466), .ZN(
        n13045) );
  AOI221_X1 U5181 ( .B1(\registers[12][22] ), .B2(n16410), .C1(
        \registers[17][22] ), .C2(n16407), .A(n12987), .ZN(n12986) );
  OAI22_X1 U5182 ( .A1(n16404), .A2(n15113), .B1(n16401), .B2(n14467), .ZN(
        n12987) );
  AOI221_X1 U5183 ( .B1(net227308), .B2(n16314), .C1(\registers[44][22] ), 
        .C2(n16311), .A(n13003), .ZN(n13002) );
  OAI22_X1 U5184 ( .A1(n16308), .A2(n15114), .B1(n16305), .B2(n14468), .ZN(
        n13003) );
  AOI221_X1 U5185 ( .B1(\registers[12][23] ), .B2(n16410), .C1(
        \registers[17][23] ), .C2(n16407), .A(n12945), .ZN(n12944) );
  OAI22_X1 U5186 ( .A1(n16404), .A2(n15115), .B1(n16401), .B2(n14469), .ZN(
        n12945) );
  AOI221_X1 U5187 ( .B1(net227326), .B2(n16314), .C1(\registers[44][23] ), 
        .C2(n16311), .A(n12961), .ZN(n12960) );
  OAI22_X1 U5188 ( .A1(n16308), .A2(n15116), .B1(n16305), .B2(n14470), .ZN(
        n12961) );
  AOI221_X1 U5189 ( .B1(\registers[12][0] ), .B2(n16661), .C1(
        \registers[15][0] ), .C2(n16658), .A(n12435), .ZN(n12434) );
  OAI22_X1 U5190 ( .A1(n16655), .A2(n15072), .B1(n16652), .B2(n14426), .ZN(
        n12435) );
  AOI221_X1 U5191 ( .B1(net226850), .B2(n16565), .C1(\registers[44][0] ), .C2(
        n16562), .A(n12471), .ZN(n12470) );
  OAI22_X1 U5192 ( .A1(n16559), .A2(n15073), .B1(n16556), .B2(n14427), .ZN(
        n12471) );
  AOI221_X1 U5193 ( .B1(\registers[12][1] ), .B2(n16661), .C1(
        \registers[15][1] ), .C2(n16658), .A(n12273), .ZN(n12272) );
  OAI22_X1 U5194 ( .A1(n16655), .A2(n15074), .B1(n16652), .B2(n14428), .ZN(
        n12273) );
  AOI221_X1 U5195 ( .B1(net226870), .B2(n16565), .C1(\registers[44][1] ), .C2(
        n16562), .A(n12289), .ZN(n12288) );
  OAI22_X1 U5196 ( .A1(n16559), .A2(n15075), .B1(n16556), .B2(n14429), .ZN(
        n12289) );
  AOI221_X1 U5197 ( .B1(\registers[12][2] ), .B2(n16661), .C1(
        \registers[15][2] ), .C2(n16658), .A(n12120), .ZN(n12119) );
  OAI22_X1 U5198 ( .A1(n16655), .A2(n15076), .B1(n16652), .B2(n14430), .ZN(
        n12120) );
  AOI221_X1 U5199 ( .B1(net226883), .B2(n16565), .C1(\registers[44][2] ), .C2(
        n16562), .A(n12136), .ZN(n12135) );
  OAI22_X1 U5200 ( .A1(n16559), .A2(n15077), .B1(n16556), .B2(n14431), .ZN(
        n12136) );
  AOI221_X1 U5201 ( .B1(\registers[12][3] ), .B2(n16661), .C1(
        \registers[15][3] ), .C2(n16658), .A(n11967), .ZN(n11966) );
  OAI22_X1 U5202 ( .A1(n16655), .A2(n14994), .B1(n16652), .B2(n14291), .ZN(
        n11967) );
  AOI221_X1 U5203 ( .B1(net226903), .B2(n16565), .C1(\registers[44][3] ), .C2(
        n16562), .A(n11983), .ZN(n11982) );
  OAI22_X1 U5204 ( .A1(n16559), .A2(n14995), .B1(n16556), .B2(n14292), .ZN(
        n11983) );
  AOI221_X1 U5205 ( .B1(\registers[12][4] ), .B2(n16661), .C1(
        \registers[15][4] ), .C2(n16658), .A(n11814), .ZN(n11813) );
  OAI22_X1 U5206 ( .A1(n16655), .A2(n15078), .B1(n16652), .B2(n14432), .ZN(
        n11814) );
  AOI221_X1 U5207 ( .B1(net226976), .B2(n16565), .C1(\registers[44][4] ), .C2(
        n16562), .A(n11830), .ZN(n11829) );
  OAI22_X1 U5208 ( .A1(n16559), .A2(n15079), .B1(n16556), .B2(n14433), .ZN(
        n11830) );
  AOI221_X1 U5209 ( .B1(\registers[12][5] ), .B2(n16661), .C1(
        \registers[15][5] ), .C2(n16658), .A(n11771), .ZN(n11770) );
  OAI22_X1 U5210 ( .A1(n16655), .A2(n15080), .B1(n16652), .B2(n14434), .ZN(
        n11771) );
  AOI221_X1 U5211 ( .B1(net226996), .B2(n16565), .C1(\registers[44][5] ), .C2(
        n16562), .A(n11787), .ZN(n11786) );
  OAI22_X1 U5212 ( .A1(n16559), .A2(n14996), .B1(n16556), .B2(n14293), .ZN(
        n11787) );
  AOI221_X1 U5213 ( .B1(\registers[12][6] ), .B2(n16661), .C1(
        \registers[15][6] ), .C2(n16658), .A(n11728), .ZN(n11727) );
  OAI22_X1 U5214 ( .A1(n16655), .A2(n15081), .B1(n16652), .B2(n14435), .ZN(
        n11728) );
  AOI221_X1 U5215 ( .B1(net227020), .B2(n16565), .C1(\registers[44][6] ), .C2(
        n16562), .A(n11744), .ZN(n11743) );
  OAI22_X1 U5216 ( .A1(n16559), .A2(n15082), .B1(n16556), .B2(n14436), .ZN(
        n11744) );
  AOI221_X1 U5217 ( .B1(\registers[12][7] ), .B2(n16661), .C1(
        \registers[15][7] ), .C2(n16658), .A(n11685), .ZN(n11684) );
  OAI22_X1 U5218 ( .A1(n16655), .A2(n15083), .B1(n16652), .B2(n14437), .ZN(
        n11685) );
  AOI221_X1 U5219 ( .B1(net227038), .B2(n16565), .C1(\registers[44][7] ), .C2(
        n16562), .A(n11701), .ZN(n11700) );
  OAI22_X1 U5220 ( .A1(n16559), .A2(n15084), .B1(n16556), .B2(n14438), .ZN(
        n11701) );
  AOI221_X1 U5221 ( .B1(\registers[12][8] ), .B2(n16661), .C1(
        \registers[15][8] ), .C2(n16658), .A(n11642), .ZN(n11641) );
  OAI22_X1 U5222 ( .A1(n16655), .A2(n15085), .B1(n16652), .B2(n14439), .ZN(
        n11642) );
  AOI221_X1 U5223 ( .B1(net227056), .B2(n16565), .C1(\registers[44][8] ), .C2(
        n16562), .A(n11658), .ZN(n11657) );
  OAI22_X1 U5224 ( .A1(n16559), .A2(n15086), .B1(n16556), .B2(n14440), .ZN(
        n11658) );
  AOI221_X1 U5225 ( .B1(\registers[12][9] ), .B2(n16661), .C1(
        \registers[15][9] ), .C2(n16658), .A(n11599), .ZN(n11598) );
  OAI22_X1 U5226 ( .A1(n16655), .A2(n15087), .B1(n16652), .B2(n14441), .ZN(
        n11599) );
  AOI221_X1 U5227 ( .B1(net227074), .B2(n16565), .C1(\registers[44][9] ), .C2(
        n16562), .A(n11615), .ZN(n11614) );
  OAI22_X1 U5228 ( .A1(n16559), .A2(n15088), .B1(n16556), .B2(n14442), .ZN(
        n11615) );
  AOI221_X1 U5229 ( .B1(\registers[12][10] ), .B2(n16661), .C1(
        \registers[15][10] ), .C2(n16658), .A(n11556), .ZN(n11555) );
  OAI22_X1 U5230 ( .A1(n16655), .A2(n15089), .B1(n16652), .B2(n14443), .ZN(
        n11556) );
  AOI221_X1 U5231 ( .B1(net227092), .B2(n16565), .C1(\registers[44][10] ), 
        .C2(n16562), .A(n11572), .ZN(n11571) );
  OAI22_X1 U5232 ( .A1(n16559), .A2(n15090), .B1(n16556), .B2(n14444), .ZN(
        n11572) );
  AOI221_X1 U5233 ( .B1(\registers[12][11] ), .B2(n16661), .C1(
        \registers[15][11] ), .C2(n16658), .A(n11513), .ZN(n11512) );
  OAI22_X1 U5234 ( .A1(n16655), .A2(n15091), .B1(n16652), .B2(n14445), .ZN(
        n11513) );
  AOI221_X1 U5235 ( .B1(net227110), .B2(n16565), .C1(\registers[44][11] ), 
        .C2(n16562), .A(n11529), .ZN(n11528) );
  OAI22_X1 U5236 ( .A1(n16559), .A2(n15092), .B1(n16556), .B2(n14446), .ZN(
        n11529) );
  AOI221_X1 U5237 ( .B1(\registers[12][12] ), .B2(n16662), .C1(
        \registers[15][12] ), .C2(n16659), .A(n11470), .ZN(n11469) );
  OAI22_X1 U5238 ( .A1(n16656), .A2(n15093), .B1(n16653), .B2(n14447), .ZN(
        n11470) );
  AOI221_X1 U5239 ( .B1(net227128), .B2(n16566), .C1(\registers[44][12] ), 
        .C2(n16563), .A(n11486), .ZN(n11485) );
  OAI22_X1 U5240 ( .A1(n16560), .A2(n15094), .B1(n16557), .B2(n14448), .ZN(
        n11486) );
  AOI221_X1 U5241 ( .B1(\registers[12][13] ), .B2(n16662), .C1(
        \registers[15][13] ), .C2(n16659), .A(n11426), .ZN(n11425) );
  OAI22_X1 U5242 ( .A1(n16656), .A2(n15095), .B1(n16653), .B2(n14449), .ZN(
        n11426) );
  AOI221_X1 U5243 ( .B1(net227146), .B2(n16566), .C1(\registers[44][13] ), 
        .C2(n16563), .A(n11442), .ZN(n11441) );
  OAI22_X1 U5244 ( .A1(n16560), .A2(n15096), .B1(n16557), .B2(n14450), .ZN(
        n11442) );
  AOI221_X1 U5245 ( .B1(\registers[12][14] ), .B2(n16662), .C1(
        \registers[15][14] ), .C2(n16659), .A(n11383), .ZN(n11382) );
  OAI22_X1 U5246 ( .A1(n16656), .A2(n15097), .B1(n16653), .B2(n14451), .ZN(
        n11383) );
  AOI221_X1 U5247 ( .B1(net227164), .B2(n16566), .C1(\registers[44][14] ), 
        .C2(n16563), .A(n11399), .ZN(n11398) );
  OAI22_X1 U5248 ( .A1(n16560), .A2(n15098), .B1(n16557), .B2(n14452), .ZN(
        n11399) );
  AOI221_X1 U5249 ( .B1(\registers[12][15] ), .B2(n16662), .C1(
        \registers[15][15] ), .C2(n16659), .A(n11340), .ZN(n11339) );
  OAI22_X1 U5250 ( .A1(n16656), .A2(n15099), .B1(n16653), .B2(n14453), .ZN(
        n11340) );
  AOI221_X1 U5251 ( .B1(net227182), .B2(n16566), .C1(\registers[44][15] ), 
        .C2(n16563), .A(n11356), .ZN(n11355) );
  OAI22_X1 U5252 ( .A1(n16560), .A2(n15100), .B1(n16557), .B2(n14454), .ZN(
        n11356) );
  AOI221_X1 U5253 ( .B1(\registers[12][16] ), .B2(n16662), .C1(
        \registers[15][16] ), .C2(n16659), .A(n11297), .ZN(n11296) );
  OAI22_X1 U5254 ( .A1(n16656), .A2(n15101), .B1(n16653), .B2(n14455), .ZN(
        n11297) );
  AOI221_X1 U5255 ( .B1(net227200), .B2(n16566), .C1(\registers[44][16] ), 
        .C2(n16563), .A(n11313), .ZN(n11312) );
  OAI22_X1 U5256 ( .A1(n16560), .A2(n15102), .B1(n16557), .B2(n14456), .ZN(
        n11313) );
  AOI221_X1 U5257 ( .B1(\registers[12][17] ), .B2(n16662), .C1(
        \registers[15][17] ), .C2(n16659), .A(n11254), .ZN(n11253) );
  OAI22_X1 U5258 ( .A1(n16656), .A2(n15103), .B1(n16653), .B2(n14457), .ZN(
        n11254) );
  AOI221_X1 U5259 ( .B1(net227218), .B2(n16566), .C1(\registers[44][17] ), 
        .C2(n16563), .A(n11270), .ZN(n11269) );
  OAI22_X1 U5260 ( .A1(n16560), .A2(n15104), .B1(n16557), .B2(n14458), .ZN(
        n11270) );
  AOI221_X1 U5261 ( .B1(\registers[12][18] ), .B2(n16662), .C1(
        \registers[15][18] ), .C2(n16659), .A(n11211), .ZN(n11210) );
  OAI22_X1 U5262 ( .A1(n16656), .A2(n15105), .B1(n16653), .B2(n14459), .ZN(
        n11211) );
  AOI221_X1 U5263 ( .B1(net227236), .B2(n16566), .C1(\registers[44][18] ), 
        .C2(n16563), .A(n11227), .ZN(n11226) );
  OAI22_X1 U5264 ( .A1(n16560), .A2(n15106), .B1(n16557), .B2(n14460), .ZN(
        n11227) );
  AOI221_X1 U5265 ( .B1(\registers[12][19] ), .B2(n16662), .C1(
        \registers[15][19] ), .C2(n16659), .A(n11168), .ZN(n11167) );
  OAI22_X1 U5266 ( .A1(n16656), .A2(n15107), .B1(n16653), .B2(n14461), .ZN(
        n11168) );
  AOI221_X1 U5267 ( .B1(net227254), .B2(n16566), .C1(\registers[44][19] ), 
        .C2(n16563), .A(n11184), .ZN(n11183) );
  OAI22_X1 U5268 ( .A1(n16560), .A2(n15108), .B1(n16557), .B2(n14462), .ZN(
        n11184) );
  AOI221_X1 U5269 ( .B1(\registers[12][20] ), .B2(n16662), .C1(
        \registers[15][20] ), .C2(n16659), .A(n11125), .ZN(n11124) );
  OAI22_X1 U5270 ( .A1(n16656), .A2(n15109), .B1(n16653), .B2(n14463), .ZN(
        n11125) );
  AOI221_X1 U5271 ( .B1(net227272), .B2(n16566), .C1(\registers[44][20] ), 
        .C2(n16563), .A(n11141), .ZN(n11140) );
  OAI22_X1 U5272 ( .A1(n16560), .A2(n15110), .B1(n16557), .B2(n14464), .ZN(
        n11141) );
  AOI221_X1 U5273 ( .B1(\registers[12][21] ), .B2(n16662), .C1(
        \registers[15][21] ), .C2(n16659), .A(n11082), .ZN(n11081) );
  OAI22_X1 U5274 ( .A1(n16656), .A2(n15111), .B1(n16653), .B2(n14465), .ZN(
        n11082) );
  AOI221_X1 U5275 ( .B1(net227290), .B2(n16566), .C1(\registers[44][21] ), 
        .C2(n16563), .A(n11098), .ZN(n11097) );
  OAI22_X1 U5276 ( .A1(n16560), .A2(n15112), .B1(n16557), .B2(n14466), .ZN(
        n11098) );
  AOI221_X1 U5277 ( .B1(\registers[12][22] ), .B2(n16662), .C1(
        \registers[15][22] ), .C2(n16659), .A(n11039), .ZN(n11038) );
  OAI22_X1 U5278 ( .A1(n16656), .A2(n15113), .B1(n16653), .B2(n14467), .ZN(
        n11039) );
  AOI221_X1 U5279 ( .B1(net227308), .B2(n16566), .C1(\registers[44][22] ), 
        .C2(n16563), .A(n11055), .ZN(n11054) );
  OAI22_X1 U5280 ( .A1(n16560), .A2(n15114), .B1(n16557), .B2(n14468), .ZN(
        n11055) );
  AOI221_X1 U5281 ( .B1(\registers[12][23] ), .B2(n16662), .C1(
        \registers[15][23] ), .C2(n16659), .A(n10996), .ZN(n10995) );
  OAI22_X1 U5282 ( .A1(n16656), .A2(n15115), .B1(n16653), .B2(n14469), .ZN(
        n10996) );
  AOI221_X1 U5283 ( .B1(net227326), .B2(n16566), .C1(\registers[44][23] ), 
        .C2(n16563), .A(n11012), .ZN(n11011) );
  OAI22_X1 U5284 ( .A1(n16560), .A2(n15116), .B1(n16557), .B2(n14470), .ZN(
        n11012) );
  AOI221_X1 U5285 ( .B1(\registers[56][0] ), .B2(n17673), .C1(
        \registers[55][0] ), .C2(n17670), .A(n12403), .ZN(n12402) );
  OAI22_X1 U5286 ( .A1(n17667), .A2(n15432), .B1(n17664), .B2(n14711), .ZN(
        n12403) );
  AOI221_X1 U5287 ( .B1(\registers[37][0] ), .B2(n17817), .C1(
        \registers[0][0] ), .C2(n17814), .A(n12379), .ZN(n12378) );
  OAI22_X1 U5288 ( .A1(n17811), .A2(n15669), .B1(n17808), .B2(n14712), .ZN(
        n12379) );
  AOI221_X1 U5289 ( .B1(\registers[56][1] ), .B2(n17673), .C1(
        \registers[55][1] ), .C2(n17670), .A(n12249), .ZN(n12248) );
  OAI22_X1 U5290 ( .A1(n17667), .A2(n15433), .B1(n17664), .B2(n14713), .ZN(
        n12249) );
  AOI221_X1 U5291 ( .B1(\registers[37][1] ), .B2(n17817), .C1(
        \registers[0][1] ), .C2(n17814), .A(n12225), .ZN(n12224) );
  OAI22_X1 U5292 ( .A1(n17811), .A2(n15670), .B1(n17808), .B2(n14714), .ZN(
        n12225) );
  AOI221_X1 U5293 ( .B1(\registers[56][2] ), .B2(n17673), .C1(
        \registers[55][2] ), .C2(n17670), .A(n12094), .ZN(n12093) );
  OAI22_X1 U5294 ( .A1(n17667), .A2(n15434), .B1(n17664), .B2(n14715), .ZN(
        n12094) );
  AOI221_X1 U5295 ( .B1(\registers[37][2] ), .B2(n17817), .C1(
        \registers[0][2] ), .C2(n17814), .A(n12070), .ZN(n12069) );
  OAI22_X1 U5296 ( .A1(n17811), .A2(n15671), .B1(n17808), .B2(n14716), .ZN(
        n12070) );
  AOI221_X1 U5297 ( .B1(\registers[56][3] ), .B2(n17673), .C1(
        \registers[55][3] ), .C2(n17670), .A(n11941), .ZN(n11940) );
  OAI22_X1 U5298 ( .A1(n17667), .A2(n15353), .B1(n17664), .B2(n14717), .ZN(
        n11941) );
  AOI221_X1 U5299 ( .B1(\registers[37][3] ), .B2(n17817), .C1(
        \registers[0][3] ), .C2(n17814), .A(n11917), .ZN(n11916) );
  OAI22_X1 U5300 ( .A1(n17811), .A2(n15365), .B1(n17808), .B2(n14640), .ZN(
        n11917) );
  AOI221_X1 U5301 ( .B1(\registers[56][4] ), .B2(n17673), .C1(
        \registers[55][4] ), .C2(n17670), .A(n10498), .ZN(n10497) );
  OAI22_X1 U5302 ( .A1(n17667), .A2(n15354), .B1(n17664), .B2(n14718), .ZN(
        n10498) );
  AOI221_X1 U5303 ( .B1(\registers[37][4] ), .B2(n17817), .C1(
        \registers[0][4] ), .C2(n17814), .A(n10474), .ZN(n10473) );
  OAI22_X1 U5304 ( .A1(n17811), .A2(n15672), .B1(n17808), .B2(n14719), .ZN(
        n10474) );
  AOI221_X1 U5305 ( .B1(\registers[56][5] ), .B2(n17673), .C1(
        \registers[55][5] ), .C2(n17670), .A(n10388), .ZN(n10387) );
  OAI22_X1 U5306 ( .A1(n17667), .A2(n15355), .B1(n17664), .B2(n14720), .ZN(
        n10388) );
  AOI221_X1 U5307 ( .B1(\registers[37][5] ), .B2(n17817), .C1(
        \registers[0][5] ), .C2(n17814), .A(n10364), .ZN(n10363) );
  OAI22_X1 U5308 ( .A1(n17811), .A2(n15673), .B1(n17808), .B2(n14721), .ZN(
        n10364) );
  AOI221_X1 U5309 ( .B1(\registers[56][6] ), .B2(n17673), .C1(
        \registers[55][6] ), .C2(n17670), .A(n10276), .ZN(n10275) );
  OAI22_X1 U5310 ( .A1(n17667), .A2(n15435), .B1(n17664), .B2(n14722), .ZN(
        n10276) );
  AOI221_X1 U5311 ( .B1(\registers[37][6] ), .B2(n17817), .C1(
        \registers[0][6] ), .C2(n17814), .A(n10252), .ZN(n10251) );
  OAI22_X1 U5312 ( .A1(n17811), .A2(n15674), .B1(n17808), .B2(n14723), .ZN(
        n10252) );
  AOI221_X1 U5313 ( .B1(\registers[56][7] ), .B2(n17673), .C1(
        \registers[55][7] ), .C2(n17670), .A(n7640), .ZN(n7639) );
  OAI22_X1 U5314 ( .A1(n17667), .A2(n15436), .B1(n17664), .B2(n14724), .ZN(
        n7640) );
  AOI221_X1 U5315 ( .B1(\registers[37][7] ), .B2(n17817), .C1(
        \registers[0][7] ), .C2(n17814), .A(n7616), .ZN(n7615) );
  OAI22_X1 U5316 ( .A1(n17811), .A2(n15675), .B1(n17808), .B2(n14725), .ZN(
        n7616) );
  AOI221_X1 U5317 ( .B1(\registers[56][8] ), .B2(n17673), .C1(
        \registers[55][8] ), .C2(n17670), .A(n7525), .ZN(n7524) );
  OAI22_X1 U5318 ( .A1(n17667), .A2(n15437), .B1(n17664), .B2(n14726), .ZN(
        n7525) );
  AOI221_X1 U5319 ( .B1(\registers[37][8] ), .B2(n17817), .C1(
        \registers[0][8] ), .C2(n17814), .A(n7501), .ZN(n7500) );
  OAI22_X1 U5320 ( .A1(n17811), .A2(n15676), .B1(n17808), .B2(n14727), .ZN(
        n7501) );
  AOI221_X1 U5321 ( .B1(\registers[56][9] ), .B2(n17673), .C1(
        \registers[55][9] ), .C2(n17670), .A(n7416), .ZN(n7415) );
  OAI22_X1 U5322 ( .A1(n17667), .A2(n15438), .B1(n17664), .B2(n14728), .ZN(
        n7416) );
  AOI221_X1 U5323 ( .B1(\registers[37][9] ), .B2(n17817), .C1(
        \registers[0][9] ), .C2(n17814), .A(n7392), .ZN(n7391) );
  OAI22_X1 U5324 ( .A1(n17811), .A2(n15677), .B1(n17808), .B2(n14729), .ZN(
        n7392) );
  AOI221_X1 U5325 ( .B1(\registers[56][10] ), .B2(n17673), .C1(
        \registers[55][10] ), .C2(n17670), .A(n7307), .ZN(n7306) );
  OAI22_X1 U5326 ( .A1(n17667), .A2(n15439), .B1(n17664), .B2(n14730), .ZN(
        n7307) );
  AOI221_X1 U5327 ( .B1(\registers[37][10] ), .B2(n17817), .C1(
        \registers[0][10] ), .C2(n17814), .A(n7283), .ZN(n7282) );
  OAI22_X1 U5328 ( .A1(n17811), .A2(n15678), .B1(n17808), .B2(n14731), .ZN(
        n7283) );
  AOI221_X1 U5329 ( .B1(\registers[56][11] ), .B2(n17674), .C1(
        \registers[55][11] ), .C2(n17671), .A(n7193), .ZN(n7192) );
  OAI22_X1 U5330 ( .A1(n17668), .A2(n15440), .B1(n17665), .B2(n14732), .ZN(
        n7193) );
  AOI221_X1 U5331 ( .B1(\registers[37][11] ), .B2(n17818), .C1(
        \registers[0][11] ), .C2(n17815), .A(n7169), .ZN(n7168) );
  OAI22_X1 U5332 ( .A1(n17812), .A2(n15679), .B1(n17809), .B2(n14733), .ZN(
        n7169) );
  AOI221_X1 U5333 ( .B1(\registers[56][12] ), .B2(n17674), .C1(
        \registers[55][12] ), .C2(n17671), .A(n7084), .ZN(n7083) );
  OAI22_X1 U5334 ( .A1(n17668), .A2(n15441), .B1(n17665), .B2(n14734), .ZN(
        n7084) );
  AOI221_X1 U5335 ( .B1(\registers[37][12] ), .B2(n17818), .C1(
        \registers[0][12] ), .C2(n17815), .A(n7060), .ZN(n7059) );
  OAI22_X1 U5336 ( .A1(n17812), .A2(n15680), .B1(n17809), .B2(n14735), .ZN(
        n7060) );
  AOI221_X1 U5337 ( .B1(\registers[56][13] ), .B2(n17674), .C1(
        \registers[55][13] ), .C2(n17671), .A(n6975), .ZN(n6974) );
  OAI22_X1 U5338 ( .A1(n17668), .A2(n15442), .B1(n17665), .B2(n14736), .ZN(
        n6975) );
  AOI221_X1 U5339 ( .B1(\registers[37][13] ), .B2(n17818), .C1(
        \registers[0][13] ), .C2(n17815), .A(n6951), .ZN(n6950) );
  OAI22_X1 U5340 ( .A1(n17812), .A2(n15681), .B1(n17809), .B2(n14737), .ZN(
        n6951) );
  AOI221_X1 U5341 ( .B1(\registers[56][14] ), .B2(n17674), .C1(
        \registers[55][14] ), .C2(n17671), .A(n6866), .ZN(n6865) );
  OAI22_X1 U5342 ( .A1(n17668), .A2(n15443), .B1(n17665), .B2(n14738), .ZN(
        n6866) );
  AOI221_X1 U5343 ( .B1(\registers[37][14] ), .B2(n17818), .C1(
        \registers[0][14] ), .C2(n17815), .A(n6842), .ZN(n6841) );
  OAI22_X1 U5344 ( .A1(n17812), .A2(n15682), .B1(n17809), .B2(n14739), .ZN(
        n6842) );
  AOI221_X1 U5345 ( .B1(\registers[56][15] ), .B2(n17674), .C1(
        \registers[55][15] ), .C2(n17671), .A(n6757), .ZN(n6756) );
  OAI22_X1 U5346 ( .A1(n17668), .A2(n15444), .B1(n17665), .B2(n14740), .ZN(
        n6757) );
  AOI221_X1 U5347 ( .B1(\registers[37][15] ), .B2(n17818), .C1(
        \registers[0][15] ), .C2(n17815), .A(n6733), .ZN(n6732) );
  OAI22_X1 U5348 ( .A1(n17812), .A2(n15683), .B1(n17809), .B2(n14741), .ZN(
        n6733) );
  AOI221_X1 U5349 ( .B1(\registers[56][16] ), .B2(n17674), .C1(
        \registers[55][16] ), .C2(n17671), .A(n6617), .ZN(n6616) );
  OAI22_X1 U5350 ( .A1(n17668), .A2(n15445), .B1(n17665), .B2(n14742), .ZN(
        n6617) );
  AOI221_X1 U5351 ( .B1(\registers[37][16] ), .B2(n17818), .C1(
        \registers[0][16] ), .C2(n17815), .A(n6573), .ZN(n6572) );
  OAI22_X1 U5352 ( .A1(n17812), .A2(n15684), .B1(n17809), .B2(n14743), .ZN(
        n6573) );
  AOI221_X1 U5353 ( .B1(\registers[56][17] ), .B2(n17674), .C1(
        \registers[55][17] ), .C2(n17671), .A(n6430), .ZN(n6429) );
  OAI22_X1 U5354 ( .A1(n17668), .A2(n15446), .B1(n17665), .B2(n14744), .ZN(
        n6430) );
  AOI221_X1 U5355 ( .B1(\registers[37][17] ), .B2(n17818), .C1(
        \registers[0][17] ), .C2(n17815), .A(n6386), .ZN(n6385) );
  OAI22_X1 U5356 ( .A1(n17812), .A2(n15685), .B1(n17809), .B2(n14745), .ZN(
        n6386) );
  AOI221_X1 U5357 ( .B1(\registers[56][18] ), .B2(n17674), .C1(
        \registers[55][18] ), .C2(n17671), .A(n6245), .ZN(n6244) );
  OAI22_X1 U5358 ( .A1(n17668), .A2(n15447), .B1(n17665), .B2(n14746), .ZN(
        n6245) );
  AOI221_X1 U5359 ( .B1(\registers[37][18] ), .B2(n17818), .C1(
        \registers[0][18] ), .C2(n17815), .A(n6199), .ZN(n6198) );
  OAI22_X1 U5360 ( .A1(n17812), .A2(n15686), .B1(n17809), .B2(n14747), .ZN(
        n6199) );
  AOI221_X1 U5361 ( .B1(\registers[56][19] ), .B2(n17674), .C1(
        \registers[55][19] ), .C2(n17671), .A(n6059), .ZN(n6058) );
  OAI22_X1 U5362 ( .A1(n17668), .A2(n15448), .B1(n17665), .B2(n14748), .ZN(
        n6059) );
  AOI221_X1 U5363 ( .B1(\registers[37][19] ), .B2(n17818), .C1(
        \registers[0][19] ), .C2(n17815), .A(n6014), .ZN(n6013) );
  OAI22_X1 U5364 ( .A1(n17812), .A2(n15687), .B1(n17809), .B2(n14749), .ZN(
        n6014) );
  AOI221_X1 U5365 ( .B1(\registers[56][20] ), .B2(n17674), .C1(
        \registers[55][20] ), .C2(n17671), .A(n5872), .ZN(n5871) );
  OAI22_X1 U5366 ( .A1(n17668), .A2(n15449), .B1(n17665), .B2(n14750), .ZN(
        n5872) );
  AOI221_X1 U5367 ( .B1(\registers[37][20] ), .B2(n17818), .C1(
        \registers[0][20] ), .C2(n17815), .A(n5842), .ZN(n5826) );
  OAI22_X1 U5368 ( .A1(n17812), .A2(n15688), .B1(n17809), .B2(n14751), .ZN(
        n5842) );
  AOI221_X1 U5369 ( .B1(\registers[56][21] ), .B2(n17674), .C1(
        \registers[55][21] ), .C2(n17671), .A(n5686), .ZN(n5684) );
  OAI22_X1 U5370 ( .A1(n17668), .A2(n15450), .B1(n17665), .B2(n14752), .ZN(
        n5686) );
  AOI221_X1 U5371 ( .B1(\registers[37][21] ), .B2(n17818), .C1(
        \registers[0][21] ), .C2(n17815), .A(n5655), .ZN(n5654) );
  OAI22_X1 U5372 ( .A1(n17812), .A2(n15689), .B1(n17809), .B2(n14753), .ZN(
        n5655) );
  AOI221_X1 U5373 ( .B1(\registers[56][22] ), .B2(n17674), .C1(
        \registers[55][22] ), .C2(n17671), .A(n5501), .ZN(n5499) );
  OAI22_X1 U5374 ( .A1(n17668), .A2(n15451), .B1(n17665), .B2(n14754), .ZN(
        n5501) );
  AOI221_X1 U5375 ( .B1(\registers[37][22] ), .B2(n17818), .C1(
        \registers[0][22] ), .C2(n17815), .A(n5468), .ZN(n5467) );
  OAI22_X1 U5376 ( .A1(n17812), .A2(n15690), .B1(n17809), .B2(n14755), .ZN(
        n5468) );
  AOI221_X1 U5377 ( .B1(\registers[56][31] ), .B2(n17673), .C1(
        \registers[55][31] ), .C2(n17670), .A(n14191), .ZN(n14190) );
  OAI22_X1 U5378 ( .A1(n17667), .A2(n14670), .B1(n17664), .B2(n15318), .ZN(
        n14191) );
  AOI221_X1 U5379 ( .B1(\registers[37][31] ), .B2(n17817), .C1(
        \registers[0][31] ), .C2(n17814), .A(n14084), .ZN(n14083) );
  OAI22_X1 U5380 ( .A1(n17811), .A2(n15691), .B1(n17808), .B2(n14756), .ZN(
        n14084) );
  AOI221_X1 U5381 ( .B1(\registers[45][24] ), .B2(n16303), .C1(
        \registers[4][24] ), .C2(n16300), .A(n12920), .ZN(n12917) );
  OAI22_X1 U5382 ( .A1(n16297), .A2(n11907), .B1(n16294), .B2(n14875), .ZN(
        n12920) );
  AOI221_X1 U5383 ( .B1(\registers[5][24] ), .B2(n16252), .C1(
        \registers[59][24] ), .C2(n16249), .A(n12928), .ZN(n12925) );
  OAI22_X1 U5384 ( .A1(n16246), .A2(n12342), .B1(n16243), .B2(n14876), .ZN(
        n12928) );
  AOI221_X1 U5385 ( .B1(\registers[45][25] ), .B2(n16303), .C1(
        \registers[4][25] ), .C2(n16300), .A(n12878), .ZN(n12875) );
  OAI22_X1 U5386 ( .A1(n16297), .A2(n11945), .B1(n16294), .B2(n14877), .ZN(
        n12878) );
  AOI221_X1 U5387 ( .B1(\registers[5][25] ), .B2(n16252), .C1(
        \registers[59][25] ), .C2(n16249), .A(n12886), .ZN(n12883) );
  OAI22_X1 U5388 ( .A1(n16246), .A2(n12343), .B1(n16243), .B2(n14878), .ZN(
        n12886) );
  AOI221_X1 U5389 ( .B1(\registers[45][26] ), .B2(n16303), .C1(
        \registers[4][26] ), .C2(n16300), .A(n12836), .ZN(n12833) );
  OAI22_X1 U5390 ( .A1(n16297), .A2(n11946), .B1(n16294), .B2(n14879), .ZN(
        n12836) );
  AOI221_X1 U5391 ( .B1(\registers[5][26] ), .B2(n16252), .C1(
        \registers[59][26] ), .C2(n16249), .A(n12844), .ZN(n12841) );
  OAI22_X1 U5392 ( .A1(n16246), .A2(n12344), .B1(n16243), .B2(n14880), .ZN(
        n12844) );
  AOI221_X1 U5393 ( .B1(\registers[45][27] ), .B2(n16303), .C1(
        \registers[4][27] ), .C2(n16300), .A(n12794), .ZN(n12791) );
  OAI22_X1 U5394 ( .A1(n16297), .A2(n11947), .B1(n16294), .B2(n14881), .ZN(
        n12794) );
  AOI221_X1 U5395 ( .B1(\registers[5][27] ), .B2(n16252), .C1(
        \registers[59][27] ), .C2(n16249), .A(n12802), .ZN(n12799) );
  OAI22_X1 U5396 ( .A1(n16246), .A2(n12345), .B1(n16243), .B2(n14882), .ZN(
        n12802) );
  AOI221_X1 U5397 ( .B1(\registers[45][28] ), .B2(n16303), .C1(
        \registers[4][28] ), .C2(n16300), .A(n12752), .ZN(n12749) );
  OAI22_X1 U5398 ( .A1(n16297), .A2(n11948), .B1(n16294), .B2(n14883), .ZN(
        n12752) );
  AOI221_X1 U5399 ( .B1(\registers[5][28] ), .B2(n16252), .C1(
        \registers[59][28] ), .C2(n16249), .A(n12760), .ZN(n12757) );
  OAI22_X1 U5400 ( .A1(n16246), .A2(n12346), .B1(n16243), .B2(n14884), .ZN(
        n12760) );
  AOI221_X1 U5401 ( .B1(\registers[45][29] ), .B2(n16303), .C1(
        \registers[4][29] ), .C2(n16300), .A(n12710), .ZN(n12707) );
  OAI22_X1 U5402 ( .A1(n16297), .A2(n11949), .B1(n16294), .B2(n14885), .ZN(
        n12710) );
  AOI221_X1 U5403 ( .B1(\registers[5][29] ), .B2(n16252), .C1(
        \registers[59][29] ), .C2(n16249), .A(n12718), .ZN(n12715) );
  OAI22_X1 U5404 ( .A1(n16246), .A2(n12347), .B1(n16243), .B2(n14886), .ZN(
        n12718) );
  AOI221_X1 U5405 ( .B1(\registers[45][30] ), .B2(n16303), .C1(
        \registers[4][30] ), .C2(n16300), .A(n12667), .ZN(n12664) );
  OAI22_X1 U5406 ( .A1(n16297), .A2(n11670), .B1(n16294), .B2(n14854), .ZN(
        n12667) );
  AOI221_X1 U5407 ( .B1(\registers[5][30] ), .B2(n16252), .C1(
        \registers[59][30] ), .C2(n16249), .A(n12676), .ZN(n12673) );
  OAI22_X1 U5408 ( .A1(n16246), .A2(n12196), .B1(n16243), .B2(n14858), .ZN(
        n12676) );
  AOI221_X1 U5409 ( .B1(\registers[45][31] ), .B2(n16303), .C1(
        \registers[4][31] ), .C2(n16300), .A(n12593), .ZN(n12584) );
  OAI22_X1 U5410 ( .A1(n16297), .A2(n11950), .B1(n16294), .B2(n14887), .ZN(
        n12593) );
  AOI221_X1 U5411 ( .B1(\registers[5][31] ), .B2(n16252), .C1(
        \registers[59][31] ), .C2(n16249), .A(n12620), .ZN(n12610) );
  OAI22_X1 U5412 ( .A1(n16246), .A2(n12348), .B1(n16243), .B2(n14859), .ZN(
        n12620) );
  AOI221_X1 U5413 ( .B1(\registers[45][24] ), .B2(n16555), .C1(
        \registers[48][24] ), .C2(n16552), .A(n10970), .ZN(n10967) );
  OAI22_X1 U5414 ( .A1(n16549), .A2(n11907), .B1(n16546), .B2(n14875), .ZN(
        n10970) );
  AOI221_X1 U5415 ( .B1(\registers[5][24] ), .B2(n16504), .C1(
        \registers[59][24] ), .C2(n16501), .A(n10978), .ZN(n10975) );
  OAI22_X1 U5416 ( .A1(n16498), .A2(n12342), .B1(n16495), .B2(n14876), .ZN(
        n10978) );
  AOI221_X1 U5417 ( .B1(\registers[45][25] ), .B2(n16555), .C1(
        \registers[48][25] ), .C2(n16552), .A(n10927), .ZN(n10924) );
  OAI22_X1 U5418 ( .A1(n16549), .A2(n11945), .B1(n16546), .B2(n14877), .ZN(
        n10927) );
  AOI221_X1 U5419 ( .B1(\registers[5][25] ), .B2(n16504), .C1(
        \registers[59][25] ), .C2(n16501), .A(n10935), .ZN(n10932) );
  OAI22_X1 U5420 ( .A1(n16498), .A2(n12343), .B1(n16495), .B2(n14878), .ZN(
        n10935) );
  AOI221_X1 U5421 ( .B1(\registers[45][26] ), .B2(n16555), .C1(
        \registers[48][26] ), .C2(n16552), .A(n10884), .ZN(n10881) );
  OAI22_X1 U5422 ( .A1(n16549), .A2(n11946), .B1(n16546), .B2(n14879), .ZN(
        n10884) );
  AOI221_X1 U5423 ( .B1(\registers[5][26] ), .B2(n16504), .C1(
        \registers[59][26] ), .C2(n16501), .A(n10892), .ZN(n10889) );
  OAI22_X1 U5424 ( .A1(n16498), .A2(n12344), .B1(n16495), .B2(n14880), .ZN(
        n10892) );
  AOI221_X1 U5425 ( .B1(\registers[45][27] ), .B2(n16555), .C1(
        \registers[48][27] ), .C2(n16552), .A(n10841), .ZN(n10838) );
  OAI22_X1 U5426 ( .A1(n16549), .A2(n11947), .B1(n16546), .B2(n14881), .ZN(
        n10841) );
  AOI221_X1 U5427 ( .B1(\registers[5][27] ), .B2(n16504), .C1(
        \registers[59][27] ), .C2(n16501), .A(n10849), .ZN(n10846) );
  OAI22_X1 U5428 ( .A1(n16498), .A2(n12345), .B1(n16495), .B2(n14882), .ZN(
        n10849) );
  AOI221_X1 U5429 ( .B1(\registers[45][28] ), .B2(n16555), .C1(
        \registers[48][28] ), .C2(n16552), .A(n10798), .ZN(n10795) );
  OAI22_X1 U5430 ( .A1(n16549), .A2(n11948), .B1(n16546), .B2(n14883), .ZN(
        n10798) );
  AOI221_X1 U5431 ( .B1(\registers[5][28] ), .B2(n16504), .C1(
        \registers[59][28] ), .C2(n16501), .A(n10806), .ZN(n10803) );
  OAI22_X1 U5432 ( .A1(n16498), .A2(n12346), .B1(n16495), .B2(n14884), .ZN(
        n10806) );
  AOI221_X1 U5433 ( .B1(\registers[45][29] ), .B2(n16555), .C1(
        \registers[48][29] ), .C2(n16552), .A(n10755), .ZN(n10752) );
  OAI22_X1 U5434 ( .A1(n16549), .A2(n11949), .B1(n16546), .B2(n14885), .ZN(
        n10755) );
  AOI221_X1 U5435 ( .B1(\registers[5][29] ), .B2(n16504), .C1(
        \registers[59][29] ), .C2(n16501), .A(n10763), .ZN(n10760) );
  OAI22_X1 U5436 ( .A1(n16498), .A2(n12347), .B1(n16495), .B2(n14886), .ZN(
        n10763) );
  AOI221_X1 U5437 ( .B1(\registers[45][30] ), .B2(n16555), .C1(
        \registers[48][30] ), .C2(n16552), .A(n10707), .ZN(n10702) );
  OAI22_X1 U5438 ( .A1(n16549), .A2(n11670), .B1(n16546), .B2(n14854), .ZN(
        n10707) );
  AOI221_X1 U5439 ( .B1(\registers[5][30] ), .B2(n16504), .C1(
        \registers[59][30] ), .C2(n16501), .A(n10718), .ZN(n10715) );
  OAI22_X1 U5440 ( .A1(n16498), .A2(n12196), .B1(n16495), .B2(n14858), .ZN(
        n10718) );
  AOI221_X1 U5441 ( .B1(\registers[45][31] ), .B2(n16555), .C1(
        \registers[48][31] ), .C2(n16552), .A(n10609), .ZN(n10598) );
  OAI22_X1 U5442 ( .A1(n16549), .A2(n11950), .B1(n16546), .B2(n14887), .ZN(
        n10609) );
  AOI221_X1 U5443 ( .B1(\registers[5][31] ), .B2(n16504), .C1(
        \registers[59][31] ), .C2(n16501), .A(n10643), .ZN(n10630) );
  OAI22_X1 U5444 ( .A1(n16498), .A2(n12348), .B1(n16495), .B2(n14859), .ZN(
        n10643) );
  AOI221_X1 U5445 ( .B1(\registers[63][23] ), .B2(n17663), .C1(
        \registers[62][23] ), .C2(n17660), .A(n5315), .ZN(n5312) );
  OAI22_X1 U5446 ( .A1(n17657), .A2(n14050), .B1(n17654), .B2(n15319), .ZN(
        n5315) );
  AOI221_X1 U5447 ( .B1(\registers[11][23] ), .B2(n17807), .C1(net227324), 
        .C2(n17804), .A(n5282), .ZN(n5279) );
  OAI22_X1 U5448 ( .A1(n17801), .A2(n15692), .B1(n17798), .B2(n11874), .ZN(
        n5282) );
  AOI221_X1 U5449 ( .B1(\registers[63][24] ), .B2(n17663), .C1(
        \registers[62][24] ), .C2(n17660), .A(n5143), .ZN(n5140) );
  OAI22_X1 U5450 ( .A1(n17657), .A2(n12342), .B1(n17654), .B2(n15320), .ZN(
        n5143) );
  AOI221_X1 U5451 ( .B1(\registers[11][24] ), .B2(n17807), .C1(net227342), 
        .C2(n17804), .A(n5117), .ZN(n5113) );
  OAI22_X1 U5452 ( .A1(n17801), .A2(n15693), .B1(n17798), .B2(n11875), .ZN(
        n5117) );
  AOI221_X1 U5453 ( .B1(\registers[63][25] ), .B2(n17663), .C1(
        \registers[62][25] ), .C2(n17660), .A(n5029), .ZN(n5026) );
  OAI22_X1 U5454 ( .A1(n17657), .A2(n12343), .B1(n17654), .B2(n15321), .ZN(
        n5029) );
  AOI221_X1 U5455 ( .B1(\registers[11][25] ), .B2(n17807), .C1(net227360), 
        .C2(n17804), .A(n5003), .ZN(n5000) );
  OAI22_X1 U5456 ( .A1(n17801), .A2(n15694), .B1(n17798), .B2(n11876), .ZN(
        n5003) );
  AOI221_X1 U5457 ( .B1(\registers[63][26] ), .B2(n17663), .C1(
        \registers[62][26] ), .C2(n17660), .A(n4911), .ZN(n4908) );
  OAI22_X1 U5458 ( .A1(n17657), .A2(n12344), .B1(n17654), .B2(n15322), .ZN(
        n4911) );
  AOI221_X1 U5459 ( .B1(\registers[11][26] ), .B2(n17807), .C1(net227378), 
        .C2(n17804), .A(n4881), .ZN(n4878) );
  OAI22_X1 U5460 ( .A1(n17801), .A2(n15695), .B1(n17798), .B2(n11877), .ZN(
        n4881) );
  AOI221_X1 U5461 ( .B1(\registers[63][27] ), .B2(n17663), .C1(
        \registers[62][27] ), .C2(n17660), .A(n4780), .ZN(n4777) );
  OAI22_X1 U5462 ( .A1(n17657), .A2(n12345), .B1(n17654), .B2(n15323), .ZN(
        n4780) );
  AOI221_X1 U5463 ( .B1(\registers[11][27] ), .B2(n17807), .C1(net227396), 
        .C2(n17804), .A(n4752), .ZN(n4749) );
  OAI22_X1 U5464 ( .A1(n17801), .A2(n15696), .B1(n17798), .B2(n11878), .ZN(
        n4752) );
  AOI221_X1 U5465 ( .B1(\registers[63][28] ), .B2(n17663), .C1(
        \registers[62][28] ), .C2(n17660), .A(n4651), .ZN(n4648) );
  OAI22_X1 U5466 ( .A1(n17657), .A2(n12346), .B1(n17654), .B2(n15324), .ZN(
        n4651) );
  AOI221_X1 U5467 ( .B1(\registers[11][28] ), .B2(n17807), .C1(net227414), 
        .C2(n17804), .A(n4623), .ZN(n4620) );
  OAI22_X1 U5468 ( .A1(n17801), .A2(n15697), .B1(n17798), .B2(n11879), .ZN(
        n4623) );
  AOI221_X1 U5469 ( .B1(\registers[63][29] ), .B2(n17663), .C1(
        \registers[62][29] ), .C2(n17660), .A(n4522), .ZN(n4519) );
  OAI22_X1 U5470 ( .A1(n17657), .A2(n12347), .B1(n17654), .B2(n15325), .ZN(
        n4522) );
  AOI221_X1 U5471 ( .B1(\registers[11][29] ), .B2(n17807), .C1(net227432), 
        .C2(n17804), .A(n4490), .ZN(n4487) );
  OAI22_X1 U5472 ( .A1(n17801), .A2(n15698), .B1(n17798), .B2(n11880), .ZN(
        n4490) );
  AOI221_X1 U5473 ( .B1(\registers[63][30] ), .B2(n17663), .C1(
        \registers[62][30] ), .C2(n17660), .A(n4227), .ZN(n4217) );
  OAI22_X1 U5474 ( .A1(n17657), .A2(n12196), .B1(n17654), .B2(n15271), .ZN(
        n4227) );
  AOI221_X1 U5475 ( .B1(\registers[11][30] ), .B2(n17807), .C1(net227450), 
        .C2(n17804), .A(n4118), .ZN(n4103) );
  OAI22_X1 U5476 ( .A1(n17801), .A2(n15281), .B1(n17798), .B2(n11541), .ZN(
        n4118) );
  AOI221_X1 U5477 ( .B1(\registers[45][0] ), .B2(n16301), .C1(
        \registers[4][0] ), .C2(n16298), .A(n13954), .ZN(n13950) );
  OAI22_X1 U5478 ( .A1(n16295), .A2(n11951), .B1(n16292), .B2(n14888), .ZN(
        n13954) );
  AOI221_X1 U5479 ( .B1(\registers[45][1] ), .B2(n16301), .C1(
        \registers[4][1] ), .C2(n16298), .A(n13886), .ZN(n13883) );
  OAI22_X1 U5480 ( .A1(n16295), .A2(n11952), .B1(n16292), .B2(n14889), .ZN(
        n13886) );
  AOI221_X1 U5481 ( .B1(\registers[45][2] ), .B2(n16301), .C1(
        \registers[4][2] ), .C2(n16298), .A(n13844), .ZN(n13841) );
  OAI22_X1 U5482 ( .A1(n16295), .A2(n11995), .B1(n16292), .B2(n14890), .ZN(
        n13844) );
  AOI221_X1 U5483 ( .B1(\registers[45][3] ), .B2(n16301), .C1(
        \registers[4][3] ), .C2(n16298), .A(n13802), .ZN(n13799) );
  OAI22_X1 U5484 ( .A1(n16295), .A2(n11905), .B1(n16292), .B2(n14861), .ZN(
        n13802) );
  AOI221_X1 U5485 ( .B1(\registers[45][4] ), .B2(n16301), .C1(
        \registers[4][4] ), .C2(n16298), .A(n13760), .ZN(n13757) );
  OAI22_X1 U5486 ( .A1(n16295), .A2(n11997), .B1(n16292), .B2(n14891), .ZN(
        n13760) );
  AOI221_X1 U5487 ( .B1(\registers[45][5] ), .B2(n16301), .C1(
        \registers[4][5] ), .C2(n16298), .A(n13718), .ZN(n13715) );
  OAI22_X1 U5488 ( .A1(n16295), .A2(n11906), .B1(n16292), .B2(n14862), .ZN(
        n13718) );
  AOI221_X1 U5489 ( .B1(\registers[45][6] ), .B2(n16301), .C1(
        \registers[4][6] ), .C2(n16298), .A(n13676), .ZN(n13673) );
  OAI22_X1 U5490 ( .A1(n16295), .A2(n11998), .B1(n16292), .B2(n14892), .ZN(
        n13676) );
  AOI221_X1 U5491 ( .B1(\registers[45][7] ), .B2(n16301), .C1(
        \registers[4][7] ), .C2(n16298), .A(n13634), .ZN(n13631) );
  OAI22_X1 U5492 ( .A1(n16295), .A2(n11999), .B1(n16292), .B2(n14893), .ZN(
        n13634) );
  AOI221_X1 U5493 ( .B1(\registers[45][8] ), .B2(n16301), .C1(
        \registers[4][8] ), .C2(n16298), .A(n13592), .ZN(n13589) );
  OAI22_X1 U5494 ( .A1(n16295), .A2(n12000), .B1(n16292), .B2(n14894), .ZN(
        n13592) );
  AOI221_X1 U5495 ( .B1(\registers[45][9] ), .B2(n16301), .C1(
        \registers[4][9] ), .C2(n16298), .A(n13550), .ZN(n13547) );
  OAI22_X1 U5496 ( .A1(n16295), .A2(n12001), .B1(n16292), .B2(n14895), .ZN(
        n13550) );
  AOI221_X1 U5497 ( .B1(\registers[45][10] ), .B2(n16301), .C1(
        \registers[4][10] ), .C2(n16298), .A(n13508), .ZN(n13505) );
  OAI22_X1 U5498 ( .A1(n16295), .A2(n12002), .B1(n16292), .B2(n14896), .ZN(
        n13508) );
  AOI221_X1 U5499 ( .B1(\registers[45][11] ), .B2(n16301), .C1(
        \registers[4][11] ), .C2(n16298), .A(n13466), .ZN(n13463) );
  OAI22_X1 U5500 ( .A1(n16295), .A2(n12003), .B1(n16292), .B2(n14897), .ZN(
        n13466) );
  AOI221_X1 U5501 ( .B1(\registers[45][12] ), .B2(n16302), .C1(
        \registers[4][12] ), .C2(n16299), .A(n13424), .ZN(n13421) );
  OAI22_X1 U5502 ( .A1(n16296), .A2(n12004), .B1(n16293), .B2(n14898), .ZN(
        n13424) );
  AOI221_X1 U5503 ( .B1(\registers[45][13] ), .B2(n16302), .C1(
        \registers[4][13] ), .C2(n16299), .A(n13382), .ZN(n13379) );
  OAI22_X1 U5504 ( .A1(n16296), .A2(n12005), .B1(n16293), .B2(n14899), .ZN(
        n13382) );
  AOI221_X1 U5505 ( .B1(\registers[45][14] ), .B2(n16302), .C1(
        \registers[4][14] ), .C2(n16299), .A(n13340), .ZN(n13337) );
  OAI22_X1 U5506 ( .A1(n16296), .A2(n12006), .B1(n16293), .B2(n14900), .ZN(
        n13340) );
  AOI221_X1 U5507 ( .B1(\registers[45][15] ), .B2(n16302), .C1(
        \registers[4][15] ), .C2(n16299), .A(n13298), .ZN(n13295) );
  OAI22_X1 U5508 ( .A1(n16296), .A2(n12007), .B1(n16293), .B2(n14901), .ZN(
        n13298) );
  AOI221_X1 U5509 ( .B1(\registers[45][16] ), .B2(n16302), .C1(
        \registers[4][16] ), .C2(n16299), .A(n13256), .ZN(n13253) );
  OAI22_X1 U5510 ( .A1(n16296), .A2(n12008), .B1(n16293), .B2(n14902), .ZN(
        n13256) );
  AOI221_X1 U5511 ( .B1(\registers[45][17] ), .B2(n16302), .C1(
        \registers[4][17] ), .C2(n16299), .A(n13214), .ZN(n13211) );
  OAI22_X1 U5512 ( .A1(n16296), .A2(n12009), .B1(n16293), .B2(n14903), .ZN(
        n13214) );
  AOI221_X1 U5513 ( .B1(\registers[45][18] ), .B2(n16302), .C1(
        \registers[4][18] ), .C2(n16299), .A(n13172), .ZN(n13169) );
  OAI22_X1 U5514 ( .A1(n16296), .A2(n12010), .B1(n16293), .B2(n14904), .ZN(
        n13172) );
  AOI221_X1 U5515 ( .B1(\registers[45][19] ), .B2(n16302), .C1(
        \registers[4][19] ), .C2(n16299), .A(n13130), .ZN(n13127) );
  OAI22_X1 U5516 ( .A1(n16296), .A2(n12011), .B1(n16293), .B2(n14905), .ZN(
        n13130) );
  AOI221_X1 U5517 ( .B1(\registers[45][20] ), .B2(n16302), .C1(
        \registers[4][20] ), .C2(n16299), .A(n13088), .ZN(n13085) );
  OAI22_X1 U5518 ( .A1(n16296), .A2(n12012), .B1(n16293), .B2(n14906), .ZN(
        n13088) );
  AOI221_X1 U5519 ( .B1(\registers[45][21] ), .B2(n16302), .C1(
        \registers[4][21] ), .C2(n16299), .A(n13046), .ZN(n13043) );
  OAI22_X1 U5520 ( .A1(n16296), .A2(n12013), .B1(n16293), .B2(n14907), .ZN(
        n13046) );
  AOI221_X1 U5521 ( .B1(\registers[45][22] ), .B2(n16302), .C1(
        \registers[4][22] ), .C2(n16299), .A(n13004), .ZN(n13001) );
  OAI22_X1 U5522 ( .A1(n16296), .A2(n12014), .B1(n16293), .B2(n14908), .ZN(
        n13004) );
  AOI221_X1 U5523 ( .B1(\registers[45][23] ), .B2(n16302), .C1(
        \registers[4][23] ), .C2(n16299), .A(n12962), .ZN(n12959) );
  OAI22_X1 U5524 ( .A1(n16296), .A2(n12015), .B1(n16293), .B2(n14909), .ZN(
        n12962) );
  AOI221_X1 U5525 ( .B1(\registers[45][0] ), .B2(n16553), .C1(
        \registers[48][0] ), .C2(n16550), .A(n12473), .ZN(n12469) );
  OAI22_X1 U5526 ( .A1(n16547), .A2(n11951), .B1(n16544), .B2(n14888), .ZN(
        n12473) );
  AOI221_X1 U5527 ( .B1(\registers[5][0] ), .B2(n16502), .C1(
        \registers[59][0] ), .C2(n16499), .A(n12490), .ZN(n12485) );
  OAI22_X1 U5528 ( .A1(n16496), .A2(n12357), .B1(n16493), .B2(n14910), .ZN(
        n12490) );
  AOI221_X1 U5529 ( .B1(\registers[45][1] ), .B2(n16553), .C1(
        \registers[48][1] ), .C2(n16550), .A(n12290), .ZN(n12287) );
  OAI22_X1 U5530 ( .A1(n16547), .A2(n11952), .B1(n16544), .B2(n14889), .ZN(
        n12290) );
  AOI221_X1 U5531 ( .B1(\registers[5][1] ), .B2(n16502), .C1(
        \registers[59][1] ), .C2(n16499), .A(n12298), .ZN(n12295) );
  OAI22_X1 U5532 ( .A1(n16496), .A2(n12359), .B1(n16493), .B2(n14911), .ZN(
        n12298) );
  AOI221_X1 U5533 ( .B1(\registers[45][2] ), .B2(n16553), .C1(
        \registers[48][2] ), .C2(n16550), .A(n12137), .ZN(n12134) );
  OAI22_X1 U5534 ( .A1(n16547), .A2(n11995), .B1(n16544), .B2(n14890), .ZN(
        n12137) );
  AOI221_X1 U5535 ( .B1(\registers[5][2] ), .B2(n16502), .C1(
        \registers[59][2] ), .C2(n16499), .A(n12145), .ZN(n12142) );
  OAI22_X1 U5536 ( .A1(n16496), .A2(n12361), .B1(n16493), .B2(n14912), .ZN(
        n12145) );
  AOI221_X1 U5537 ( .B1(\registers[45][3] ), .B2(n16553), .C1(
        \registers[48][3] ), .C2(n16550), .A(n11984), .ZN(n11981) );
  OAI22_X1 U5538 ( .A1(n16547), .A2(n11905), .B1(n16544), .B2(n14861), .ZN(
        n11984) );
  AOI221_X1 U5539 ( .B1(\registers[5][3] ), .B2(n16502), .C1(
        \registers[59][3] ), .C2(n16499), .A(n11992), .ZN(n11989) );
  OAI22_X1 U5540 ( .A1(n16496), .A2(n12362), .B1(n16493), .B2(n14863), .ZN(
        n11992) );
  AOI221_X1 U5541 ( .B1(\registers[45][4] ), .B2(n16553), .C1(
        \registers[48][4] ), .C2(n16550), .A(n11831), .ZN(n11828) );
  OAI22_X1 U5542 ( .A1(n16547), .A2(n11997), .B1(n16544), .B2(n14891), .ZN(
        n11831) );
  AOI221_X1 U5543 ( .B1(\registers[5][4] ), .B2(n16502), .C1(
        \registers[59][4] ), .C2(n16499), .A(n11839), .ZN(n11836) );
  OAI22_X1 U5544 ( .A1(n16496), .A2(n12363), .B1(n16493), .B2(n14864), .ZN(
        n11839) );
  AOI221_X1 U5545 ( .B1(\registers[45][5] ), .B2(n16553), .C1(
        \registers[48][5] ), .C2(n16550), .A(n11788), .ZN(n11785) );
  OAI22_X1 U5546 ( .A1(n16547), .A2(n11906), .B1(n16544), .B2(n14862), .ZN(
        n11788) );
  AOI221_X1 U5547 ( .B1(\registers[5][5] ), .B2(n16502), .C1(
        \registers[59][5] ), .C2(n16499), .A(n11796), .ZN(n11793) );
  OAI22_X1 U5548 ( .A1(n16496), .A2(n12365), .B1(n16493), .B2(n14865), .ZN(
        n11796) );
  AOI221_X1 U5549 ( .B1(\registers[45][6] ), .B2(n16553), .C1(
        \registers[48][6] ), .C2(n16550), .A(n11745), .ZN(n11742) );
  OAI22_X1 U5550 ( .A1(n16547), .A2(n11998), .B1(n16544), .B2(n14892), .ZN(
        n11745) );
  AOI221_X1 U5551 ( .B1(\registers[5][6] ), .B2(n16502), .C1(
        \registers[59][6] ), .C2(n16499), .A(n11753), .ZN(n11750) );
  OAI22_X1 U5552 ( .A1(n16496), .A2(n12367), .B1(n16493), .B2(n14913), .ZN(
        n11753) );
  AOI221_X1 U5553 ( .B1(\registers[45][7] ), .B2(n16553), .C1(
        \registers[48][7] ), .C2(n16550), .A(n11702), .ZN(n11699) );
  OAI22_X1 U5554 ( .A1(n16547), .A2(n11999), .B1(n16544), .B2(n14893), .ZN(
        n11702) );
  AOI221_X1 U5555 ( .B1(\registers[5][7] ), .B2(n16502), .C1(
        \registers[59][7] ), .C2(n16499), .A(n11710), .ZN(n11707) );
  OAI22_X1 U5556 ( .A1(n16496), .A2(n12369), .B1(n16493), .B2(n14914), .ZN(
        n11710) );
  AOI221_X1 U5557 ( .B1(\registers[45][8] ), .B2(n16553), .C1(
        \registers[48][8] ), .C2(n16550), .A(n11659), .ZN(n11656) );
  OAI22_X1 U5558 ( .A1(n16547), .A2(n12000), .B1(n16544), .B2(n14894), .ZN(
        n11659) );
  AOI221_X1 U5559 ( .B1(\registers[5][8] ), .B2(n16502), .C1(
        \registers[59][8] ), .C2(n16499), .A(n11667), .ZN(n11664) );
  OAI22_X1 U5560 ( .A1(n16496), .A2(n12408), .B1(n16493), .B2(n14915), .ZN(
        n11667) );
  AOI221_X1 U5561 ( .B1(\registers[45][9] ), .B2(n16553), .C1(
        \registers[48][9] ), .C2(n16550), .A(n11616), .ZN(n11613) );
  OAI22_X1 U5562 ( .A1(n16547), .A2(n12001), .B1(n16544), .B2(n14895), .ZN(
        n11616) );
  AOI221_X1 U5563 ( .B1(\registers[5][9] ), .B2(n16502), .C1(
        \registers[59][9] ), .C2(n16499), .A(n11624), .ZN(n11621) );
  OAI22_X1 U5564 ( .A1(n16496), .A2(n12410), .B1(n16493), .B2(n14916), .ZN(
        n11624) );
  AOI221_X1 U5565 ( .B1(\registers[45][10] ), .B2(n16553), .C1(
        \registers[48][10] ), .C2(n16550), .A(n11573), .ZN(n11570) );
  OAI22_X1 U5566 ( .A1(n16547), .A2(n12002), .B1(n16544), .B2(n14896), .ZN(
        n11573) );
  AOI221_X1 U5567 ( .B1(\registers[5][10] ), .B2(n16502), .C1(
        \registers[59][10] ), .C2(n16499), .A(n11581), .ZN(n11578) );
  OAI22_X1 U5568 ( .A1(n16496), .A2(n12551), .B1(n16493), .B2(n14917), .ZN(
        n11581) );
  AOI221_X1 U5569 ( .B1(\registers[45][11] ), .B2(n16553), .C1(
        \registers[48][11] ), .C2(n16550), .A(n11530), .ZN(n11527) );
  OAI22_X1 U5570 ( .A1(n16547), .A2(n12003), .B1(n16544), .B2(n14897), .ZN(
        n11530) );
  AOI221_X1 U5571 ( .B1(\registers[5][11] ), .B2(n16502), .C1(
        \registers[59][11] ), .C2(n16499), .A(n11538), .ZN(n11535) );
  OAI22_X1 U5572 ( .A1(n16496), .A2(n12602), .B1(n16493), .B2(n14918), .ZN(
        n11538) );
  AOI221_X1 U5573 ( .B1(\registers[45][12] ), .B2(n16554), .C1(
        \registers[48][12] ), .C2(n16551), .A(n11487), .ZN(n11484) );
  OAI22_X1 U5574 ( .A1(n16548), .A2(n12004), .B1(n16545), .B2(n14898), .ZN(
        n11487) );
  AOI221_X1 U5575 ( .B1(\registers[5][12] ), .B2(n16503), .C1(
        \registers[59][12] ), .C2(n16500), .A(n11495), .ZN(n11492) );
  OAI22_X1 U5576 ( .A1(n16497), .A2(n12669), .B1(n16494), .B2(n14919), .ZN(
        n11495) );
  AOI221_X1 U5577 ( .B1(\registers[45][13] ), .B2(n16554), .C1(
        \registers[48][13] ), .C2(n16551), .A(n11443), .ZN(n11440) );
  OAI22_X1 U5578 ( .A1(n16548), .A2(n12005), .B1(n16545), .B2(n14899), .ZN(
        n11443) );
  AOI221_X1 U5579 ( .B1(\registers[5][13] ), .B2(n16503), .C1(
        \registers[59][13] ), .C2(n16500), .A(n11451), .ZN(n11448) );
  OAI22_X1 U5580 ( .A1(n16497), .A2(n13999), .B1(n16494), .B2(n14920), .ZN(
        n11451) );
  AOI221_X1 U5581 ( .B1(\registers[45][14] ), .B2(n16554), .C1(
        \registers[48][14] ), .C2(n16551), .A(n11400), .ZN(n11397) );
  OAI22_X1 U5582 ( .A1(n16548), .A2(n12006), .B1(n16545), .B2(n14900), .ZN(
        n11400) );
  AOI221_X1 U5583 ( .B1(\registers[5][14] ), .B2(n16503), .C1(
        \registers[59][14] ), .C2(n16500), .A(n11408), .ZN(n11405) );
  OAI22_X1 U5584 ( .A1(n16497), .A2(n14014), .B1(n16494), .B2(n14921), .ZN(
        n11408) );
  AOI221_X1 U5585 ( .B1(\registers[45][15] ), .B2(n16554), .C1(
        \registers[48][15] ), .C2(n16551), .A(n11357), .ZN(n11354) );
  OAI22_X1 U5586 ( .A1(n16548), .A2(n12007), .B1(n16545), .B2(n14901), .ZN(
        n11357) );
  AOI221_X1 U5587 ( .B1(\registers[5][15] ), .B2(n16503), .C1(
        \registers[59][15] ), .C2(n16500), .A(n11365), .ZN(n11362) );
  OAI22_X1 U5588 ( .A1(n16497), .A2(n14032), .B1(n16494), .B2(n14922), .ZN(
        n11365) );
  AOI221_X1 U5589 ( .B1(\registers[45][16] ), .B2(n16554), .C1(
        \registers[48][16] ), .C2(n16551), .A(n11314), .ZN(n11311) );
  OAI22_X1 U5590 ( .A1(n16548), .A2(n12008), .B1(n16545), .B2(n14902), .ZN(
        n11314) );
  AOI221_X1 U5591 ( .B1(\registers[5][16] ), .B2(n16503), .C1(
        \registers[59][16] ), .C2(n16500), .A(n11322), .ZN(n11319) );
  OAI22_X1 U5592 ( .A1(n16497), .A2(n14036), .B1(n16494), .B2(n14923), .ZN(
        n11322) );
  AOI221_X1 U5593 ( .B1(\registers[45][17] ), .B2(n16554), .C1(
        \registers[48][17] ), .C2(n16551), .A(n11271), .ZN(n11268) );
  OAI22_X1 U5594 ( .A1(n16548), .A2(n12009), .B1(n16545), .B2(n14903), .ZN(
        n11271) );
  AOI221_X1 U5595 ( .B1(\registers[5][17] ), .B2(n16503), .C1(
        \registers[59][17] ), .C2(n16500), .A(n11279), .ZN(n11276) );
  OAI22_X1 U5596 ( .A1(n16497), .A2(n14038), .B1(n16494), .B2(n14924), .ZN(
        n11279) );
  AOI221_X1 U5597 ( .B1(\registers[45][18] ), .B2(n16554), .C1(
        \registers[48][18] ), .C2(n16551), .A(n11228), .ZN(n11225) );
  OAI22_X1 U5598 ( .A1(n16548), .A2(n12010), .B1(n16545), .B2(n14904), .ZN(
        n11228) );
  AOI221_X1 U5599 ( .B1(\registers[5][18] ), .B2(n16503), .C1(
        \registers[59][18] ), .C2(n16500), .A(n11236), .ZN(n11233) );
  OAI22_X1 U5600 ( .A1(n16497), .A2(n14040), .B1(n16494), .B2(n14925), .ZN(
        n11236) );
  AOI221_X1 U5601 ( .B1(\registers[45][19] ), .B2(n16554), .C1(
        \registers[48][19] ), .C2(n16551), .A(n11185), .ZN(n11182) );
  OAI22_X1 U5602 ( .A1(n16548), .A2(n12011), .B1(n16545), .B2(n14905), .ZN(
        n11185) );
  AOI221_X1 U5603 ( .B1(\registers[5][19] ), .B2(n16503), .C1(
        \registers[59][19] ), .C2(n16500), .A(n11193), .ZN(n11190) );
  OAI22_X1 U5604 ( .A1(n16497), .A2(n14042), .B1(n16494), .B2(n14926), .ZN(
        n11193) );
  AOI221_X1 U5605 ( .B1(\registers[45][20] ), .B2(n16554), .C1(
        \registers[48][20] ), .C2(n16551), .A(n11142), .ZN(n11139) );
  OAI22_X1 U5606 ( .A1(n16548), .A2(n12012), .B1(n16545), .B2(n14906), .ZN(
        n11142) );
  AOI221_X1 U5607 ( .B1(\registers[5][20] ), .B2(n16503), .C1(
        \registers[59][20] ), .C2(n16500), .A(n11150), .ZN(n11147) );
  OAI22_X1 U5608 ( .A1(n16497), .A2(n14044), .B1(n16494), .B2(n14927), .ZN(
        n11150) );
  AOI221_X1 U5609 ( .B1(\registers[45][21] ), .B2(n16554), .C1(
        \registers[48][21] ), .C2(n16551), .A(n11099), .ZN(n11096) );
  OAI22_X1 U5610 ( .A1(n16548), .A2(n12013), .B1(n16545), .B2(n14907), .ZN(
        n11099) );
  AOI221_X1 U5611 ( .B1(\registers[5][21] ), .B2(n16503), .C1(
        \registers[59][21] ), .C2(n16500), .A(n11107), .ZN(n11104) );
  OAI22_X1 U5612 ( .A1(n16497), .A2(n14046), .B1(n16494), .B2(n14928), .ZN(
        n11107) );
  AOI221_X1 U5613 ( .B1(\registers[45][22] ), .B2(n16554), .C1(
        \registers[48][22] ), .C2(n16551), .A(n11056), .ZN(n11053) );
  OAI22_X1 U5614 ( .A1(n16548), .A2(n12014), .B1(n16545), .B2(n14908), .ZN(
        n11056) );
  AOI221_X1 U5615 ( .B1(\registers[5][22] ), .B2(n16503), .C1(
        \registers[59][22] ), .C2(n16500), .A(n11064), .ZN(n11061) );
  OAI22_X1 U5616 ( .A1(n16497), .A2(n14048), .B1(n16494), .B2(n14929), .ZN(
        n11064) );
  AOI221_X1 U5617 ( .B1(\registers[45][23] ), .B2(n16554), .C1(
        \registers[48][23] ), .C2(n16551), .A(n11013), .ZN(n11010) );
  OAI22_X1 U5618 ( .A1(n16548), .A2(n12015), .B1(n16545), .B2(n14909), .ZN(
        n11013) );
  AOI221_X1 U5619 ( .B1(\registers[5][23] ), .B2(n16503), .C1(
        \registers[59][23] ), .C2(n16500), .A(n11021), .ZN(n11018) );
  OAI22_X1 U5620 ( .A1(n16497), .A2(n14050), .B1(n16494), .B2(n14930), .ZN(
        n11021) );
  AOI221_X1 U5621 ( .B1(\registers[63][0] ), .B2(n17661), .C1(
        \registers[62][0] ), .C2(n17658), .A(n12404), .ZN(n12401) );
  OAI22_X1 U5622 ( .A1(n17655), .A2(n12357), .B1(n17652), .B2(n15326), .ZN(
        n12404) );
  AOI221_X1 U5623 ( .B1(\registers[11][0] ), .B2(n17805), .C1(net226849), .C2(
        n17802), .A(n12380), .ZN(n12377) );
  OAI22_X1 U5624 ( .A1(n17799), .A2(n15699), .B1(n17796), .B2(n11881), .ZN(
        n12380) );
  AOI221_X1 U5625 ( .B1(\registers[63][1] ), .B2(n17661), .C1(
        \registers[62][1] ), .C2(n17658), .A(n12250), .ZN(n12247) );
  OAI22_X1 U5626 ( .A1(n17655), .A2(n12359), .B1(n17652), .B2(n15327), .ZN(
        n12250) );
  AOI221_X1 U5627 ( .B1(\registers[11][1] ), .B2(n17805), .C1(net226863), .C2(
        n17802), .A(n12226), .ZN(n12223) );
  OAI22_X1 U5628 ( .A1(n17799), .A2(n15700), .B1(n17796), .B2(n11882), .ZN(
        n12226) );
  AOI221_X1 U5629 ( .B1(\registers[63][2] ), .B2(n17661), .C1(
        \registers[62][2] ), .C2(n17658), .A(n12095), .ZN(n12092) );
  OAI22_X1 U5630 ( .A1(n17655), .A2(n12361), .B1(n17652), .B2(n15328), .ZN(
        n12095) );
  AOI221_X1 U5631 ( .B1(\registers[11][2] ), .B2(n17805), .C1(net226890), .C2(
        n17802), .A(n12071), .ZN(n12068) );
  OAI22_X1 U5632 ( .A1(n17799), .A2(n15701), .B1(n17796), .B2(n11883), .ZN(
        n12071) );
  AOI221_X1 U5633 ( .B1(\registers[63][3] ), .B2(n17661), .C1(
        \registers[62][3] ), .C2(n17658), .A(n11942), .ZN(n11939) );
  OAI22_X1 U5634 ( .A1(n17655), .A2(n12362), .B1(n17652), .B2(n15329), .ZN(
        n11942) );
  AOI221_X1 U5635 ( .B1(\registers[11][3] ), .B2(n17805), .C1(net226901), .C2(
        n17802), .A(n11918), .ZN(n11915) );
  OAI22_X1 U5636 ( .A1(n17799), .A2(n15702), .B1(n17796), .B2(n11627), .ZN(
        n11918) );
  AOI221_X1 U5637 ( .B1(\registers[63][4] ), .B2(n17661), .C1(
        \registers[62][4] ), .C2(n17658), .A(n10499), .ZN(n10496) );
  OAI22_X1 U5638 ( .A1(n17655), .A2(n12363), .B1(n17652), .B2(n15330), .ZN(
        n10499) );
  AOI221_X1 U5639 ( .B1(\registers[11][4] ), .B2(n17805), .C1(net226974), .C2(
        n17802), .A(n10475), .ZN(n10472) );
  OAI22_X1 U5640 ( .A1(n17799), .A2(n15366), .B1(n17796), .B2(n11884), .ZN(
        n10475) );
  AOI221_X1 U5641 ( .B1(\registers[63][5] ), .B2(n17661), .C1(
        \registers[62][5] ), .C2(n17658), .A(n10389), .ZN(n10386) );
  OAI22_X1 U5642 ( .A1(n17655), .A2(n12365), .B1(n17652), .B2(n15331), .ZN(
        n10389) );
  AOI221_X1 U5643 ( .B1(\registers[11][5] ), .B2(n17805), .C1(net226994), .C2(
        n17802), .A(n10365), .ZN(n10362) );
  OAI22_X1 U5644 ( .A1(n17799), .A2(n15703), .B1(n17796), .B2(n11885), .ZN(
        n10365) );
  AOI221_X1 U5645 ( .B1(\registers[63][6] ), .B2(n17661), .C1(
        \registers[62][6] ), .C2(n17658), .A(n10277), .ZN(n10274) );
  OAI22_X1 U5646 ( .A1(n17655), .A2(n12367), .B1(n17652), .B2(n15332), .ZN(
        n10277) );
  AOI221_X1 U5647 ( .B1(\registers[11][6] ), .B2(n17805), .C1(net227018), .C2(
        n17802), .A(n10253), .ZN(n10250) );
  OAI22_X1 U5648 ( .A1(n17799), .A2(n15704), .B1(n17796), .B2(n11886), .ZN(
        n10253) );
  AOI221_X1 U5649 ( .B1(\registers[63][7] ), .B2(n17661), .C1(
        \registers[62][7] ), .C2(n17658), .A(n7641), .ZN(n7638) );
  OAI22_X1 U5650 ( .A1(n17655), .A2(n12369), .B1(n17652), .B2(n15333), .ZN(
        n7641) );
  AOI221_X1 U5651 ( .B1(\registers[11][7] ), .B2(n17805), .C1(net227036), .C2(
        n17802), .A(n7617), .ZN(n7614) );
  OAI22_X1 U5652 ( .A1(n17799), .A2(n15705), .B1(n17796), .B2(n11887), .ZN(
        n7617) );
  AOI221_X1 U5653 ( .B1(\registers[63][8] ), .B2(n17661), .C1(
        \registers[62][8] ), .C2(n17658), .A(n7526), .ZN(n7523) );
  OAI22_X1 U5654 ( .A1(n17655), .A2(n12408), .B1(n17652), .B2(n15334), .ZN(
        n7526) );
  AOI221_X1 U5655 ( .B1(\registers[11][8] ), .B2(n17805), .C1(net227054), .C2(
        n17802), .A(n7502), .ZN(n7499) );
  OAI22_X1 U5656 ( .A1(n17799), .A2(n15706), .B1(n17796), .B2(n11888), .ZN(
        n7502) );
  AOI221_X1 U5657 ( .B1(\registers[63][9] ), .B2(n17661), .C1(
        \registers[62][9] ), .C2(n17658), .A(n7417), .ZN(n7414) );
  OAI22_X1 U5658 ( .A1(n17655), .A2(n12410), .B1(n17652), .B2(n15335), .ZN(
        n7417) );
  AOI221_X1 U5659 ( .B1(\registers[11][9] ), .B2(n17805), .C1(net227072), .C2(
        n17802), .A(n7393), .ZN(n7390) );
  OAI22_X1 U5660 ( .A1(n17799), .A2(n15707), .B1(n17796), .B2(n11889), .ZN(
        n7393) );
  AOI221_X1 U5661 ( .B1(\registers[63][10] ), .B2(n17661), .C1(
        \registers[62][10] ), .C2(n17658), .A(n7308), .ZN(n7305) );
  OAI22_X1 U5662 ( .A1(n17655), .A2(n12551), .B1(n17652), .B2(n15336), .ZN(
        n7308) );
  AOI221_X1 U5663 ( .B1(\registers[11][10] ), .B2(n17805), .C1(net227090), 
        .C2(n17802), .A(n7284), .ZN(n7281) );
  OAI22_X1 U5664 ( .A1(n17799), .A2(n15708), .B1(n17796), .B2(n11890), .ZN(
        n7284) );
  AOI221_X1 U5665 ( .B1(\registers[63][11] ), .B2(n17662), .C1(
        \registers[62][11] ), .C2(n17659), .A(n7194), .ZN(n7191) );
  OAI22_X1 U5666 ( .A1(n17656), .A2(n12602), .B1(n17653), .B2(n15337), .ZN(
        n7194) );
  AOI221_X1 U5667 ( .B1(\registers[11][11] ), .B2(n17806), .C1(net227108), 
        .C2(n17803), .A(n7170), .ZN(n7167) );
  OAI22_X1 U5668 ( .A1(n17800), .A2(n15709), .B1(n17797), .B2(n11891), .ZN(
        n7170) );
  AOI221_X1 U5669 ( .B1(\registers[63][12] ), .B2(n17662), .C1(
        \registers[62][12] ), .C2(n17659), .A(n7085), .ZN(n7082) );
  OAI22_X1 U5670 ( .A1(n17656), .A2(n12669), .B1(n17653), .B2(n15338), .ZN(
        n7085) );
  AOI221_X1 U5671 ( .B1(\registers[11][12] ), .B2(n17806), .C1(net227126), 
        .C2(n17803), .A(n7061), .ZN(n7058) );
  OAI22_X1 U5672 ( .A1(n17800), .A2(n15710), .B1(n17797), .B2(n11892), .ZN(
        n7061) );
  AOI221_X1 U5673 ( .B1(\registers[63][13] ), .B2(n17662), .C1(
        \registers[62][13] ), .C2(n17659), .A(n6976), .ZN(n6973) );
  OAI22_X1 U5674 ( .A1(n17656), .A2(n13999), .B1(n17653), .B2(n15339), .ZN(
        n6976) );
  AOI221_X1 U5675 ( .B1(\registers[11][13] ), .B2(n17806), .C1(net227144), 
        .C2(n17803), .A(n6952), .ZN(n6949) );
  OAI22_X1 U5676 ( .A1(n17800), .A2(n15711), .B1(n17797), .B2(n11893), .ZN(
        n6952) );
  AOI221_X1 U5677 ( .B1(\registers[63][14] ), .B2(n17662), .C1(
        \registers[62][14] ), .C2(n17659), .A(n6867), .ZN(n6864) );
  OAI22_X1 U5678 ( .A1(n17656), .A2(n14014), .B1(n17653), .B2(n15340), .ZN(
        n6867) );
  AOI221_X1 U5679 ( .B1(\registers[11][14] ), .B2(n17806), .C1(net227162), 
        .C2(n17803), .A(n6843), .ZN(n6840) );
  OAI22_X1 U5680 ( .A1(n17800), .A2(n15712), .B1(n17797), .B2(n11894), .ZN(
        n6843) );
  AOI221_X1 U5681 ( .B1(\registers[63][15] ), .B2(n17662), .C1(
        \registers[62][15] ), .C2(n17659), .A(n6758), .ZN(n6755) );
  OAI22_X1 U5682 ( .A1(n17656), .A2(n14032), .B1(n17653), .B2(n15341), .ZN(
        n6758) );
  AOI221_X1 U5683 ( .B1(\registers[11][15] ), .B2(n17806), .C1(net227180), 
        .C2(n17803), .A(n6734), .ZN(n6731) );
  OAI22_X1 U5684 ( .A1(n17800), .A2(n15713), .B1(n17797), .B2(n11895), .ZN(
        n6734) );
  AOI221_X1 U5685 ( .B1(\registers[63][16] ), .B2(n17662), .C1(
        \registers[62][16] ), .C2(n17659), .A(n6618), .ZN(n6615) );
  OAI22_X1 U5686 ( .A1(n17656), .A2(n14036), .B1(n17653), .B2(n15342), .ZN(
        n6618) );
  AOI221_X1 U5687 ( .B1(\registers[11][16] ), .B2(n17806), .C1(net227198), 
        .C2(n17803), .A(n6574), .ZN(n6570) );
  OAI22_X1 U5688 ( .A1(n17800), .A2(n15714), .B1(n17797), .B2(n11896), .ZN(
        n6574) );
  AOI221_X1 U5689 ( .B1(\registers[63][17] ), .B2(n17662), .C1(
        \registers[62][17] ), .C2(n17659), .A(n6433), .ZN(n6428) );
  OAI22_X1 U5690 ( .A1(n17656), .A2(n14038), .B1(n17653), .B2(n15343), .ZN(
        n6433) );
  AOI221_X1 U5691 ( .B1(\registers[11][17] ), .B2(n17806), .C1(net227216), 
        .C2(n17803), .A(n6387), .ZN(n6384) );
  OAI22_X1 U5692 ( .A1(n17800), .A2(n15715), .B1(n17797), .B2(n11897), .ZN(
        n6387) );
  AOI221_X1 U5693 ( .B1(\registers[63][18] ), .B2(n17662), .C1(
        \registers[62][18] ), .C2(n17659), .A(n6247), .ZN(n6241) );
  OAI22_X1 U5694 ( .A1(n17656), .A2(n14040), .B1(n17653), .B2(n15344), .ZN(
        n6247) );
  AOI221_X1 U5695 ( .B1(\registers[11][18] ), .B2(n17806), .C1(net227234), 
        .C2(n17803), .A(n6202), .ZN(n6197) );
  OAI22_X1 U5696 ( .A1(n17800), .A2(n15716), .B1(n17797), .B2(n11898), .ZN(
        n6202) );
  AOI221_X1 U5697 ( .B1(\registers[63][19] ), .B2(n17662), .C1(
        \registers[62][19] ), .C2(n17659), .A(n6060), .ZN(n6056) );
  OAI22_X1 U5698 ( .A1(n17656), .A2(n14042), .B1(n17653), .B2(n15345), .ZN(
        n6060) );
  AOI221_X1 U5699 ( .B1(\registers[11][19] ), .B2(n17806), .C1(net227252), 
        .C2(n17803), .A(n6015), .ZN(n6010) );
  OAI22_X1 U5700 ( .A1(n17800), .A2(n15717), .B1(n17797), .B2(n11899), .ZN(
        n6015) );
  AOI221_X1 U5701 ( .B1(\registers[63][20] ), .B2(n17662), .C1(
        \registers[62][20] ), .C2(n17659), .A(n5873), .ZN(n5870) );
  OAI22_X1 U5702 ( .A1(n17656), .A2(n14044), .B1(n17653), .B2(n15346), .ZN(
        n5873) );
  AOI221_X1 U5703 ( .B1(\registers[11][20] ), .B2(n17806), .C1(net227270), 
        .C2(n17803), .A(n5843), .ZN(n5825) );
  OAI22_X1 U5704 ( .A1(n17800), .A2(n15718), .B1(n17797), .B2(n11900), .ZN(
        n5843) );
  AOI221_X1 U5705 ( .B1(\registers[63][21] ), .B2(n17662), .C1(
        \registers[62][21] ), .C2(n17659), .A(n5688), .ZN(n5683) );
  OAI22_X1 U5706 ( .A1(n17656), .A2(n14046), .B1(n17653), .B2(n15347), .ZN(
        n5688) );
  AOI221_X1 U5707 ( .B1(\registers[11][21] ), .B2(n17806), .C1(net227288), 
        .C2(n17803), .A(n5656), .ZN(n5653) );
  OAI22_X1 U5708 ( .A1(n17800), .A2(n15719), .B1(n17797), .B2(n11901), .ZN(
        n5656) );
  AOI221_X1 U5709 ( .B1(\registers[63][22] ), .B2(n17662), .C1(
        \registers[62][22] ), .C2(n17659), .A(n5502), .ZN(n5497) );
  OAI22_X1 U5710 ( .A1(n17656), .A2(n14048), .B1(n17653), .B2(n15348), .ZN(
        n5502) );
  AOI221_X1 U5711 ( .B1(\registers[11][22] ), .B2(n17806), .C1(net227306), 
        .C2(n17803), .A(n5469), .ZN(n5466) );
  OAI22_X1 U5712 ( .A1(n17800), .A2(n15720), .B1(n17797), .B2(n11902), .ZN(
        n5469) );
  AOI221_X1 U5713 ( .B1(\registers[63][31] ), .B2(n17661), .C1(
        \registers[62][31] ), .C2(n17658), .A(n14198), .ZN(n14189) );
  OAI22_X1 U5714 ( .A1(n17655), .A2(n12348), .B1(n17652), .B2(n15349), .ZN(
        n14198) );
  AOI221_X1 U5715 ( .B1(\registers[11][31] ), .B2(n17805), .C1(net227468), 
        .C2(n17802), .A(n14093), .ZN(n14082) );
  OAI22_X1 U5716 ( .A1(n17799), .A2(n15721), .B1(n17796), .B2(n11903), .ZN(
        n14093) );
  OAI22_X1 U5717 ( .A1(n7699), .A2(n17827), .B1(n4871), .B2(n17825), .ZN(n9701) );
  NOR4_X1 U5718 ( .A1(n4872), .A2(n4873), .A3(n4874), .A4(n4875), .ZN(n4871)
         );
  NAND4_X1 U5719 ( .A1(n4876), .A2(n4877), .A3(n4878), .A4(n4879), .ZN(n4875)
         );
  NAND4_X1 U5720 ( .A1(n4906), .A2(n4907), .A3(n4908), .A4(n4909), .ZN(n4872)
         );
  OAI22_X1 U5721 ( .A1(n7698), .A2(n17826), .B1(n4738), .B2(n17825), .ZN(n9773) );
  NOR4_X1 U5722 ( .A1(n4739), .A2(n4740), .A3(n4741), .A4(n4742), .ZN(n4738)
         );
  NAND4_X1 U5723 ( .A1(n4745), .A2(n4748), .A3(n4749), .A4(n4750), .ZN(n4742)
         );
  NAND4_X1 U5724 ( .A1(n4775), .A2(n4776), .A3(n4777), .A4(n4778), .ZN(n4739)
         );
  OAI22_X1 U5725 ( .A1(n7697), .A2(n17826), .B1(n4611), .B2(n17825), .ZN(n9845) );
  NOR4_X1 U5726 ( .A1(n4612), .A2(n4613), .A3(n4614), .A4(n4617), .ZN(n4611)
         );
  NAND4_X1 U5727 ( .A1(n4618), .A2(n4619), .A3(n4620), .A4(n4621), .ZN(n4617)
         );
  NAND4_X1 U5728 ( .A1(n4642), .A2(n4645), .A3(n4648), .A4(n4649), .ZN(n4612)
         );
  OAI22_X1 U5729 ( .A1(n7696), .A2(n17826), .B1(n4480), .B2(n17825), .ZN(n9917) );
  NOR4_X1 U5730 ( .A1(n4481), .A2(n4482), .A3(n4483), .A4(n4484), .ZN(n4480)
         );
  NAND4_X1 U5731 ( .A1(n4485), .A2(n4486), .A3(n4487), .A4(n4488), .ZN(n4484)
         );
  NAND4_X1 U5732 ( .A1(n4517), .A2(n4518), .A3(n4519), .A4(n4520), .ZN(n4481)
         );
  OAI22_X1 U5733 ( .A1(n7694), .A2(n17833), .B1(n14075), .B2(n17825), .ZN(
        n10061) );
  NOR4_X1 U5734 ( .A1(n14076), .A2(n14077), .A3(n14078), .A4(n14079), .ZN(
        n14075) );
  NAND4_X1 U5735 ( .A1(n14080), .A2(n14081), .A3(n14082), .A4(n14083), .ZN(
        n14079) );
  NAND4_X1 U5736 ( .A1(n14187), .A2(n14188), .A3(n14189), .A4(n14190), .ZN(
        n14076) );
  AOI211_X1 U5737 ( .C1(add_wr[4]), .C2(\sub_71/carry[4] ), .A(n14267), .B(
        n12514), .ZN(n14232) );
  NOR4_X1 U5738 ( .A1(n14213), .A2(N192), .A3(add_wr[4]), .A4(
        \sub_71/carry[4] ), .ZN(n14267) );
  AOI221_X1 U5739 ( .B1(\registers[47][24] ), .B2(n16291), .C1(
        \registers[51][24] ), .C2(n16288), .A(n12921), .ZN(n12916) );
  OAI22_X1 U5740 ( .A1(n16285), .A2(n15545), .B1(n16282), .B2(n14471), .ZN(
        n12921) );
  AOI221_X1 U5741 ( .B1(net227332), .B2(n16240), .C1(n16237), .C2(datain[24]), 
        .A(n12929), .ZN(n12924) );
  OAI22_X1 U5742 ( .A1(n16234), .A2(n15117), .B1(n16231), .B2(n14478), .ZN(
        n12929) );
  AOI221_X1 U5743 ( .B1(\registers[47][25] ), .B2(n16291), .C1(
        \registers[51][25] ), .C2(n16288), .A(n12879), .ZN(n12874) );
  OAI22_X1 U5744 ( .A1(n16285), .A2(n15546), .B1(n16282), .B2(n14472), .ZN(
        n12879) );
  AOI221_X1 U5745 ( .B1(net227350), .B2(n16240), .C1(n16237), .C2(datain[25]), 
        .A(n12887), .ZN(n12882) );
  OAI22_X1 U5746 ( .A1(n16234), .A2(n15118), .B1(n16231), .B2(n14479), .ZN(
        n12887) );
  AOI221_X1 U5747 ( .B1(\registers[47][26] ), .B2(n16291), .C1(
        \registers[51][26] ), .C2(n16288), .A(n12837), .ZN(n12832) );
  OAI22_X1 U5748 ( .A1(n16285), .A2(n15547), .B1(n16282), .B2(n14473), .ZN(
        n12837) );
  AOI221_X1 U5749 ( .B1(net227368), .B2(n16240), .C1(n16237), .C2(datain[26]), 
        .A(n12845), .ZN(n12840) );
  OAI22_X1 U5750 ( .A1(n16234), .A2(n15119), .B1(n16231), .B2(n14480), .ZN(
        n12845) );
  AOI221_X1 U5751 ( .B1(\registers[47][27] ), .B2(n16291), .C1(
        \registers[51][27] ), .C2(n16288), .A(n12795), .ZN(n12790) );
  OAI22_X1 U5752 ( .A1(n16285), .A2(n15548), .B1(n16282), .B2(n14474), .ZN(
        n12795) );
  AOI221_X1 U5753 ( .B1(net227386), .B2(n16240), .C1(n16237), .C2(datain[27]), 
        .A(n12803), .ZN(n12798) );
  OAI22_X1 U5754 ( .A1(n16234), .A2(n15120), .B1(n16231), .B2(n14481), .ZN(
        n12803) );
  AOI221_X1 U5755 ( .B1(\registers[47][28] ), .B2(n16291), .C1(
        \registers[51][28] ), .C2(n16288), .A(n12753), .ZN(n12748) );
  OAI22_X1 U5756 ( .A1(n16285), .A2(n15549), .B1(n16282), .B2(n14475), .ZN(
        n12753) );
  AOI221_X1 U5757 ( .B1(net227404), .B2(n16240), .C1(n16237), .C2(datain[28]), 
        .A(n12761), .ZN(n12756) );
  OAI22_X1 U5758 ( .A1(n16234), .A2(n15121), .B1(n16231), .B2(n14482), .ZN(
        n12761) );
  AOI221_X1 U5759 ( .B1(\registers[47][29] ), .B2(n16291), .C1(
        \registers[51][29] ), .C2(n16288), .A(n12711), .ZN(n12706) );
  OAI22_X1 U5760 ( .A1(n16285), .A2(n15550), .B1(n16282), .B2(n14476), .ZN(
        n12711) );
  AOI221_X1 U5761 ( .B1(net227422), .B2(n16240), .C1(n16237), .C2(datain[29]), 
        .A(n12719), .ZN(n12714) );
  OAI22_X1 U5762 ( .A1(n16234), .A2(n15122), .B1(n16231), .B2(n14483), .ZN(
        n12719) );
  AOI221_X1 U5763 ( .B1(\registers[47][30] ), .B2(n16291), .C1(
        \registers[51][30] ), .C2(n16288), .A(n12668), .ZN(n12663) );
  OAI22_X1 U5764 ( .A1(n16285), .A2(n15277), .B1(n16282), .B2(n14065), .ZN(
        n12668) );
  AOI221_X1 U5765 ( .B1(net227440), .B2(n16240), .C1(n16237), .C2(datain[30]), 
        .A(n12677), .ZN(n12672) );
  OAI22_X1 U5766 ( .A1(n16234), .A2(n14991), .B1(n16231), .B2(n14280), .ZN(
        n12677) );
  AOI221_X1 U5767 ( .B1(\registers[47][31] ), .B2(n16291), .C1(
        \registers[51][31] ), .C2(n16288), .A(n12598), .ZN(n12583) );
  OAI22_X1 U5768 ( .A1(n16285), .A2(n15551), .B1(n16282), .B2(n14477), .ZN(
        n12598) );
  AOI221_X1 U5769 ( .B1(net227458), .B2(n16240), .C1(n16237), .C2(datain[31]), 
        .A(n12625), .ZN(n12609) );
  OAI22_X1 U5770 ( .A1(n16234), .A2(n14992), .B1(n16231), .B2(n14281), .ZN(
        n12625) );
  AOI221_X1 U5771 ( .B1(\registers[49][24] ), .B2(n16543), .C1(
        \registers[51][24] ), .C2(n16540), .A(n10971), .ZN(n10966) );
  OAI22_X1 U5772 ( .A1(n16537), .A2(n15452), .B1(n16534), .B2(n14540), .ZN(
        n10971) );
  AOI221_X1 U5773 ( .B1(net227332), .B2(n16492), .C1(n16488), .C2(datain[24]), 
        .A(n10979), .ZN(n10974) );
  OAI22_X1 U5774 ( .A1(n16486), .A2(n15117), .B1(n16483), .B2(n14478), .ZN(
        n10979) );
  AOI221_X1 U5775 ( .B1(\registers[49][25] ), .B2(n16543), .C1(
        \registers[51][25] ), .C2(n16540), .A(n10928), .ZN(n10923) );
  OAI22_X1 U5776 ( .A1(n16537), .A2(n15453), .B1(n16534), .B2(n14541), .ZN(
        n10928) );
  AOI221_X1 U5777 ( .B1(net227350), .B2(n16492), .C1(n16488), .C2(datain[25]), 
        .A(n10936), .ZN(n10931) );
  OAI22_X1 U5778 ( .A1(n16486), .A2(n15118), .B1(n16483), .B2(n14479), .ZN(
        n10936) );
  AOI221_X1 U5779 ( .B1(\registers[49][26] ), .B2(n16543), .C1(
        \registers[51][26] ), .C2(n16540), .A(n10885), .ZN(n10880) );
  OAI22_X1 U5780 ( .A1(n16537), .A2(n15454), .B1(n16534), .B2(n14542), .ZN(
        n10885) );
  AOI221_X1 U5781 ( .B1(net227368), .B2(n16492), .C1(n16489), .C2(datain[26]), 
        .A(n10893), .ZN(n10888) );
  OAI22_X1 U5782 ( .A1(n16486), .A2(n15119), .B1(n16483), .B2(n14480), .ZN(
        n10893) );
  AOI221_X1 U5783 ( .B1(\registers[49][27] ), .B2(n16543), .C1(
        \registers[51][27] ), .C2(n16540), .A(n10842), .ZN(n10837) );
  OAI22_X1 U5784 ( .A1(n16537), .A2(n15455), .B1(n16534), .B2(n14543), .ZN(
        n10842) );
  AOI221_X1 U5785 ( .B1(net227386), .B2(n16492), .C1(n16489), .C2(datain[27]), 
        .A(n10850), .ZN(n10845) );
  OAI22_X1 U5786 ( .A1(n16486), .A2(n15120), .B1(n16483), .B2(n14481), .ZN(
        n10850) );
  AOI221_X1 U5787 ( .B1(\registers[49][28] ), .B2(n16543), .C1(
        \registers[51][28] ), .C2(n16540), .A(n10799), .ZN(n10794) );
  OAI22_X1 U5788 ( .A1(n16537), .A2(n15456), .B1(n16534), .B2(n14544), .ZN(
        n10799) );
  AOI221_X1 U5789 ( .B1(net227404), .B2(n16492), .C1(n16489), .C2(datain[28]), 
        .A(n10807), .ZN(n10802) );
  OAI22_X1 U5790 ( .A1(n16486), .A2(n15121), .B1(n16483), .B2(n14482), .ZN(
        n10807) );
  AOI221_X1 U5791 ( .B1(\registers[49][29] ), .B2(n16543), .C1(
        \registers[51][29] ), .C2(n16540), .A(n10756), .ZN(n10751) );
  OAI22_X1 U5792 ( .A1(n16537), .A2(n15457), .B1(n16534), .B2(n14545), .ZN(
        n10756) );
  AOI221_X1 U5793 ( .B1(net227422), .B2(n16492), .C1(n16489), .C2(datain[29]), 
        .A(n10764), .ZN(n10759) );
  OAI22_X1 U5794 ( .A1(n16486), .A2(n15122), .B1(n16483), .B2(n14483), .ZN(
        n10764) );
  AOI221_X1 U5795 ( .B1(\registers[49][30] ), .B2(n16543), .C1(
        \registers[51][30] ), .C2(n16540), .A(n10709), .ZN(n10701) );
  OAI22_X1 U5796 ( .A1(n16537), .A2(n15274), .B1(n16534), .B2(n14279), .ZN(
        n10709) );
  AOI221_X1 U5797 ( .B1(net227440), .B2(n16492), .C1(n16489), .C2(datain[30]), 
        .A(n10719), .ZN(n10714) );
  OAI22_X1 U5798 ( .A1(n16486), .A2(n14991), .B1(n16483), .B2(n14280), .ZN(
        n10719) );
  AOI221_X1 U5799 ( .B1(\registers[49][31] ), .B2(n16543), .C1(
        \registers[51][31] ), .C2(n16540), .A(n10616), .ZN(n10597) );
  OAI22_X1 U5800 ( .A1(n16537), .A2(n15458), .B1(n16534), .B2(n14546), .ZN(
        n10616) );
  AOI221_X1 U5801 ( .B1(net227458), .B2(n16492), .C1(n16489), .C2(datain[31]), 
        .A(n10650), .ZN(n10629) );
  OAI22_X1 U5802 ( .A1(n16486), .A2(n14992), .B1(n16483), .B2(n14281), .ZN(
        n10650) );
  AOI221_X1 U5803 ( .B1(net227322), .B2(n17747), .C1(\registers[29][23] ), 
        .C2(n17744), .A(n5294), .ZN(n5288) );
  OAI22_X1 U5804 ( .A1(n17741), .A2(n15722), .B1(n17738), .B2(n14757), .ZN(
        n5294) );
  AOI221_X1 U5805 ( .B1(net227325), .B2(n17699), .C1(\registers[9][23] ), .C2(
        n17696), .A(n5305), .ZN(n5299) );
  OAI22_X1 U5806 ( .A1(n17693), .A2(n15723), .B1(n17690), .B2(n12164), .ZN(
        n5305) );
  AOI221_X1 U5807 ( .B1(\registers[41][23] ), .B2(n17651), .C1(
        \registers[40][23] ), .C2(n17648), .A(n5316), .ZN(n5311) );
  OAI22_X1 U5808 ( .A1(n17645), .A2(n15459), .B1(n17642), .B2(n14758), .ZN(
        n5316) );
  AOI221_X1 U5809 ( .B1(\registers[18][23] ), .B2(n17795), .C1(
        \registers[19][23] ), .C2(n17792), .A(n5283), .ZN(n5278) );
  OAI22_X1 U5810 ( .A1(n17789), .A2(n14598), .B1(n17786), .B2(n15285), .ZN(
        n5283) );
  AOI221_X1 U5811 ( .B1(net227340), .B2(n17747), .C1(\registers[29][24] ), 
        .C2(n17744), .A(n5128), .ZN(n5121) );
  OAI22_X1 U5812 ( .A1(n17741), .A2(n15724), .B1(n17738), .B2(n14759), .ZN(
        n5128) );
  AOI221_X1 U5813 ( .B1(net227343), .B2(n17699), .C1(\registers[9][24] ), .C2(
        n17696), .A(n5136), .ZN(n5131) );
  OAI22_X1 U5814 ( .A1(n17693), .A2(n15725), .B1(n17690), .B2(n12165), .ZN(
        n5136) );
  AOI221_X1 U5815 ( .B1(\registers[41][24] ), .B2(n17651), .C1(
        \registers[40][24] ), .C2(n17648), .A(n5146), .ZN(n5139) );
  OAI22_X1 U5816 ( .A1(n17645), .A2(n15460), .B1(n17642), .B2(n14760), .ZN(
        n5146) );
  AOI221_X1 U5817 ( .B1(\registers[18][24] ), .B2(n17795), .C1(
        \registers[19][24] ), .C2(n17792), .A(n5118), .ZN(n5112) );
  OAI22_X1 U5818 ( .A1(n17789), .A2(n14599), .B1(n17786), .B2(n15286), .ZN(
        n5118) );
  AOI221_X1 U5819 ( .B1(net227358), .B2(n17747), .C1(\registers[29][25] ), 
        .C2(n17744), .A(n5012), .ZN(n5007) );
  OAI22_X1 U5820 ( .A1(n17741), .A2(n15726), .B1(n17738), .B2(n14761), .ZN(
        n5012) );
  AOI221_X1 U5821 ( .B1(net227361), .B2(n17699), .C1(\registers[9][25] ), .C2(
        n17696), .A(n5022), .ZN(n5015) );
  OAI22_X1 U5822 ( .A1(n17693), .A2(n15727), .B1(n17690), .B2(n12166), .ZN(
        n5022) );
  AOI221_X1 U5823 ( .B1(\registers[41][25] ), .B2(n17651), .C1(
        \registers[40][25] ), .C2(n17648), .A(n5030), .ZN(n5025) );
  OAI22_X1 U5824 ( .A1(n17645), .A2(n15461), .B1(n17642), .B2(n14762), .ZN(
        n5030) );
  AOI221_X1 U5825 ( .B1(\registers[18][25] ), .B2(n17795), .C1(
        \registers[19][25] ), .C2(n17792), .A(n5004), .ZN(n4999) );
  OAI22_X1 U5826 ( .A1(n17789), .A2(n14600), .B1(n17786), .B2(n15287), .ZN(
        n5004) );
  AOI221_X1 U5827 ( .B1(net227376), .B2(n17747), .C1(\registers[29][26] ), 
        .C2(n17744), .A(n4890), .ZN(n4885) );
  OAI22_X1 U5828 ( .A1(n17741), .A2(n15728), .B1(n17738), .B2(n14763), .ZN(
        n4890) );
  AOI221_X1 U5829 ( .B1(net227379), .B2(n17699), .C1(\registers[9][26] ), .C2(
        n17696), .A(n4902), .ZN(n4895) );
  OAI22_X1 U5830 ( .A1(n17693), .A2(n15729), .B1(n17690), .B2(n12167), .ZN(
        n4902) );
  AOI221_X1 U5831 ( .B1(\registers[41][26] ), .B2(n17651), .C1(
        \registers[40][26] ), .C2(n17648), .A(n4912), .ZN(n4907) );
  OAI22_X1 U5832 ( .A1(n17645), .A2(n15462), .B1(n17642), .B2(n14764), .ZN(
        n4912) );
  AOI221_X1 U5833 ( .B1(\registers[18][26] ), .B2(n17795), .C1(
        \registers[19][26] ), .C2(n17792), .A(n4882), .ZN(n4877) );
  OAI22_X1 U5834 ( .A1(n17789), .A2(n14601), .B1(n17786), .B2(n15288), .ZN(
        n4882) );
  AOI221_X1 U5835 ( .B1(net227394), .B2(n17747), .C1(\registers[29][27] ), 
        .C2(n17744), .A(n4763), .ZN(n4758) );
  OAI22_X1 U5836 ( .A1(n17741), .A2(n15730), .B1(n17738), .B2(n14765), .ZN(
        n4763) );
  AOI221_X1 U5837 ( .B1(net227397), .B2(n17699), .C1(\registers[9][27] ), .C2(
        n17696), .A(n4773), .ZN(n4768) );
  OAI22_X1 U5838 ( .A1(n17693), .A2(n15731), .B1(n17690), .B2(n12168), .ZN(
        n4773) );
  AOI221_X1 U5839 ( .B1(\registers[41][27] ), .B2(n17651), .C1(
        \registers[40][27] ), .C2(n17648), .A(n4781), .ZN(n4776) );
  OAI22_X1 U5840 ( .A1(n17645), .A2(n15463), .B1(n17642), .B2(n14766), .ZN(
        n4781) );
  AOI221_X1 U5841 ( .B1(\registers[18][27] ), .B2(n17795), .C1(
        \registers[19][27] ), .C2(n17792), .A(n4753), .ZN(n4748) );
  OAI22_X1 U5842 ( .A1(n17789), .A2(n14602), .B1(n17786), .B2(n15289), .ZN(
        n4753) );
  AOI221_X1 U5843 ( .B1(net227412), .B2(n17747), .C1(\registers[29][28] ), 
        .C2(n17744), .A(n4632), .ZN(n4627) );
  OAI22_X1 U5844 ( .A1(n17741), .A2(n15732), .B1(n17738), .B2(n14767), .ZN(
        n4632) );
  AOI221_X1 U5845 ( .B1(net227415), .B2(n17699), .C1(\registers[9][28] ), .C2(
        n17696), .A(n4640), .ZN(n4635) );
  OAI22_X1 U5846 ( .A1(n17693), .A2(n15733), .B1(n17690), .B2(n12169), .ZN(
        n4640) );
  AOI221_X1 U5847 ( .B1(\registers[41][28] ), .B2(n17651), .C1(
        \registers[40][28] ), .C2(n17648), .A(n4652), .ZN(n4645) );
  OAI22_X1 U5848 ( .A1(n17645), .A2(n15464), .B1(n17642), .B2(n14768), .ZN(
        n4652) );
  AOI221_X1 U5849 ( .B1(\registers[18][28] ), .B2(n17795), .C1(
        \registers[19][28] ), .C2(n17792), .A(n4624), .ZN(n4619) );
  OAI22_X1 U5850 ( .A1(n17789), .A2(n14603), .B1(n17786), .B2(n15290), .ZN(
        n4624) );
  AOI221_X1 U5851 ( .B1(net227430), .B2(n17747), .C1(\registers[29][29] ), 
        .C2(n17744), .A(n4503), .ZN(n4498) );
  OAI22_X1 U5852 ( .A1(n17741), .A2(n15734), .B1(n17738), .B2(n14769), .ZN(
        n4503) );
  AOI221_X1 U5853 ( .B1(net227433), .B2(n17699), .C1(\registers[9][29] ), .C2(
        n17696), .A(n4513), .ZN(n4508) );
  OAI22_X1 U5854 ( .A1(n17693), .A2(n15735), .B1(n17690), .B2(n12170), .ZN(
        n4513) );
  AOI221_X1 U5855 ( .B1(\registers[41][29] ), .B2(n17651), .C1(
        \registers[40][29] ), .C2(n17648), .A(n4523), .ZN(n4518) );
  OAI22_X1 U5856 ( .A1(n17645), .A2(n15465), .B1(n17642), .B2(n14770), .ZN(
        n4523) );
  AOI221_X1 U5857 ( .B1(\registers[18][29] ), .B2(n17795), .C1(
        \registers[19][29] ), .C2(n17792), .A(n4491), .ZN(n4486) );
  OAI22_X1 U5858 ( .A1(n17789), .A2(n14604), .B1(n17786), .B2(n15291), .ZN(
        n4491) );
  AOI221_X1 U5859 ( .B1(net227448), .B2(n17747), .C1(\registers[29][30] ), 
        .C2(n17744), .A(n4163), .ZN(n4138) );
  OAI22_X1 U5860 ( .A1(n17741), .A2(n15282), .B1(n17738), .B2(n14630), .ZN(
        n4163) );
  AOI221_X1 U5861 ( .B1(net227451), .B2(n17699), .C1(\registers[9][30] ), .C2(
        n17696), .A(n4199), .ZN(n4178) );
  OAI22_X1 U5862 ( .A1(n17693), .A2(n15283), .B1(n17690), .B2(n12160), .ZN(
        n4199) );
  AOI221_X1 U5863 ( .B1(\registers[41][30] ), .B2(n17651), .C1(
        \registers[40][30] ), .C2(n17648), .A(n4234), .ZN(n4214) );
  OAI22_X1 U5864 ( .A1(n17645), .A2(n15275), .B1(n17642), .B2(n14631), .ZN(
        n4234) );
  AOI221_X1 U5865 ( .B1(\registers[18][30] ), .B2(n17795), .C1(
        \registers[19][30] ), .C2(n17792), .A(n4125), .ZN(n4102) );
  OAI22_X1 U5866 ( .A1(n17789), .A2(n14299), .B1(n17786), .B2(n15270), .ZN(
        n4125) );
  AOI221_X1 U5867 ( .B1(\registers[47][0] ), .B2(n16289), .C1(
        \registers[51][0] ), .C2(n16286), .A(n13956), .ZN(n13949) );
  OAI22_X1 U5868 ( .A1(n16283), .A2(n15552), .B1(n16280), .B2(n14484), .ZN(
        n13956) );
  AOI221_X1 U5869 ( .B1(net226844), .B2(n16238), .C1(n16235), .C2(datain[0]), 
        .A(n13972), .ZN(n13965) );
  OAI22_X1 U5870 ( .A1(n16232), .A2(n15123), .B1(n16229), .B2(n14506), .ZN(
        n13972) );
  AOI221_X1 U5871 ( .B1(\registers[47][1] ), .B2(n16289), .C1(
        \registers[51][1] ), .C2(n16286), .A(n13887), .ZN(n13882) );
  OAI22_X1 U5872 ( .A1(n16283), .A2(n15553), .B1(n16280), .B2(n14485), .ZN(
        n13887) );
  AOI221_X1 U5873 ( .B1(net226857), .B2(n16238), .C1(n16235), .C2(datain[1]), 
        .A(n13895), .ZN(n13890) );
  OAI22_X1 U5874 ( .A1(n16232), .A2(n15124), .B1(n16229), .B2(n14507), .ZN(
        n13895) );
  AOI221_X1 U5875 ( .B1(\registers[47][2] ), .B2(n16289), .C1(
        \registers[51][2] ), .C2(n16286), .A(n13845), .ZN(n13840) );
  OAI22_X1 U5876 ( .A1(n16283), .A2(n15554), .B1(n16280), .B2(n14486), .ZN(
        n13845) );
  AOI221_X1 U5877 ( .B1(net226884), .B2(n16238), .C1(n16235), .C2(datain[2]), 
        .A(n13853), .ZN(n13848) );
  OAI22_X1 U5878 ( .A1(n16232), .A2(n15125), .B1(n16229), .B2(n14508), .ZN(
        n13853) );
  AOI221_X1 U5879 ( .B1(\registers[47][3] ), .B2(n16289), .C1(
        \registers[51][3] ), .C2(n16286), .A(n13803), .ZN(n13798) );
  OAI22_X1 U5880 ( .A1(n16283), .A2(n15555), .B1(n16280), .B2(n14487), .ZN(
        n13803) );
  AOI221_X1 U5881 ( .B1(net226904), .B2(n16238), .C1(n16235), .C2(datain[3]), 
        .A(n13811), .ZN(n13806) );
  OAI22_X1 U5882 ( .A1(n16232), .A2(n14997), .B1(n16229), .B2(n14296), .ZN(
        n13811) );
  AOI221_X1 U5883 ( .B1(\registers[47][4] ), .B2(n16289), .C1(
        \registers[51][4] ), .C2(n16286), .A(n13761), .ZN(n13756) );
  OAI22_X1 U5884 ( .A1(n16283), .A2(n15359), .B1(n16280), .B2(n14294), .ZN(
        n13761) );
  AOI221_X1 U5885 ( .B1(net226977), .B2(n16238), .C1(n16235), .C2(datain[4]), 
        .A(n13769), .ZN(n13764) );
  OAI22_X1 U5886 ( .A1(n16232), .A2(n14998), .B1(n16229), .B2(n14297), .ZN(
        n13769) );
  AOI221_X1 U5887 ( .B1(\registers[47][5] ), .B2(n16289), .C1(
        \registers[51][5] ), .C2(n16286), .A(n13719), .ZN(n13714) );
  OAI22_X1 U5888 ( .A1(n16283), .A2(n15360), .B1(n16280), .B2(n14295), .ZN(
        n13719) );
  AOI221_X1 U5889 ( .B1(net226997), .B2(n16238), .C1(n16235), .C2(datain[5]), 
        .A(n13727), .ZN(n13722) );
  OAI22_X1 U5890 ( .A1(n16232), .A2(n14999), .B1(n16229), .B2(n14298), .ZN(
        n13727) );
  AOI221_X1 U5891 ( .B1(\registers[47][6] ), .B2(n16289), .C1(
        \registers[51][6] ), .C2(n16286), .A(n13677), .ZN(n13672) );
  OAI22_X1 U5892 ( .A1(n16283), .A2(n15556), .B1(n16280), .B2(n14488), .ZN(
        n13677) );
  AOI221_X1 U5893 ( .B1(net227008), .B2(n16238), .C1(n16235), .C2(datain[6]), 
        .A(n13685), .ZN(n13680) );
  OAI22_X1 U5894 ( .A1(n16232), .A2(n15126), .B1(n16229), .B2(n14509), .ZN(
        n13685) );
  AOI221_X1 U5895 ( .B1(\registers[47][7] ), .B2(n16289), .C1(
        \registers[51][7] ), .C2(n16286), .A(n13635), .ZN(n13630) );
  OAI22_X1 U5896 ( .A1(n16283), .A2(n15557), .B1(n16280), .B2(n14489), .ZN(
        n13635) );
  AOI221_X1 U5897 ( .B1(net227026), .B2(n16238), .C1(n16235), .C2(datain[7]), 
        .A(n13643), .ZN(n13638) );
  OAI22_X1 U5898 ( .A1(n16232), .A2(n15127), .B1(n16229), .B2(n14510), .ZN(
        n13643) );
  AOI221_X1 U5899 ( .B1(\registers[47][8] ), .B2(n16289), .C1(
        \registers[51][8] ), .C2(n16286), .A(n13593), .ZN(n13588) );
  OAI22_X1 U5900 ( .A1(n16283), .A2(n15558), .B1(n16280), .B2(n14490), .ZN(
        n13593) );
  AOI221_X1 U5901 ( .B1(net227044), .B2(n16238), .C1(n16235), .C2(datain[8]), 
        .A(n13601), .ZN(n13596) );
  OAI22_X1 U5902 ( .A1(n16232), .A2(n15128), .B1(n16229), .B2(n14511), .ZN(
        n13601) );
  AOI221_X1 U5903 ( .B1(\registers[47][9] ), .B2(n16289), .C1(
        \registers[51][9] ), .C2(n16286), .A(n13551), .ZN(n13546) );
  OAI22_X1 U5904 ( .A1(n16283), .A2(n15559), .B1(n16280), .B2(n14491), .ZN(
        n13551) );
  AOI221_X1 U5905 ( .B1(net227062), .B2(n16238), .C1(n16235), .C2(datain[9]), 
        .A(n13559), .ZN(n13554) );
  OAI22_X1 U5906 ( .A1(n16232), .A2(n15129), .B1(n16229), .B2(n14512), .ZN(
        n13559) );
  AOI221_X1 U5907 ( .B1(\registers[47][10] ), .B2(n16289), .C1(
        \registers[51][10] ), .C2(n16286), .A(n13509), .ZN(n13504) );
  OAI22_X1 U5908 ( .A1(n16283), .A2(n15560), .B1(n16280), .B2(n14492), .ZN(
        n13509) );
  AOI221_X1 U5909 ( .B1(net227080), .B2(n16238), .C1(n16235), .C2(datain[10]), 
        .A(n13517), .ZN(n13512) );
  OAI22_X1 U5910 ( .A1(n16232), .A2(n15130), .B1(n16229), .B2(n14513), .ZN(
        n13517) );
  AOI221_X1 U5911 ( .B1(\registers[47][11] ), .B2(n16289), .C1(
        \registers[51][11] ), .C2(n16286), .A(n13467), .ZN(n13462) );
  OAI22_X1 U5912 ( .A1(n16283), .A2(n15561), .B1(n16280), .B2(n14493), .ZN(
        n13467) );
  AOI221_X1 U5913 ( .B1(net227098), .B2(n16238), .C1(n16235), .C2(datain[11]), 
        .A(n13475), .ZN(n13470) );
  OAI22_X1 U5914 ( .A1(n16232), .A2(n15131), .B1(n16229), .B2(n14514), .ZN(
        n13475) );
  AOI221_X1 U5915 ( .B1(\registers[47][12] ), .B2(n16290), .C1(
        \registers[51][12] ), .C2(n16287), .A(n13425), .ZN(n13420) );
  OAI22_X1 U5916 ( .A1(n16284), .A2(n15562), .B1(n16281), .B2(n14494), .ZN(
        n13425) );
  AOI221_X1 U5917 ( .B1(net227116), .B2(n16239), .C1(n16236), .C2(datain[12]), 
        .A(n13433), .ZN(n13428) );
  OAI22_X1 U5918 ( .A1(n16233), .A2(n15132), .B1(n16230), .B2(n14515), .ZN(
        n13433) );
  AOI221_X1 U5919 ( .B1(\registers[47][13] ), .B2(n16290), .C1(
        \registers[51][13] ), .C2(n16287), .A(n13383), .ZN(n13378) );
  OAI22_X1 U5920 ( .A1(n16284), .A2(n15563), .B1(n16281), .B2(n14495), .ZN(
        n13383) );
  AOI221_X1 U5921 ( .B1(net227134), .B2(n16239), .C1(n16236), .C2(datain[13]), 
        .A(n13391), .ZN(n13386) );
  OAI22_X1 U5922 ( .A1(n16233), .A2(n15133), .B1(n16230), .B2(n14516), .ZN(
        n13391) );
  AOI221_X1 U5923 ( .B1(\registers[47][14] ), .B2(n16290), .C1(
        \registers[51][14] ), .C2(n16287), .A(n13341), .ZN(n13336) );
  OAI22_X1 U5924 ( .A1(n16284), .A2(n15564), .B1(n16281), .B2(n14496), .ZN(
        n13341) );
  AOI221_X1 U5925 ( .B1(net227152), .B2(n16239), .C1(n16236), .C2(datain[14]), 
        .A(n13349), .ZN(n13344) );
  OAI22_X1 U5926 ( .A1(n16233), .A2(n15134), .B1(n16230), .B2(n14517), .ZN(
        n13349) );
  AOI221_X1 U5927 ( .B1(\registers[47][15] ), .B2(n16290), .C1(
        \registers[51][15] ), .C2(n16287), .A(n13299), .ZN(n13294) );
  OAI22_X1 U5928 ( .A1(n16284), .A2(n15565), .B1(n16281), .B2(n14497), .ZN(
        n13299) );
  AOI221_X1 U5929 ( .B1(net227170), .B2(n16239), .C1(n16236), .C2(datain[15]), 
        .A(n13307), .ZN(n13302) );
  OAI22_X1 U5930 ( .A1(n16233), .A2(n15135), .B1(n16230), .B2(n14518), .ZN(
        n13307) );
  AOI221_X1 U5931 ( .B1(\registers[47][16] ), .B2(n16290), .C1(
        \registers[51][16] ), .C2(n16287), .A(n13257), .ZN(n13252) );
  OAI22_X1 U5932 ( .A1(n16284), .A2(n15566), .B1(n16281), .B2(n14498), .ZN(
        n13257) );
  AOI221_X1 U5933 ( .B1(net227188), .B2(n16239), .C1(n16236), .C2(datain[16]), 
        .A(n13265), .ZN(n13260) );
  OAI22_X1 U5934 ( .A1(n16233), .A2(n15136), .B1(n16230), .B2(n14519), .ZN(
        n13265) );
  AOI221_X1 U5935 ( .B1(\registers[47][17] ), .B2(n16290), .C1(
        \registers[51][17] ), .C2(n16287), .A(n13215), .ZN(n13210) );
  OAI22_X1 U5936 ( .A1(n16284), .A2(n15567), .B1(n16281), .B2(n14499), .ZN(
        n13215) );
  AOI221_X1 U5937 ( .B1(net227206), .B2(n16239), .C1(n16236), .C2(datain[17]), 
        .A(n13223), .ZN(n13218) );
  OAI22_X1 U5938 ( .A1(n16233), .A2(n15137), .B1(n16230), .B2(n14520), .ZN(
        n13223) );
  AOI221_X1 U5939 ( .B1(\registers[47][18] ), .B2(n16290), .C1(
        \registers[51][18] ), .C2(n16287), .A(n13173), .ZN(n13168) );
  OAI22_X1 U5940 ( .A1(n16284), .A2(n15568), .B1(n16281), .B2(n14500), .ZN(
        n13173) );
  AOI221_X1 U5941 ( .B1(net227224), .B2(n16239), .C1(n16236), .C2(datain[18]), 
        .A(n13181), .ZN(n13176) );
  OAI22_X1 U5942 ( .A1(n16233), .A2(n15138), .B1(n16230), .B2(n14521), .ZN(
        n13181) );
  AOI221_X1 U5943 ( .B1(\registers[47][19] ), .B2(n16290), .C1(
        \registers[51][19] ), .C2(n16287), .A(n13131), .ZN(n13126) );
  OAI22_X1 U5944 ( .A1(n16284), .A2(n15569), .B1(n16281), .B2(n14501), .ZN(
        n13131) );
  AOI221_X1 U5945 ( .B1(net227242), .B2(n16239), .C1(n16236), .C2(datain[19]), 
        .A(n13139), .ZN(n13134) );
  OAI22_X1 U5946 ( .A1(n16233), .A2(n15139), .B1(n16230), .B2(n14522), .ZN(
        n13139) );
  AOI221_X1 U5947 ( .B1(\registers[47][20] ), .B2(n16290), .C1(
        \registers[51][20] ), .C2(n16287), .A(n13089), .ZN(n13084) );
  OAI22_X1 U5948 ( .A1(n16284), .A2(n15570), .B1(n16281), .B2(n14502), .ZN(
        n13089) );
  AOI221_X1 U5949 ( .B1(net227260), .B2(n16239), .C1(n16236), .C2(datain[20]), 
        .A(n13097), .ZN(n13092) );
  OAI22_X1 U5950 ( .A1(n16233), .A2(n15140), .B1(n16230), .B2(n14523), .ZN(
        n13097) );
  AOI221_X1 U5951 ( .B1(\registers[47][21] ), .B2(n16290), .C1(
        \registers[51][21] ), .C2(n16287), .A(n13047), .ZN(n13042) );
  OAI22_X1 U5952 ( .A1(n16284), .A2(n15571), .B1(n16281), .B2(n14503), .ZN(
        n13047) );
  AOI221_X1 U5953 ( .B1(net227278), .B2(n16239), .C1(n16236), .C2(datain[21]), 
        .A(n13055), .ZN(n13050) );
  OAI22_X1 U5954 ( .A1(n16233), .A2(n15141), .B1(n16230), .B2(n14524), .ZN(
        n13055) );
  AOI221_X1 U5955 ( .B1(\registers[47][22] ), .B2(n16290), .C1(
        \registers[51][22] ), .C2(n16287), .A(n13005), .ZN(n13000) );
  OAI22_X1 U5956 ( .A1(n16284), .A2(n15572), .B1(n16281), .B2(n14504), .ZN(
        n13005) );
  AOI221_X1 U5957 ( .B1(net227296), .B2(n16239), .C1(n16236), .C2(datain[22]), 
        .A(n13013), .ZN(n13008) );
  OAI22_X1 U5958 ( .A1(n16233), .A2(n15142), .B1(n16230), .B2(n14525), .ZN(
        n13013) );
  AOI221_X1 U5959 ( .B1(\registers[47][23] ), .B2(n16290), .C1(
        \registers[51][23] ), .C2(n16287), .A(n12963), .ZN(n12958) );
  OAI22_X1 U5960 ( .A1(n16284), .A2(n15573), .B1(n16281), .B2(n14505), .ZN(
        n12963) );
  AOI221_X1 U5961 ( .B1(net227314), .B2(n16239), .C1(n16236), .C2(datain[23]), 
        .A(n12971), .ZN(n12966) );
  OAI22_X1 U5962 ( .A1(n16233), .A2(n15143), .B1(n16230), .B2(n14526), .ZN(
        n12971) );
  AOI221_X1 U5963 ( .B1(net226844), .B2(n16490), .C1(datain[0]), .C2(n16487), 
        .A(n12491), .ZN(n12484) );
  OAI22_X1 U5964 ( .A1(n16484), .A2(n15123), .B1(n16481), .B2(n14506), .ZN(
        n12491) );
  AOI221_X1 U5965 ( .B1(net226857), .B2(n16490), .C1(datain[1]), .C2(n16487), 
        .A(n12299), .ZN(n12294) );
  OAI22_X1 U5966 ( .A1(n16484), .A2(n15124), .B1(n16481), .B2(n14507), .ZN(
        n12299) );
  AOI221_X1 U5967 ( .B1(net226884), .B2(n16490), .C1(datain[2]), .C2(n16487), 
        .A(n12146), .ZN(n12141) );
  OAI22_X1 U5968 ( .A1(n16484), .A2(n15125), .B1(n16481), .B2(n14508), .ZN(
        n12146) );
  AOI221_X1 U5969 ( .B1(net226904), .B2(n16490), .C1(datain[3]), .C2(n16487), 
        .A(n11993), .ZN(n11988) );
  OAI22_X1 U5970 ( .A1(n16484), .A2(n14997), .B1(n16481), .B2(n14296), .ZN(
        n11993) );
  AOI221_X1 U5971 ( .B1(net226977), .B2(n16490), .C1(n16487), .C2(datain[4]), 
        .A(n11840), .ZN(n11835) );
  OAI22_X1 U5972 ( .A1(n16484), .A2(n14998), .B1(n16481), .B2(n14297), .ZN(
        n11840) );
  AOI221_X1 U5973 ( .B1(net226997), .B2(n16490), .C1(n16487), .C2(datain[5]), 
        .A(n11797), .ZN(n11792) );
  OAI22_X1 U5974 ( .A1(n16484), .A2(n14999), .B1(n16481), .B2(n14298), .ZN(
        n11797) );
  AOI221_X1 U5975 ( .B1(net227008), .B2(n16490), .C1(n16487), .C2(datain[6]), 
        .A(n11754), .ZN(n11749) );
  OAI22_X1 U5976 ( .A1(n16484), .A2(n15126), .B1(n16481), .B2(n14509), .ZN(
        n11754) );
  AOI221_X1 U5977 ( .B1(net227026), .B2(n16490), .C1(n16487), .C2(datain[7]), 
        .A(n11711), .ZN(n11706) );
  OAI22_X1 U5978 ( .A1(n16484), .A2(n15127), .B1(n16481), .B2(n14510), .ZN(
        n11711) );
  AOI221_X1 U5979 ( .B1(net227044), .B2(n16490), .C1(n16487), .C2(datain[8]), 
        .A(n11668), .ZN(n11663) );
  OAI22_X1 U5980 ( .A1(n16484), .A2(n15128), .B1(n16481), .B2(n14511), .ZN(
        n11668) );
  AOI221_X1 U5981 ( .B1(net227062), .B2(n16490), .C1(n16487), .C2(datain[9]), 
        .A(n11625), .ZN(n11620) );
  OAI22_X1 U5982 ( .A1(n16484), .A2(n15129), .B1(n16481), .B2(n14512), .ZN(
        n11625) );
  AOI221_X1 U5983 ( .B1(net227080), .B2(n16490), .C1(n16487), .C2(datain[10]), 
        .A(n11582), .ZN(n11577) );
  OAI22_X1 U5984 ( .A1(n16484), .A2(n15130), .B1(n16481), .B2(n14513), .ZN(
        n11582) );
  AOI221_X1 U5985 ( .B1(net227098), .B2(n16490), .C1(n16487), .C2(datain[11]), 
        .A(n11539), .ZN(n11534) );
  OAI22_X1 U5986 ( .A1(n16484), .A2(n15131), .B1(n16481), .B2(n14514), .ZN(
        n11539) );
  AOI221_X1 U5987 ( .B1(net227116), .B2(n16491), .C1(n16487), .C2(datain[12]), 
        .A(n11496), .ZN(n11491) );
  OAI22_X1 U5988 ( .A1(n16485), .A2(n15132), .B1(n16482), .B2(n14515), .ZN(
        n11496) );
  AOI221_X1 U5989 ( .B1(net227134), .B2(n16491), .C1(n16488), .C2(datain[13]), 
        .A(n11452), .ZN(n11447) );
  OAI22_X1 U5990 ( .A1(n16485), .A2(n15133), .B1(n16482), .B2(n14516), .ZN(
        n11452) );
  AOI221_X1 U5991 ( .B1(net227152), .B2(n16491), .C1(n16488), .C2(datain[14]), 
        .A(n11409), .ZN(n11404) );
  OAI22_X1 U5992 ( .A1(n16485), .A2(n15134), .B1(n16482), .B2(n14517), .ZN(
        n11409) );
  AOI221_X1 U5993 ( .B1(net227170), .B2(n16491), .C1(n16488), .C2(datain[15]), 
        .A(n11366), .ZN(n11361) );
  OAI22_X1 U5994 ( .A1(n16485), .A2(n15135), .B1(n16482), .B2(n14518), .ZN(
        n11366) );
  AOI221_X1 U5995 ( .B1(net227188), .B2(n16491), .C1(n16488), .C2(datain[16]), 
        .A(n11323), .ZN(n11318) );
  OAI22_X1 U5996 ( .A1(n16485), .A2(n15136), .B1(n16482), .B2(n14519), .ZN(
        n11323) );
  AOI221_X1 U5997 ( .B1(net227206), .B2(n16491), .C1(n16488), .C2(datain[17]), 
        .A(n11280), .ZN(n11275) );
  OAI22_X1 U5998 ( .A1(n16485), .A2(n15137), .B1(n16482), .B2(n14520), .ZN(
        n11280) );
  AOI221_X1 U5999 ( .B1(net227224), .B2(n16491), .C1(n16488), .C2(datain[18]), 
        .A(n11237), .ZN(n11232) );
  OAI22_X1 U6000 ( .A1(n16485), .A2(n15138), .B1(n16482), .B2(n14521), .ZN(
        n11237) );
  AOI221_X1 U6001 ( .B1(net227242), .B2(n16491), .C1(n16488), .C2(datain[19]), 
        .A(n11194), .ZN(n11189) );
  OAI22_X1 U6002 ( .A1(n16485), .A2(n15139), .B1(n16482), .B2(n14522), .ZN(
        n11194) );
  AOI221_X1 U6003 ( .B1(net227260), .B2(n16491), .C1(n16488), .C2(datain[20]), 
        .A(n11151), .ZN(n11146) );
  OAI22_X1 U6004 ( .A1(n16485), .A2(n15140), .B1(n16482), .B2(n14523), .ZN(
        n11151) );
  AOI221_X1 U6005 ( .B1(net227278), .B2(n16491), .C1(n16488), .C2(datain[21]), 
        .A(n11108), .ZN(n11103) );
  OAI22_X1 U6006 ( .A1(n16485), .A2(n15141), .B1(n16482), .B2(n14524), .ZN(
        n11108) );
  AOI221_X1 U6007 ( .B1(net227296), .B2(n16491), .C1(n16488), .C2(datain[22]), 
        .A(n11065), .ZN(n11060) );
  OAI22_X1 U6008 ( .A1(n16485), .A2(n15142), .B1(n16482), .B2(n14525), .ZN(
        n11065) );
  AOI221_X1 U6009 ( .B1(net227314), .B2(n16491), .C1(n16488), .C2(datain[23]), 
        .A(n11022), .ZN(n11017) );
  OAI22_X1 U6010 ( .A1(n16485), .A2(n15143), .B1(n16482), .B2(n14526), .ZN(
        n11022) );
  AOI221_X1 U6011 ( .B1(net226839), .B2(n17745), .C1(\registers[29][0] ), .C2(
        n17742), .A(n12389), .ZN(n12384) );
  OAI22_X1 U6012 ( .A1(n17739), .A2(n15736), .B1(n17736), .B2(n14771), .ZN(
        n12389) );
  AOI221_X1 U6013 ( .B1(\registers[41][0] ), .B2(n17649), .C1(
        \registers[40][0] ), .C2(n17646), .A(n12405), .ZN(n12400) );
  OAI22_X1 U6014 ( .A1(n17643), .A2(n15466), .B1(n17640), .B2(n14772), .ZN(
        n12405) );
  AOI221_X1 U6015 ( .B1(\registers[18][0] ), .B2(n17793), .C1(
        \registers[19][0] ), .C2(n17790), .A(n12381), .ZN(n12376) );
  OAI22_X1 U6016 ( .A1(n17787), .A2(n14605), .B1(n17784), .B2(n15292), .ZN(
        n12381) );
  AOI221_X1 U6017 ( .B1(net226861), .B2(n17745), .C1(\registers[29][1] ), .C2(
        n17742), .A(n12235), .ZN(n12230) );
  OAI22_X1 U6018 ( .A1(n17739), .A2(n15737), .B1(n17736), .B2(n14773), .ZN(
        n12235) );
  AOI221_X1 U6019 ( .B1(\registers[41][1] ), .B2(n17649), .C1(
        \registers[40][1] ), .C2(n17646), .A(n12251), .ZN(n12246) );
  OAI22_X1 U6020 ( .A1(n17643), .A2(n15467), .B1(n17640), .B2(n14774), .ZN(
        n12251) );
  AOI221_X1 U6021 ( .B1(\registers[18][1] ), .B2(n17793), .C1(
        \registers[19][1] ), .C2(n17790), .A(n12227), .ZN(n12222) );
  OAI22_X1 U6022 ( .A1(n17787), .A2(n14606), .B1(n17784), .B2(n15293), .ZN(
        n12227) );
  AOI221_X1 U6023 ( .B1(net226889), .B2(n17745), .C1(\registers[29][2] ), .C2(
        n17742), .A(n12080), .ZN(n12075) );
  OAI22_X1 U6024 ( .A1(n17739), .A2(n15738), .B1(n17736), .B2(n14775), .ZN(
        n12080) );
  AOI221_X1 U6025 ( .B1(\registers[41][2] ), .B2(n17649), .C1(
        \registers[40][2] ), .C2(n17646), .A(n12096), .ZN(n12091) );
  OAI22_X1 U6026 ( .A1(n17643), .A2(n15468), .B1(n17640), .B2(n14776), .ZN(
        n12096) );
  AOI221_X1 U6027 ( .B1(\registers[18][2] ), .B2(n17793), .C1(
        \registers[19][2] ), .C2(n17790), .A(n12072), .ZN(n12067) );
  OAI22_X1 U6028 ( .A1(n17787), .A2(n14607), .B1(n17784), .B2(n15294), .ZN(
        n12072) );
  AOI221_X1 U6029 ( .B1(net226909), .B2(n17745), .C1(\registers[29][3] ), .C2(
        n17742), .A(n11927), .ZN(n11922) );
  OAI22_X1 U6030 ( .A1(n17739), .A2(n15367), .B1(n17736), .B2(n14777), .ZN(
        n11927) );
  AOI221_X1 U6031 ( .B1(\registers[41][3] ), .B2(n17649), .C1(
        \registers[40][3] ), .C2(n17646), .A(n11943), .ZN(n11938) );
  OAI22_X1 U6032 ( .A1(n17643), .A2(n15356), .B1(n17640), .B2(n14641), .ZN(
        n11943) );
  AOI221_X1 U6033 ( .B1(\registers[18][3] ), .B2(n17793), .C1(
        \registers[19][3] ), .C2(n17790), .A(n11919), .ZN(n11914) );
  OAI22_X1 U6034 ( .A1(n17787), .A2(n14608), .B1(n17784), .B2(n15284), .ZN(
        n11919) );
  AOI221_X1 U6035 ( .B1(net226983), .B2(n17745), .C1(\registers[29][4] ), .C2(
        n17742), .A(n10484), .ZN(n10479) );
  OAI22_X1 U6036 ( .A1(n17739), .A2(n15368), .B1(n17736), .B2(n14778), .ZN(
        n10484) );
  AOI221_X1 U6037 ( .B1(\registers[41][4] ), .B2(n17649), .C1(
        \registers[40][4] ), .C2(n17646), .A(n10500), .ZN(n10495) );
  OAI22_X1 U6038 ( .A1(n17643), .A2(n15469), .B1(n17640), .B2(n14779), .ZN(
        n10500) );
  AOI221_X1 U6039 ( .B1(\registers[18][4] ), .B2(n17793), .C1(
        \registers[19][4] ), .C2(n17790), .A(n10476), .ZN(n10471) );
  OAI22_X1 U6040 ( .A1(n17787), .A2(n14569), .B1(n17784), .B2(n15295), .ZN(
        n10476) );
  AOI221_X1 U6041 ( .B1(net226992), .B2(n17745), .C1(\registers[29][5] ), .C2(
        n17742), .A(n10374), .ZN(n10369) );
  OAI22_X1 U6042 ( .A1(n17739), .A2(n15739), .B1(n17736), .B2(n14780), .ZN(
        n10374) );
  AOI221_X1 U6043 ( .B1(\registers[41][5] ), .B2(n17649), .C1(
        \registers[40][5] ), .C2(n17646), .A(n10390), .ZN(n10385) );
  OAI22_X1 U6044 ( .A1(n17643), .A2(n15357), .B1(n17640), .B2(n14642), .ZN(
        n10390) );
  AOI221_X1 U6045 ( .B1(\registers[18][5] ), .B2(n17793), .C1(
        \registers[19][5] ), .C2(n17790), .A(n10366), .ZN(n10361) );
  OAI22_X1 U6046 ( .A1(n17787), .A2(n14609), .B1(n17784), .B2(n15296), .ZN(
        n10366) );
  AOI221_X1 U6047 ( .B1(net227016), .B2(n17745), .C1(\registers[29][6] ), .C2(
        n17742), .A(n10262), .ZN(n10257) );
  OAI22_X1 U6048 ( .A1(n17739), .A2(n15740), .B1(n17736), .B2(n14781), .ZN(
        n10262) );
  AOI221_X1 U6049 ( .B1(\registers[41][6] ), .B2(n17649), .C1(
        \registers[40][6] ), .C2(n17646), .A(n10278), .ZN(n10273) );
  OAI22_X1 U6050 ( .A1(n17643), .A2(n15470), .B1(n17640), .B2(n14782), .ZN(
        n10278) );
  AOI221_X1 U6051 ( .B1(\registers[18][6] ), .B2(n17793), .C1(
        \registers[19][6] ), .C2(n17790), .A(n10254), .ZN(n10249) );
  OAI22_X1 U6052 ( .A1(n17787), .A2(n14610), .B1(n17784), .B2(n15297), .ZN(
        n10254) );
  AOI221_X1 U6053 ( .B1(net227034), .B2(n17745), .C1(\registers[29][7] ), .C2(
        n17742), .A(n7626), .ZN(n7621) );
  OAI22_X1 U6054 ( .A1(n17739), .A2(n15741), .B1(n17736), .B2(n14783), .ZN(
        n7626) );
  AOI221_X1 U6055 ( .B1(\registers[41][7] ), .B2(n17649), .C1(
        \registers[40][7] ), .C2(n17646), .A(n7642), .ZN(n7637) );
  OAI22_X1 U6056 ( .A1(n17643), .A2(n15471), .B1(n17640), .B2(n14784), .ZN(
        n7642) );
  AOI221_X1 U6057 ( .B1(\registers[18][7] ), .B2(n17793), .C1(
        \registers[19][7] ), .C2(n17790), .A(n7618), .ZN(n7613) );
  OAI22_X1 U6058 ( .A1(n17787), .A2(n14611), .B1(n17784), .B2(n15298), .ZN(
        n7618) );
  AOI221_X1 U6059 ( .B1(net227052), .B2(n17745), .C1(\registers[29][8] ), .C2(
        n17742), .A(n7511), .ZN(n7506) );
  OAI22_X1 U6060 ( .A1(n17739), .A2(n15742), .B1(n17736), .B2(n14785), .ZN(
        n7511) );
  AOI221_X1 U6061 ( .B1(\registers[41][8] ), .B2(n17649), .C1(
        \registers[40][8] ), .C2(n17646), .A(n7527), .ZN(n7522) );
  OAI22_X1 U6062 ( .A1(n17643), .A2(n15472), .B1(n17640), .B2(n14786), .ZN(
        n7527) );
  AOI221_X1 U6063 ( .B1(\registers[18][8] ), .B2(n17793), .C1(
        \registers[19][8] ), .C2(n17790), .A(n7503), .ZN(n7498) );
  OAI22_X1 U6064 ( .A1(n17787), .A2(n14612), .B1(n17784), .B2(n15299), .ZN(
        n7503) );
  AOI221_X1 U6065 ( .B1(net227070), .B2(n17745), .C1(\registers[29][9] ), .C2(
        n17742), .A(n7402), .ZN(n7397) );
  OAI22_X1 U6066 ( .A1(n17739), .A2(n15743), .B1(n17736), .B2(n14787), .ZN(
        n7402) );
  AOI221_X1 U6067 ( .B1(\registers[41][9] ), .B2(n17649), .C1(
        \registers[40][9] ), .C2(n17646), .A(n7418), .ZN(n7413) );
  OAI22_X1 U6068 ( .A1(n17643), .A2(n15473), .B1(n17640), .B2(n14788), .ZN(
        n7418) );
  AOI221_X1 U6069 ( .B1(\registers[18][9] ), .B2(n17793), .C1(
        \registers[19][9] ), .C2(n17790), .A(n7394), .ZN(n7389) );
  OAI22_X1 U6070 ( .A1(n17787), .A2(n14613), .B1(n17784), .B2(n15300), .ZN(
        n7394) );
  AOI221_X1 U6071 ( .B1(net227088), .B2(n17745), .C1(\registers[29][10] ), 
        .C2(n17742), .A(n7293), .ZN(n7288) );
  OAI22_X1 U6072 ( .A1(n17739), .A2(n15744), .B1(n17736), .B2(n14789), .ZN(
        n7293) );
  AOI221_X1 U6073 ( .B1(\registers[41][10] ), .B2(n17649), .C1(
        \registers[40][10] ), .C2(n17646), .A(n7309), .ZN(n7304) );
  OAI22_X1 U6074 ( .A1(n17643), .A2(n15474), .B1(n17640), .B2(n14790), .ZN(
        n7309) );
  AOI221_X1 U6075 ( .B1(\registers[18][10] ), .B2(n17793), .C1(
        \registers[19][10] ), .C2(n17790), .A(n7285), .ZN(n7280) );
  OAI22_X1 U6076 ( .A1(n17787), .A2(n14614), .B1(n17784), .B2(n15301), .ZN(
        n7285) );
  AOI221_X1 U6077 ( .B1(net227106), .B2(n17746), .C1(\registers[29][11] ), 
        .C2(n17743), .A(n7179), .ZN(n7174) );
  OAI22_X1 U6078 ( .A1(n17740), .A2(n15745), .B1(n17737), .B2(n14791), .ZN(
        n7179) );
  AOI221_X1 U6079 ( .B1(\registers[41][11] ), .B2(n17650), .C1(
        \registers[40][11] ), .C2(n17647), .A(n7195), .ZN(n7190) );
  OAI22_X1 U6080 ( .A1(n17644), .A2(n15475), .B1(n17641), .B2(n14792), .ZN(
        n7195) );
  AOI221_X1 U6081 ( .B1(\registers[18][11] ), .B2(n17794), .C1(
        \registers[19][11] ), .C2(n17791), .A(n7171), .ZN(n7166) );
  OAI22_X1 U6082 ( .A1(n17788), .A2(n14615), .B1(n17785), .B2(n15302), .ZN(
        n7171) );
  AOI221_X1 U6083 ( .B1(net227124), .B2(n17746), .C1(\registers[29][12] ), 
        .C2(n17743), .A(n7070), .ZN(n7065) );
  OAI22_X1 U6084 ( .A1(n17740), .A2(n15746), .B1(n17737), .B2(n14793), .ZN(
        n7070) );
  AOI221_X1 U6085 ( .B1(\registers[41][12] ), .B2(n17650), .C1(
        \registers[40][12] ), .C2(n17647), .A(n7086), .ZN(n7081) );
  OAI22_X1 U6086 ( .A1(n17644), .A2(n15476), .B1(n17641), .B2(n14794), .ZN(
        n7086) );
  AOI221_X1 U6087 ( .B1(\registers[18][12] ), .B2(n17794), .C1(
        \registers[19][12] ), .C2(n17791), .A(n7062), .ZN(n7057) );
  OAI22_X1 U6088 ( .A1(n17788), .A2(n14616), .B1(n17785), .B2(n15303), .ZN(
        n7062) );
  AOI221_X1 U6089 ( .B1(net227142), .B2(n17746), .C1(\registers[29][13] ), 
        .C2(n17743), .A(n6961), .ZN(n6956) );
  OAI22_X1 U6090 ( .A1(n17740), .A2(n15747), .B1(n17737), .B2(n14795), .ZN(
        n6961) );
  AOI221_X1 U6091 ( .B1(\registers[41][13] ), .B2(n17650), .C1(
        \registers[40][13] ), .C2(n17647), .A(n6977), .ZN(n6972) );
  OAI22_X1 U6092 ( .A1(n17644), .A2(n15477), .B1(n17641), .B2(n14796), .ZN(
        n6977) );
  AOI221_X1 U6093 ( .B1(\registers[18][13] ), .B2(n17794), .C1(
        \registers[19][13] ), .C2(n17791), .A(n6953), .ZN(n6948) );
  OAI22_X1 U6094 ( .A1(n17788), .A2(n14617), .B1(n17785), .B2(n15304), .ZN(
        n6953) );
  AOI221_X1 U6095 ( .B1(net227160), .B2(n17746), .C1(\registers[29][14] ), 
        .C2(n17743), .A(n6852), .ZN(n6847) );
  OAI22_X1 U6096 ( .A1(n17740), .A2(n15748), .B1(n17737), .B2(n14797), .ZN(
        n6852) );
  AOI221_X1 U6097 ( .B1(\registers[41][14] ), .B2(n17650), .C1(
        \registers[40][14] ), .C2(n17647), .A(n6868), .ZN(n6863) );
  OAI22_X1 U6098 ( .A1(n17644), .A2(n15478), .B1(n17641), .B2(n14798), .ZN(
        n6868) );
  AOI221_X1 U6099 ( .B1(\registers[18][14] ), .B2(n17794), .C1(
        \registers[19][14] ), .C2(n17791), .A(n6844), .ZN(n6839) );
  OAI22_X1 U6100 ( .A1(n17788), .A2(n14618), .B1(n17785), .B2(n15305), .ZN(
        n6844) );
  AOI221_X1 U6101 ( .B1(net227178), .B2(n17746), .C1(\registers[29][15] ), 
        .C2(n17743), .A(n6743), .ZN(n6738) );
  OAI22_X1 U6102 ( .A1(n17740), .A2(n15749), .B1(n17737), .B2(n14799), .ZN(
        n6743) );
  AOI221_X1 U6103 ( .B1(\registers[41][15] ), .B2(n17650), .C1(
        \registers[40][15] ), .C2(n17647), .A(n6759), .ZN(n6754) );
  OAI22_X1 U6104 ( .A1(n17644), .A2(n15479), .B1(n17641), .B2(n14800), .ZN(
        n6759) );
  AOI221_X1 U6105 ( .B1(\registers[18][15] ), .B2(n17794), .C1(
        \registers[19][15] ), .C2(n17791), .A(n6735), .ZN(n6730) );
  OAI22_X1 U6106 ( .A1(n17788), .A2(n14619), .B1(n17785), .B2(n15306), .ZN(
        n6735) );
  AOI221_X1 U6107 ( .B1(net227196), .B2(n17746), .C1(\registers[29][16] ), 
        .C2(n17743), .A(n6600), .ZN(n6580) );
  OAI22_X1 U6108 ( .A1(n17740), .A2(n15750), .B1(n17737), .B2(n14801), .ZN(
        n6600) );
  AOI221_X1 U6109 ( .B1(\registers[41][16] ), .B2(n17650), .C1(
        \registers[40][16] ), .C2(n17647), .A(n6619), .ZN(n6614) );
  OAI22_X1 U6110 ( .A1(n17644), .A2(n15480), .B1(n17641), .B2(n14802), .ZN(
        n6619) );
  AOI221_X1 U6111 ( .B1(\registers[18][16] ), .B2(n17794), .C1(
        \registers[19][16] ), .C2(n17791), .A(n6575), .ZN(n6568) );
  OAI22_X1 U6112 ( .A1(n17788), .A2(n14620), .B1(n17785), .B2(n15307), .ZN(
        n6575) );
  AOI221_X1 U6113 ( .B1(net227214), .B2(n17746), .C1(\registers[29][17] ), 
        .C2(n17743), .A(n6413), .ZN(n6393) );
  OAI22_X1 U6114 ( .A1(n17740), .A2(n15751), .B1(n17737), .B2(n14803), .ZN(
        n6413) );
  AOI221_X1 U6115 ( .B1(\registers[41][17] ), .B2(n17650), .C1(
        \registers[40][17] ), .C2(n17647), .A(n6434), .ZN(n6427) );
  OAI22_X1 U6116 ( .A1(n17644), .A2(n15481), .B1(n17641), .B2(n14804), .ZN(
        n6434) );
  AOI221_X1 U6117 ( .B1(\registers[18][17] ), .B2(n17794), .C1(
        \registers[19][17] ), .C2(n17791), .A(n6388), .ZN(n6383) );
  OAI22_X1 U6118 ( .A1(n17788), .A2(n14621), .B1(n17785), .B2(n15308), .ZN(
        n6388) );
  AOI221_X1 U6119 ( .B1(net227232), .B2(n17746), .C1(\registers[29][18] ), 
        .C2(n17743), .A(n6226), .ZN(n6221) );
  OAI22_X1 U6120 ( .A1(n17740), .A2(n15752), .B1(n17737), .B2(n14805), .ZN(
        n6226) );
  AOI221_X1 U6121 ( .B1(\registers[41][18] ), .B2(n17650), .C1(
        \registers[40][18] ), .C2(n17647), .A(n6248), .ZN(n6240) );
  OAI22_X1 U6122 ( .A1(n17644), .A2(n15482), .B1(n17641), .B2(n14806), .ZN(
        n6248) );
  AOI221_X1 U6123 ( .B1(\registers[18][18] ), .B2(n17794), .C1(
        \registers[19][18] ), .C2(n17791), .A(n6203), .ZN(n6196) );
  OAI22_X1 U6124 ( .A1(n17788), .A2(n14622), .B1(n17785), .B2(n15309), .ZN(
        n6203) );
  AOI221_X1 U6125 ( .B1(net227250), .B2(n17746), .C1(\registers[29][19] ), 
        .C2(n17743), .A(n6039), .ZN(n6034) );
  OAI22_X1 U6126 ( .A1(n17740), .A2(n15753), .B1(n17737), .B2(n14807), .ZN(
        n6039) );
  AOI221_X1 U6127 ( .B1(\registers[41][19] ), .B2(n17650), .C1(
        \registers[40][19] ), .C2(n17647), .A(n6061), .ZN(n6055) );
  OAI22_X1 U6128 ( .A1(n17644), .A2(n15483), .B1(n17641), .B2(n14808), .ZN(
        n6061) );
  AOI221_X1 U6129 ( .B1(\registers[18][19] ), .B2(n17794), .C1(
        \registers[19][19] ), .C2(n17791), .A(n6031), .ZN(n6009) );
  OAI22_X1 U6130 ( .A1(n17788), .A2(n14623), .B1(n17785), .B2(n15310), .ZN(
        n6031) );
  AOI221_X1 U6131 ( .B1(net227268), .B2(n17746), .C1(\registers[29][20] ), 
        .C2(n17743), .A(n5853), .ZN(n5847) );
  OAI22_X1 U6132 ( .A1(n17740), .A2(n15754), .B1(n17737), .B2(n14809), .ZN(
        n5853) );
  AOI221_X1 U6133 ( .B1(\registers[41][20] ), .B2(n17650), .C1(
        \registers[40][20] ), .C2(n17647), .A(n5875), .ZN(n5869) );
  OAI22_X1 U6134 ( .A1(n17644), .A2(n15484), .B1(n17641), .B2(n14810), .ZN(
        n5875) );
  AOI221_X1 U6135 ( .B1(\registers[18][20] ), .B2(n17794), .C1(
        \registers[19][20] ), .C2(n17791), .A(n5844), .ZN(n5824) );
  OAI22_X1 U6136 ( .A1(n17788), .A2(n14624), .B1(n17785), .B2(n15311), .ZN(
        n5844) );
  AOI221_X1 U6137 ( .B1(net227286), .B2(n17746), .C1(\registers[29][21] ), 
        .C2(n17743), .A(n5667), .ZN(n5660) );
  OAI22_X1 U6138 ( .A1(n17740), .A2(n15755), .B1(n17737), .B2(n14811), .ZN(
        n5667) );
  AOI221_X1 U6139 ( .B1(\registers[41][21] ), .B2(n17650), .C1(
        \registers[40][21] ), .C2(n17647), .A(n5690), .ZN(n5682) );
  OAI22_X1 U6140 ( .A1(n17644), .A2(n15485), .B1(n17641), .B2(n14812), .ZN(
        n5690) );
  AOI221_X1 U6141 ( .B1(\registers[18][21] ), .B2(n17794), .C1(
        \registers[19][21] ), .C2(n17791), .A(n5657), .ZN(n5637) );
  OAI22_X1 U6142 ( .A1(n17788), .A2(n14625), .B1(n17785), .B2(n15312), .ZN(
        n5657) );
  AOI221_X1 U6143 ( .B1(net227304), .B2(n17746), .C1(\registers[29][22] ), 
        .C2(n17743), .A(n5481), .ZN(n5473) );
  OAI22_X1 U6144 ( .A1(n17740), .A2(n15756), .B1(n17737), .B2(n14813), .ZN(
        n5481) );
  AOI221_X1 U6145 ( .B1(\registers[41][22] ), .B2(n17650), .C1(
        \registers[40][22] ), .C2(n17647), .A(n5503), .ZN(n5495) );
  OAI22_X1 U6146 ( .A1(n17644), .A2(n15486), .B1(n17641), .B2(n14814), .ZN(
        n5503) );
  AOI221_X1 U6147 ( .B1(\registers[18][22] ), .B2(n17794), .C1(
        \registers[19][22] ), .C2(n17791), .A(n5470), .ZN(n5465) );
  OAI22_X1 U6148 ( .A1(n17788), .A2(n14626), .B1(n17785), .B2(n15313), .ZN(
        n5470) );
  AOI221_X1 U6149 ( .B1(net227466), .B2(n17745), .C1(\registers[29][31] ), 
        .C2(n17742), .A(n14139), .ZN(n14110) );
  OAI22_X1 U6150 ( .A1(n17739), .A2(n15757), .B1(n17736), .B2(n14815), .ZN(
        n14139) );
  AOI221_X1 U6151 ( .B1(\registers[41][31] ), .B2(n17649), .C1(
        \registers[40][31] ), .C2(n17646), .A(n14203), .ZN(n14188) );
  OAI22_X1 U6152 ( .A1(n17643), .A2(n15487), .B1(n17640), .B2(n14816), .ZN(
        n14203) );
  AOI221_X1 U6153 ( .B1(\registers[18][31] ), .B2(n17793), .C1(
        \registers[19][31] ), .C2(n17790), .A(n14102), .ZN(n14081) );
  OAI22_X1 U6154 ( .A1(n17787), .A2(n14627), .B1(n17784), .B2(n15314), .ZN(
        n14102) );
  AOI221_X1 U6155 ( .B1(\registers[50][24] ), .B2(n16279), .C1(net227335), 
        .C2(n16276), .A(n12922), .ZN(n12915) );
  OAI22_X1 U6156 ( .A1(n16273), .A2(n12349), .B1(n16270), .B2(n14931), .ZN(
        n12922) );
  AOI221_X1 U6157 ( .B1(\registers[50][25] ), .B2(n16279), .C1(net227353), 
        .C2(n16276), .A(n12880), .ZN(n12873) );
  OAI22_X1 U6158 ( .A1(n16273), .A2(n12350), .B1(n16270), .B2(n14932), .ZN(
        n12880) );
  AOI221_X1 U6159 ( .B1(\registers[50][26] ), .B2(n16279), .C1(net227371), 
        .C2(n16276), .A(n12838), .ZN(n12831) );
  OAI22_X1 U6160 ( .A1(n16273), .A2(n12351), .B1(n16270), .B2(n14933), .ZN(
        n12838) );
  AOI221_X1 U6161 ( .B1(\registers[50][27] ), .B2(n16279), .C1(net227389), 
        .C2(n16276), .A(n12796), .ZN(n12789) );
  OAI22_X1 U6162 ( .A1(n16273), .A2(n12352), .B1(n16270), .B2(n14934), .ZN(
        n12796) );
  AOI221_X1 U6163 ( .B1(\registers[50][28] ), .B2(n16279), .C1(net227407), 
        .C2(n16276), .A(n12754), .ZN(n12747) );
  OAI22_X1 U6164 ( .A1(n16273), .A2(n12353), .B1(n16270), .B2(n14935), .ZN(
        n12754) );
  AOI221_X1 U6165 ( .B1(\registers[50][29] ), .B2(n16279), .C1(net227425), 
        .C2(n16276), .A(n12712), .ZN(n12705) );
  OAI22_X1 U6166 ( .A1(n16273), .A2(n12354), .B1(n16270), .B2(n14936), .ZN(
        n12712) );
  AOI221_X1 U6167 ( .B1(\registers[50][30] ), .B2(n16279), .C1(net227443), 
        .C2(n16276), .A(n12670), .ZN(n12662) );
  OAI22_X1 U6168 ( .A1(n16273), .A2(n12197), .B1(n16270), .B2(n14855), .ZN(
        n12670) );
  AOI221_X1 U6169 ( .B1(\registers[50][31] ), .B2(n16279), .C1(net227461), 
        .C2(n16276), .A(n12605), .ZN(n12582) );
  OAI22_X1 U6170 ( .A1(n16273), .A2(n12355), .B1(n16270), .B2(n14937), .ZN(
        n12605) );
  AOI221_X1 U6171 ( .B1(\registers[50][24] ), .B2(n16531), .C1(net227335), 
        .C2(n16528), .A(n10972), .ZN(n10965) );
  OAI22_X1 U6172 ( .A1(n16525), .A2(n12349), .B1(n16522), .B2(n14931), .ZN(
        n10972) );
  AOI221_X1 U6173 ( .B1(\registers[7][24] ), .B2(n16480), .C1(
        \registers[42][24] ), .C2(n16477), .A(n10980), .ZN(n10973) );
  OAI22_X1 U6174 ( .A1(n16474), .A2(n15233), .B1(n16471), .B2(n14352), .ZN(
        n10980) );
  AOI221_X1 U6175 ( .B1(\registers[50][25] ), .B2(n16531), .C1(net227353), 
        .C2(n16528), .A(n10929), .ZN(n10922) );
  OAI22_X1 U6176 ( .A1(n16525), .A2(n12350), .B1(n16522), .B2(n14932), .ZN(
        n10929) );
  AOI221_X1 U6177 ( .B1(\registers[7][25] ), .B2(n16480), .C1(
        \registers[42][25] ), .C2(n16477), .A(n10937), .ZN(n10930) );
  OAI22_X1 U6178 ( .A1(n16474), .A2(n15234), .B1(n16471), .B2(n14353), .ZN(
        n10937) );
  AOI221_X1 U6179 ( .B1(\registers[50][26] ), .B2(n16531), .C1(net227371), 
        .C2(n16528), .A(n10886), .ZN(n10879) );
  OAI22_X1 U6180 ( .A1(n16525), .A2(n12351), .B1(n16522), .B2(n14933), .ZN(
        n10886) );
  AOI221_X1 U6181 ( .B1(\registers[7][26] ), .B2(n16480), .C1(
        \registers[42][26] ), .C2(n16477), .A(n10894), .ZN(n10887) );
  OAI22_X1 U6182 ( .A1(n16474), .A2(n15235), .B1(n16471), .B2(n14354), .ZN(
        n10894) );
  AOI221_X1 U6183 ( .B1(\registers[50][27] ), .B2(n16531), .C1(net227389), 
        .C2(n16528), .A(n10843), .ZN(n10836) );
  OAI22_X1 U6184 ( .A1(n16525), .A2(n12352), .B1(n16522), .B2(n14934), .ZN(
        n10843) );
  AOI221_X1 U6185 ( .B1(\registers[7][27] ), .B2(n16480), .C1(
        \registers[42][27] ), .C2(n16477), .A(n10851), .ZN(n10844) );
  OAI22_X1 U6186 ( .A1(n16474), .A2(n15236), .B1(n16471), .B2(n14355), .ZN(
        n10851) );
  AOI221_X1 U6187 ( .B1(\registers[50][28] ), .B2(n16531), .C1(net227407), 
        .C2(n16528), .A(n10800), .ZN(n10793) );
  OAI22_X1 U6188 ( .A1(n16525), .A2(n12353), .B1(n16522), .B2(n14935), .ZN(
        n10800) );
  AOI221_X1 U6189 ( .B1(\registers[7][28] ), .B2(n16480), .C1(
        \registers[42][28] ), .C2(n16477), .A(n10808), .ZN(n10801) );
  OAI22_X1 U6190 ( .A1(n16474), .A2(n15237), .B1(n16471), .B2(n14356), .ZN(
        n10808) );
  AOI221_X1 U6191 ( .B1(\registers[50][29] ), .B2(n16531), .C1(net227425), 
        .C2(n16528), .A(n10757), .ZN(n10750) );
  OAI22_X1 U6192 ( .A1(n16525), .A2(n12354), .B1(n16522), .B2(n14936), .ZN(
        n10757) );
  AOI221_X1 U6193 ( .B1(\registers[7][29] ), .B2(n16480), .C1(
        \registers[42][29] ), .C2(n16477), .A(n10765), .ZN(n10758) );
  OAI22_X1 U6194 ( .A1(n16474), .A2(n15238), .B1(n16471), .B2(n14357), .ZN(
        n10765) );
  AOI221_X1 U6195 ( .B1(\registers[50][30] ), .B2(n16531), .C1(net227443), 
        .C2(n16528), .A(n10711), .ZN(n10700) );
  OAI22_X1 U6196 ( .A1(n16525), .A2(n12197), .B1(n16522), .B2(n14855), .ZN(
        n10711) );
  AOI221_X1 U6197 ( .B1(\registers[7][30] ), .B2(n16480), .C1(
        \registers[42][30] ), .C2(n16477), .A(n10720), .ZN(n10713) );
  OAI22_X1 U6198 ( .A1(n16474), .A2(n14874), .B1(n16471), .B2(n14055), .ZN(
        n10720) );
  AOI221_X1 U6199 ( .B1(\registers[50][31] ), .B2(n16531), .C1(net227461), 
        .C2(n16528), .A(n10623), .ZN(n10596) );
  OAI22_X1 U6200 ( .A1(n16525), .A2(n12355), .B1(n16522), .B2(n14937), .ZN(
        n10623) );
  AOI221_X1 U6201 ( .B1(\registers[7][31] ), .B2(n16480), .C1(
        \registers[42][31] ), .C2(n16477), .A(n10657), .ZN(n10628) );
  OAI22_X1 U6202 ( .A1(n16474), .A2(n15239), .B1(n16471), .B2(n14358), .ZN(
        n10657) );
  AOI221_X1 U6203 ( .B1(\registers[48][23] ), .B2(n17639), .C1(
        \registers[4][23] ), .C2(n17636), .A(n5319), .ZN(n5309) );
  OAI22_X1 U6204 ( .A1(n17633), .A2(n15488), .B1(n17630), .B2(n14671), .ZN(
        n5319) );
  AOI221_X1 U6205 ( .B1(\registers[23][23] ), .B2(n17783), .C1(
        \registers[22][23] ), .C2(n17780), .A(n5285), .ZN(n5277) );
  OAI22_X1 U6206 ( .A1(n17777), .A2(n12198), .B1(n17774), .B2(n14824), .ZN(
        n5285) );
  AOI221_X1 U6207 ( .B1(\registers[48][24] ), .B2(n17639), .C1(
        \registers[4][24] ), .C2(n17636), .A(n5147), .ZN(n5138) );
  OAI22_X1 U6208 ( .A1(n17633), .A2(n15489), .B1(n17630), .B2(n14672), .ZN(
        n5147) );
  AOI221_X1 U6209 ( .B1(\registers[23][24] ), .B2(n17783), .C1(
        \registers[22][24] ), .C2(n17780), .A(n5119), .ZN(n5111) );
  OAI22_X1 U6210 ( .A1(n17777), .A2(n12199), .B1(n17774), .B2(n14825), .ZN(
        n5119) );
  AOI221_X1 U6211 ( .B1(\registers[48][25] ), .B2(n17639), .C1(
        \registers[4][25] ), .C2(n17636), .A(n5031), .ZN(n5024) );
  OAI22_X1 U6212 ( .A1(n17633), .A2(n15490), .B1(n17630), .B2(n14673), .ZN(
        n5031) );
  AOI221_X1 U6213 ( .B1(\registers[23][25] ), .B2(n17783), .C1(
        \registers[22][25] ), .C2(n17780), .A(n5005), .ZN(n4998) );
  OAI22_X1 U6214 ( .A1(n17777), .A2(n12200), .B1(n17774), .B2(n14826), .ZN(
        n5005) );
  AOI221_X1 U6215 ( .B1(\registers[48][26] ), .B2(n17639), .C1(
        \registers[4][26] ), .C2(n17636), .A(n4913), .ZN(n4906) );
  OAI22_X1 U6216 ( .A1(n17633), .A2(n15491), .B1(n17630), .B2(n14674), .ZN(
        n4913) );
  AOI221_X1 U6217 ( .B1(\registers[23][26] ), .B2(n17783), .C1(
        \registers[22][26] ), .C2(n17780), .A(n4883), .ZN(n4876) );
  OAI22_X1 U6218 ( .A1(n17777), .A2(n12201), .B1(n17774), .B2(n14827), .ZN(
        n4883) );
  AOI221_X1 U6219 ( .B1(\registers[48][27] ), .B2(n17639), .C1(
        \registers[4][27] ), .C2(n17636), .A(n4782), .ZN(n4775) );
  OAI22_X1 U6220 ( .A1(n17633), .A2(n15492), .B1(n17630), .B2(n14675), .ZN(
        n4782) );
  AOI221_X1 U6221 ( .B1(\registers[23][27] ), .B2(n17783), .C1(
        \registers[22][27] ), .C2(n17780), .A(n4756), .ZN(n4745) );
  OAI22_X1 U6222 ( .A1(n17777), .A2(n12202), .B1(n17774), .B2(n14828), .ZN(
        n4756) );
  AOI221_X1 U6223 ( .B1(\registers[48][28] ), .B2(n17639), .C1(
        \registers[4][28] ), .C2(n17636), .A(n4653), .ZN(n4642) );
  OAI22_X1 U6224 ( .A1(n17633), .A2(n15493), .B1(n17630), .B2(n14676), .ZN(
        n4653) );
  AOI221_X1 U6225 ( .B1(\registers[23][28] ), .B2(n17783), .C1(
        \registers[22][28] ), .C2(n17780), .A(n4625), .ZN(n4618) );
  OAI22_X1 U6226 ( .A1(n17777), .A2(n12203), .B1(n17774), .B2(n14829), .ZN(
        n4625) );
  AOI221_X1 U6227 ( .B1(\registers[48][29] ), .B2(n17639), .C1(
        \registers[4][29] ), .C2(n17636), .A(n4524), .ZN(n4517) );
  OAI22_X1 U6228 ( .A1(n17633), .A2(n15494), .B1(n17630), .B2(n14677), .ZN(
        n4524) );
  AOI221_X1 U6229 ( .B1(\registers[23][29] ), .B2(n17783), .C1(
        \registers[22][29] ), .C2(n17780), .A(n4492), .ZN(n4485) );
  OAI22_X1 U6230 ( .A1(n17777), .A2(n12204), .B1(n17774), .B2(n14830), .ZN(
        n4492) );
  AOI221_X1 U6231 ( .B1(\registers[48][30] ), .B2(n17639), .C1(
        \registers[4][30] ), .C2(n17636), .A(n4241), .ZN(n4213) );
  OAI22_X1 U6232 ( .A1(n17633), .A2(n15276), .B1(n17630), .B2(n14628), .ZN(
        n4241) );
  AOI221_X1 U6233 ( .B1(\registers[23][30] ), .B2(n17783), .C1(
        \registers[22][30] ), .C2(n17780), .A(n4132), .ZN(n4101) );
  OAI22_X1 U6234 ( .A1(n17777), .A2(n12161), .B1(n17774), .B2(n14822), .ZN(
        n4132) );
  AOI221_X1 U6235 ( .B1(\registers[7][0] ), .B2(n16226), .C1(
        \registers[42][0] ), .C2(n16223), .A(n13977), .ZN(n13964) );
  OAI22_X1 U6236 ( .A1(n16220), .A2(n15210), .B1(n16217), .B2(n14329), .ZN(
        n13977) );
  AOI221_X1 U6237 ( .B1(\registers[7][1] ), .B2(n16226), .C1(
        \registers[42][1] ), .C2(n16223), .A(n13896), .ZN(n13889) );
  OAI22_X1 U6238 ( .A1(n16220), .A2(n15211), .B1(n16217), .B2(n14330), .ZN(
        n13896) );
  AOI221_X1 U6239 ( .B1(\registers[7][2] ), .B2(n16226), .C1(
        \registers[42][2] ), .C2(n16223), .A(n13854), .ZN(n13847) );
  OAI22_X1 U6240 ( .A1(n16220), .A2(n15212), .B1(n16217), .B2(n14331), .ZN(
        n13854) );
  AOI221_X1 U6241 ( .B1(\registers[7][3] ), .B2(n16226), .C1(
        \registers[42][3] ), .C2(n16223), .A(n13812), .ZN(n13805) );
  OAI22_X1 U6242 ( .A1(n16220), .A2(n15003), .B1(n16217), .B2(n14288), .ZN(
        n13812) );
  AOI221_X1 U6243 ( .B1(\registers[7][4] ), .B2(n16226), .C1(
        \registers[42][4] ), .C2(n16223), .A(n13770), .ZN(n13763) );
  OAI22_X1 U6244 ( .A1(n16220), .A2(n15213), .B1(n16217), .B2(n14332), .ZN(
        n13770) );
  AOI221_X1 U6245 ( .B1(\registers[7][5] ), .B2(n16226), .C1(
        \registers[42][5] ), .C2(n16223), .A(n13728), .ZN(n13721) );
  OAI22_X1 U6246 ( .A1(n16220), .A2(n15214), .B1(n16217), .B2(n14333), .ZN(
        n13728) );
  AOI221_X1 U6247 ( .B1(\registers[7][6] ), .B2(n16226), .C1(
        \registers[42][6] ), .C2(n16223), .A(n13686), .ZN(n13679) );
  OAI22_X1 U6248 ( .A1(n16220), .A2(n15215), .B1(n16217), .B2(n14334), .ZN(
        n13686) );
  AOI221_X1 U6249 ( .B1(\registers[7][7] ), .B2(n16226), .C1(
        \registers[42][7] ), .C2(n16223), .A(n13644), .ZN(n13637) );
  OAI22_X1 U6250 ( .A1(n16220), .A2(n15216), .B1(n16217), .B2(n14335), .ZN(
        n13644) );
  AOI221_X1 U6251 ( .B1(\registers[7][8] ), .B2(n16226), .C1(
        \registers[42][8] ), .C2(n16223), .A(n13602), .ZN(n13595) );
  OAI22_X1 U6252 ( .A1(n16220), .A2(n15217), .B1(n16217), .B2(n14336), .ZN(
        n13602) );
  AOI221_X1 U6253 ( .B1(\registers[7][9] ), .B2(n16226), .C1(
        \registers[42][9] ), .C2(n16223), .A(n13560), .ZN(n13553) );
  OAI22_X1 U6254 ( .A1(n16220), .A2(n15218), .B1(n16217), .B2(n14337), .ZN(
        n13560) );
  AOI221_X1 U6255 ( .B1(\registers[7][10] ), .B2(n16226), .C1(
        \registers[42][10] ), .C2(n16223), .A(n13518), .ZN(n13511) );
  OAI22_X1 U6256 ( .A1(n16220), .A2(n15219), .B1(n16217), .B2(n14338), .ZN(
        n13518) );
  AOI221_X1 U6257 ( .B1(\registers[7][11] ), .B2(n16226), .C1(
        \registers[42][11] ), .C2(n16223), .A(n13476), .ZN(n13469) );
  OAI22_X1 U6258 ( .A1(n16220), .A2(n15220), .B1(n16217), .B2(n14339), .ZN(
        n13476) );
  AOI221_X1 U6259 ( .B1(\registers[7][12] ), .B2(n16227), .C1(
        \registers[42][12] ), .C2(n16224), .A(n13434), .ZN(n13427) );
  OAI22_X1 U6260 ( .A1(n16221), .A2(n15221), .B1(n16218), .B2(n14340), .ZN(
        n13434) );
  AOI221_X1 U6261 ( .B1(\registers[7][13] ), .B2(n16227), .C1(
        \registers[42][13] ), .C2(n16224), .A(n13392), .ZN(n13385) );
  OAI22_X1 U6262 ( .A1(n16221), .A2(n15222), .B1(n16218), .B2(n14341), .ZN(
        n13392) );
  AOI221_X1 U6263 ( .B1(\registers[7][14] ), .B2(n16227), .C1(
        \registers[42][14] ), .C2(n16224), .A(n13350), .ZN(n13343) );
  OAI22_X1 U6264 ( .A1(n16221), .A2(n15223), .B1(n16218), .B2(n14342), .ZN(
        n13350) );
  AOI221_X1 U6265 ( .B1(\registers[7][15] ), .B2(n16227), .C1(
        \registers[42][15] ), .C2(n16224), .A(n13308), .ZN(n13301) );
  OAI22_X1 U6266 ( .A1(n16221), .A2(n15224), .B1(n16218), .B2(n14343), .ZN(
        n13308) );
  AOI221_X1 U6267 ( .B1(\registers[7][16] ), .B2(n16227), .C1(
        \registers[42][16] ), .C2(n16224), .A(n13266), .ZN(n13259) );
  OAI22_X1 U6268 ( .A1(n16221), .A2(n15225), .B1(n16218), .B2(n14344), .ZN(
        n13266) );
  AOI221_X1 U6269 ( .B1(\registers[7][17] ), .B2(n16227), .C1(
        \registers[42][17] ), .C2(n16224), .A(n13224), .ZN(n13217) );
  OAI22_X1 U6270 ( .A1(n16221), .A2(n15226), .B1(n16218), .B2(n14345), .ZN(
        n13224) );
  AOI221_X1 U6271 ( .B1(\registers[7][18] ), .B2(n16227), .C1(
        \registers[42][18] ), .C2(n16224), .A(n13182), .ZN(n13175) );
  OAI22_X1 U6272 ( .A1(n16221), .A2(n15227), .B1(n16218), .B2(n14346), .ZN(
        n13182) );
  AOI221_X1 U6273 ( .B1(\registers[7][19] ), .B2(n16227), .C1(
        \registers[42][19] ), .C2(n16224), .A(n13140), .ZN(n13133) );
  OAI22_X1 U6274 ( .A1(n16221), .A2(n15228), .B1(n16218), .B2(n14347), .ZN(
        n13140) );
  AOI221_X1 U6275 ( .B1(\registers[7][20] ), .B2(n16227), .C1(
        \registers[42][20] ), .C2(n16224), .A(n13098), .ZN(n13091) );
  OAI22_X1 U6276 ( .A1(n16221), .A2(n15229), .B1(n16218), .B2(n14348), .ZN(
        n13098) );
  AOI221_X1 U6277 ( .B1(\registers[7][21] ), .B2(n16227), .C1(
        \registers[42][21] ), .C2(n16224), .A(n13056), .ZN(n13049) );
  OAI22_X1 U6278 ( .A1(n16221), .A2(n15230), .B1(n16218), .B2(n14349), .ZN(
        n13056) );
  AOI221_X1 U6279 ( .B1(\registers[7][22] ), .B2(n16227), .C1(
        \registers[42][22] ), .C2(n16224), .A(n13014), .ZN(n13007) );
  OAI22_X1 U6280 ( .A1(n16221), .A2(n15231), .B1(n16218), .B2(n14350), .ZN(
        n13014) );
  AOI221_X1 U6281 ( .B1(\registers[7][23] ), .B2(n16227), .C1(
        \registers[42][23] ), .C2(n16224), .A(n12972), .ZN(n12965) );
  OAI22_X1 U6282 ( .A1(n16221), .A2(n15232), .B1(n16218), .B2(n14351), .ZN(
        n12972) );
  AOI221_X1 U6283 ( .B1(\registers[50][0] ), .B2(n16529), .C1(net226846), .C2(
        n16526), .A(n12478), .ZN(n12467) );
  OAI22_X1 U6284 ( .A1(n16523), .A2(n12356), .B1(n16520), .B2(n14938), .ZN(
        n12478) );
  AOI221_X1 U6285 ( .B1(\registers[7][0] ), .B2(n16478), .C1(
        \registers[42][0] ), .C2(n16475), .A(n12496), .ZN(n12483) );
  OAI22_X1 U6286 ( .A1(n16472), .A2(n15210), .B1(n16469), .B2(n14329), .ZN(
        n12496) );
  AOI221_X1 U6287 ( .B1(\registers[50][1] ), .B2(n16529), .C1(net226859), .C2(
        n16526), .A(n12292), .ZN(n12285) );
  OAI22_X1 U6288 ( .A1(n16523), .A2(n12358), .B1(n16520), .B2(n14939), .ZN(
        n12292) );
  AOI221_X1 U6289 ( .B1(\registers[7][1] ), .B2(n16478), .C1(
        \registers[42][1] ), .C2(n16475), .A(n12300), .ZN(n12293) );
  OAI22_X1 U6290 ( .A1(n16472), .A2(n15211), .B1(n16469), .B2(n14330), .ZN(
        n12300) );
  AOI221_X1 U6291 ( .B1(\registers[50][2] ), .B2(n16529), .C1(net226885), .C2(
        n16526), .A(n12139), .ZN(n12132) );
  OAI22_X1 U6292 ( .A1(n16523), .A2(n12360), .B1(n16520), .B2(n14940), .ZN(
        n12139) );
  AOI221_X1 U6293 ( .B1(\registers[7][2] ), .B2(n16478), .C1(
        \registers[42][2] ), .C2(n16475), .A(n12147), .ZN(n12140) );
  OAI22_X1 U6294 ( .A1(n16472), .A2(n15212), .B1(n16469), .B2(n14331), .ZN(
        n12147) );
  AOI221_X1 U6295 ( .B1(\registers[50][3] ), .B2(n16529), .C1(net226898), .C2(
        n16526), .A(n11986), .ZN(n11979) );
  OAI22_X1 U6296 ( .A1(n16523), .A2(n12340), .B1(n16520), .B2(n14941), .ZN(
        n11986) );
  AOI221_X1 U6297 ( .B1(\registers[7][3] ), .B2(n16478), .C1(
        \registers[42][3] ), .C2(n16475), .A(n11994), .ZN(n11987) );
  OAI22_X1 U6298 ( .A1(n16472), .A2(n15003), .B1(n16469), .B2(n14288), .ZN(
        n11994) );
  AOI221_X1 U6299 ( .B1(\registers[50][4] ), .B2(n16529), .C1(net226980), .C2(
        n16526), .A(n11833), .ZN(n11826) );
  OAI22_X1 U6300 ( .A1(n16523), .A2(n12341), .B1(n16520), .B2(n14866), .ZN(
        n11833) );
  AOI221_X1 U6301 ( .B1(\registers[7][4] ), .B2(n16478), .C1(
        \registers[42][4] ), .C2(n16475), .A(n11841), .ZN(n11834) );
  OAI22_X1 U6302 ( .A1(n16472), .A2(n15213), .B1(n16469), .B2(n14332), .ZN(
        n11841) );
  AOI221_X1 U6303 ( .B1(\registers[50][5] ), .B2(n16529), .C1(net227000), .C2(
        n16526), .A(n11790), .ZN(n11783) );
  OAI22_X1 U6304 ( .A1(n16523), .A2(n12364), .B1(n16520), .B2(n14867), .ZN(
        n11790) );
  AOI221_X1 U6305 ( .B1(\registers[7][5] ), .B2(n16478), .C1(
        \registers[42][5] ), .C2(n16475), .A(n11798), .ZN(n11791) );
  OAI22_X1 U6306 ( .A1(n16472), .A2(n15214), .B1(n16469), .B2(n14333), .ZN(
        n11798) );
  AOI221_X1 U6307 ( .B1(\registers[50][6] ), .B2(n16529), .C1(net227011), .C2(
        n16526), .A(n11747), .ZN(n11740) );
  OAI22_X1 U6308 ( .A1(n16523), .A2(n12366), .B1(n16520), .B2(n14942), .ZN(
        n11747) );
  AOI221_X1 U6309 ( .B1(\registers[7][6] ), .B2(n16478), .C1(
        \registers[42][6] ), .C2(n16475), .A(n11755), .ZN(n11748) );
  OAI22_X1 U6310 ( .A1(n16472), .A2(n15215), .B1(n16469), .B2(n14334), .ZN(
        n11755) );
  AOI221_X1 U6311 ( .B1(\registers[50][7] ), .B2(n16529), .C1(net227029), .C2(
        n16526), .A(n11704), .ZN(n11697) );
  OAI22_X1 U6312 ( .A1(n16523), .A2(n12368), .B1(n16520), .B2(n14943), .ZN(
        n11704) );
  AOI221_X1 U6313 ( .B1(\registers[7][7] ), .B2(n16478), .C1(
        \registers[42][7] ), .C2(n16475), .A(n11712), .ZN(n11705) );
  OAI22_X1 U6314 ( .A1(n16472), .A2(n15216), .B1(n16469), .B2(n14335), .ZN(
        n11712) );
  AOI221_X1 U6315 ( .B1(\registers[50][8] ), .B2(n16529), .C1(net227047), .C2(
        n16526), .A(n11661), .ZN(n11654) );
  OAI22_X1 U6316 ( .A1(n16523), .A2(n12407), .B1(n16520), .B2(n14944), .ZN(
        n11661) );
  AOI221_X1 U6317 ( .B1(\registers[7][8] ), .B2(n16478), .C1(
        \registers[42][8] ), .C2(n16475), .A(n11669), .ZN(n11662) );
  OAI22_X1 U6318 ( .A1(n16472), .A2(n15217), .B1(n16469), .B2(n14336), .ZN(
        n11669) );
  AOI221_X1 U6319 ( .B1(\registers[50][9] ), .B2(n16529), .C1(net227065), .C2(
        n16526), .A(n11618), .ZN(n11611) );
  OAI22_X1 U6320 ( .A1(n16523), .A2(n12409), .B1(n16520), .B2(n14945), .ZN(
        n11618) );
  AOI221_X1 U6321 ( .B1(\registers[7][9] ), .B2(n16478), .C1(
        \registers[42][9] ), .C2(n16475), .A(n11626), .ZN(n11619) );
  OAI22_X1 U6322 ( .A1(n16472), .A2(n15218), .B1(n16469), .B2(n14337), .ZN(
        n11626) );
  AOI221_X1 U6323 ( .B1(\registers[50][10] ), .B2(n16529), .C1(net227083), 
        .C2(n16526), .A(n11575), .ZN(n11568) );
  OAI22_X1 U6324 ( .A1(n16523), .A2(n12411), .B1(n16520), .B2(n14946), .ZN(
        n11575) );
  AOI221_X1 U6325 ( .B1(\registers[7][10] ), .B2(n16478), .C1(
        \registers[42][10] ), .C2(n16475), .A(n11583), .ZN(n11576) );
  OAI22_X1 U6326 ( .A1(n16472), .A2(n15219), .B1(n16469), .B2(n14338), .ZN(
        n11583) );
  AOI221_X1 U6327 ( .B1(\registers[50][11] ), .B2(n16529), .C1(net227101), 
        .C2(n16526), .A(n11532), .ZN(n11525) );
  OAI22_X1 U6328 ( .A1(n16523), .A2(n12600), .B1(n16520), .B2(n14947), .ZN(
        n11532) );
  AOI221_X1 U6329 ( .B1(\registers[7][11] ), .B2(n16478), .C1(
        \registers[42][11] ), .C2(n16475), .A(n11540), .ZN(n11533) );
  OAI22_X1 U6330 ( .A1(n16472), .A2(n15220), .B1(n16469), .B2(n14339), .ZN(
        n11540) );
  AOI221_X1 U6331 ( .B1(\registers[50][12] ), .B2(n16530), .C1(net227119), 
        .C2(n16527), .A(n11489), .ZN(n11482) );
  OAI22_X1 U6332 ( .A1(n16524), .A2(n12652), .B1(n16521), .B2(n14948), .ZN(
        n11489) );
  AOI221_X1 U6333 ( .B1(\registers[7][12] ), .B2(n16479), .C1(
        \registers[42][12] ), .C2(n16476), .A(n11497), .ZN(n11490) );
  OAI22_X1 U6334 ( .A1(n16473), .A2(n15221), .B1(n16470), .B2(n14340), .ZN(
        n11497) );
  AOI221_X1 U6335 ( .B1(\registers[50][13] ), .B2(n16530), .C1(net227137), 
        .C2(n16527), .A(n11445), .ZN(n11438) );
  OAI22_X1 U6336 ( .A1(n16524), .A2(n13996), .B1(n16521), .B2(n14949), .ZN(
        n11445) );
  AOI221_X1 U6337 ( .B1(\registers[7][13] ), .B2(n16479), .C1(
        \registers[42][13] ), .C2(n16476), .A(n11453), .ZN(n11446) );
  OAI22_X1 U6338 ( .A1(n16473), .A2(n15222), .B1(n16470), .B2(n14341), .ZN(
        n11453) );
  AOI221_X1 U6339 ( .B1(\registers[50][14] ), .B2(n16530), .C1(net227155), 
        .C2(n16527), .A(n11402), .ZN(n11395) );
  OAI22_X1 U6340 ( .A1(n16524), .A2(n14008), .B1(n16521), .B2(n14950), .ZN(
        n11402) );
  AOI221_X1 U6341 ( .B1(\registers[7][14] ), .B2(n16479), .C1(
        \registers[42][14] ), .C2(n16476), .A(n11410), .ZN(n11403) );
  OAI22_X1 U6342 ( .A1(n16473), .A2(n15223), .B1(n16470), .B2(n14342), .ZN(
        n11410) );
  AOI221_X1 U6343 ( .B1(\registers[50][15] ), .B2(n16530), .C1(net227173), 
        .C2(n16527), .A(n11359), .ZN(n11352) );
  OAI22_X1 U6344 ( .A1(n16524), .A2(n14015), .B1(n16521), .B2(n14951), .ZN(
        n11359) );
  AOI221_X1 U6345 ( .B1(\registers[7][15] ), .B2(n16479), .C1(
        \registers[42][15] ), .C2(n16476), .A(n11367), .ZN(n11360) );
  OAI22_X1 U6346 ( .A1(n16473), .A2(n15224), .B1(n16470), .B2(n14343), .ZN(
        n11367) );
  AOI221_X1 U6347 ( .B1(\registers[50][16] ), .B2(n16530), .C1(net227191), 
        .C2(n16527), .A(n11316), .ZN(n11309) );
  OAI22_X1 U6348 ( .A1(n16524), .A2(n14035), .B1(n16521), .B2(n14952), .ZN(
        n11316) );
  AOI221_X1 U6349 ( .B1(\registers[7][16] ), .B2(n16479), .C1(
        \registers[42][16] ), .C2(n16476), .A(n11324), .ZN(n11317) );
  OAI22_X1 U6350 ( .A1(n16473), .A2(n15225), .B1(n16470), .B2(n14344), .ZN(
        n11324) );
  AOI221_X1 U6351 ( .B1(\registers[50][17] ), .B2(n16530), .C1(net227209), 
        .C2(n16527), .A(n11273), .ZN(n11266) );
  OAI22_X1 U6352 ( .A1(n16524), .A2(n14037), .B1(n16521), .B2(n14953), .ZN(
        n11273) );
  AOI221_X1 U6353 ( .B1(\registers[7][17] ), .B2(n16479), .C1(
        \registers[42][17] ), .C2(n16476), .A(n11281), .ZN(n11274) );
  OAI22_X1 U6354 ( .A1(n16473), .A2(n15226), .B1(n16470), .B2(n14345), .ZN(
        n11281) );
  AOI221_X1 U6355 ( .B1(\registers[50][18] ), .B2(n16530), .C1(net227227), 
        .C2(n16527), .A(n11230), .ZN(n11223) );
  OAI22_X1 U6356 ( .A1(n16524), .A2(n14039), .B1(n16521), .B2(n14954), .ZN(
        n11230) );
  AOI221_X1 U6357 ( .B1(\registers[7][18] ), .B2(n16479), .C1(
        \registers[42][18] ), .C2(n16476), .A(n11238), .ZN(n11231) );
  OAI22_X1 U6358 ( .A1(n16473), .A2(n15227), .B1(n16470), .B2(n14346), .ZN(
        n11238) );
  AOI221_X1 U6359 ( .B1(\registers[50][19] ), .B2(n16530), .C1(net227245), 
        .C2(n16527), .A(n11187), .ZN(n11180) );
  OAI22_X1 U6360 ( .A1(n16524), .A2(n14041), .B1(n16521), .B2(n14955), .ZN(
        n11187) );
  AOI221_X1 U6361 ( .B1(\registers[7][19] ), .B2(n16479), .C1(
        \registers[42][19] ), .C2(n16476), .A(n11195), .ZN(n11188) );
  OAI22_X1 U6362 ( .A1(n16473), .A2(n15228), .B1(n16470), .B2(n14347), .ZN(
        n11195) );
  AOI221_X1 U6363 ( .B1(\registers[50][20] ), .B2(n16530), .C1(net227263), 
        .C2(n16527), .A(n11144), .ZN(n11137) );
  OAI22_X1 U6364 ( .A1(n16524), .A2(n14043), .B1(n16521), .B2(n14956), .ZN(
        n11144) );
  AOI221_X1 U6365 ( .B1(\registers[7][20] ), .B2(n16479), .C1(
        \registers[42][20] ), .C2(n16476), .A(n11152), .ZN(n11145) );
  OAI22_X1 U6366 ( .A1(n16473), .A2(n15229), .B1(n16470), .B2(n14348), .ZN(
        n11152) );
  AOI221_X1 U6367 ( .B1(\registers[50][21] ), .B2(n16530), .C1(net227281), 
        .C2(n16527), .A(n11101), .ZN(n11094) );
  OAI22_X1 U6368 ( .A1(n16524), .A2(n14045), .B1(n16521), .B2(n14957), .ZN(
        n11101) );
  AOI221_X1 U6369 ( .B1(\registers[7][21] ), .B2(n16479), .C1(
        \registers[42][21] ), .C2(n16476), .A(n11109), .ZN(n11102) );
  OAI22_X1 U6370 ( .A1(n16473), .A2(n15230), .B1(n16470), .B2(n14349), .ZN(
        n11109) );
  AOI221_X1 U6371 ( .B1(\registers[50][22] ), .B2(n16530), .C1(net227299), 
        .C2(n16527), .A(n11058), .ZN(n11051) );
  OAI22_X1 U6372 ( .A1(n16524), .A2(n14047), .B1(n16521), .B2(n14958), .ZN(
        n11058) );
  AOI221_X1 U6373 ( .B1(\registers[7][22] ), .B2(n16479), .C1(
        \registers[42][22] ), .C2(n16476), .A(n11066), .ZN(n11059) );
  OAI22_X1 U6374 ( .A1(n16473), .A2(n15231), .B1(n16470), .B2(n14350), .ZN(
        n11066) );
  AOI221_X1 U6375 ( .B1(\registers[50][23] ), .B2(n16530), .C1(net227317), 
        .C2(n16527), .A(n11015), .ZN(n11008) );
  OAI22_X1 U6376 ( .A1(n16524), .A2(n14049), .B1(n16521), .B2(n14959), .ZN(
        n11015) );
  AOI221_X1 U6377 ( .B1(\registers[7][23] ), .B2(n16479), .C1(
        \registers[42][23] ), .C2(n16476), .A(n11023), .ZN(n11016) );
  OAI22_X1 U6378 ( .A1(n16473), .A2(n15232), .B1(n16470), .B2(n14351), .ZN(
        n11023) );
  AOI221_X1 U6379 ( .B1(\registers[48][0] ), .B2(n17637), .C1(
        \registers[4][0] ), .C2(n17634), .A(n12406), .ZN(n12399) );
  OAI22_X1 U6380 ( .A1(n17631), .A2(n15495), .B1(n17628), .B2(n14678), .ZN(
        n12406) );
  AOI221_X1 U6381 ( .B1(\registers[23][0] ), .B2(n17781), .C1(
        \registers[22][0] ), .C2(n17778), .A(n12382), .ZN(n12375) );
  OAI22_X1 U6382 ( .A1(n17775), .A2(n12205), .B1(n17772), .B2(n14831), .ZN(
        n12382) );
  AOI221_X1 U6383 ( .B1(\registers[48][1] ), .B2(n17637), .C1(
        \registers[4][1] ), .C2(n17634), .A(n12252), .ZN(n12245) );
  OAI22_X1 U6384 ( .A1(n17631), .A2(n15496), .B1(n17628), .B2(n14679), .ZN(
        n12252) );
  AOI221_X1 U6385 ( .B1(\registers[23][1] ), .B2(n17781), .C1(
        \registers[22][1] ), .C2(n17778), .A(n12228), .ZN(n12221) );
  OAI22_X1 U6386 ( .A1(n17775), .A2(n12206), .B1(n17772), .B2(n14832), .ZN(
        n12228) );
  AOI221_X1 U6387 ( .B1(\registers[48][2] ), .B2(n17637), .C1(
        \registers[4][2] ), .C2(n17634), .A(n12097), .ZN(n12090) );
  OAI22_X1 U6388 ( .A1(n17631), .A2(n15497), .B1(n17628), .B2(n14680), .ZN(
        n12097) );
  AOI221_X1 U6389 ( .B1(\registers[23][2] ), .B2(n17781), .C1(
        \registers[22][2] ), .C2(n17778), .A(n12073), .ZN(n12066) );
  OAI22_X1 U6390 ( .A1(n17775), .A2(n12207), .B1(n17772), .B2(n14833), .ZN(
        n12073) );
  AOI221_X1 U6391 ( .B1(\registers[48][3] ), .B2(n17637), .C1(
        \registers[4][3] ), .C2(n17634), .A(n11944), .ZN(n11937) );
  OAI22_X1 U6392 ( .A1(n17631), .A2(n15498), .B1(n17628), .B2(n14638), .ZN(
        n11944) );
  AOI221_X1 U6393 ( .B1(\registers[23][3] ), .B2(n17781), .C1(
        \registers[22][3] ), .C2(n17778), .A(n11920), .ZN(n11913) );
  OAI22_X1 U6394 ( .A1(n17775), .A2(n12208), .B1(n17772), .B2(n14834), .ZN(
        n11920) );
  AOI221_X1 U6395 ( .B1(\registers[48][4] ), .B2(n17637), .C1(
        \registers[4][4] ), .C2(n17634), .A(n10501), .ZN(n10494) );
  OAI22_X1 U6396 ( .A1(n17631), .A2(n15499), .B1(n17628), .B2(n14639), .ZN(
        n10501) );
  AOI221_X1 U6397 ( .B1(\registers[23][4] ), .B2(n17781), .C1(
        \registers[22][4] ), .C2(n17778), .A(n10477), .ZN(n10470) );
  OAI22_X1 U6398 ( .A1(n17775), .A2(n12195), .B1(n17772), .B2(n14823), .ZN(
        n10477) );
  AOI221_X1 U6399 ( .B1(\registers[48][5] ), .B2(n17637), .C1(
        \registers[4][5] ), .C2(n17634), .A(n10391), .ZN(n10384) );
  OAI22_X1 U6400 ( .A1(n17631), .A2(n15358), .B1(n17628), .B2(n14681), .ZN(
        n10391) );
  AOI221_X1 U6401 ( .B1(\registers[23][5] ), .B2(n17781), .C1(
        \registers[22][5] ), .C2(n17778), .A(n10367), .ZN(n10360) );
  OAI22_X1 U6402 ( .A1(n17775), .A2(n12209), .B1(n17772), .B2(n14835), .ZN(
        n10367) );
  AOI221_X1 U6403 ( .B1(\registers[48][6] ), .B2(n17637), .C1(
        \registers[4][6] ), .C2(n17634), .A(n10279), .ZN(n10272) );
  OAI22_X1 U6404 ( .A1(n17631), .A2(n15500), .B1(n17628), .B2(n14682), .ZN(
        n10279) );
  AOI221_X1 U6405 ( .B1(\registers[23][6] ), .B2(n17781), .C1(
        \registers[22][6] ), .C2(n17778), .A(n10255), .ZN(n10248) );
  OAI22_X1 U6406 ( .A1(n17775), .A2(n12210), .B1(n17772), .B2(n14836), .ZN(
        n10255) );
  AOI221_X1 U6407 ( .B1(\registers[48][7] ), .B2(n17637), .C1(
        \registers[4][7] ), .C2(n17634), .A(n7643), .ZN(n7636) );
  OAI22_X1 U6408 ( .A1(n17631), .A2(n15501), .B1(n17628), .B2(n14683), .ZN(
        n7643) );
  AOI221_X1 U6409 ( .B1(\registers[23][7] ), .B2(n17781), .C1(
        \registers[22][7] ), .C2(n17778), .A(n7619), .ZN(n7612) );
  OAI22_X1 U6410 ( .A1(n17775), .A2(n12211), .B1(n17772), .B2(n14837), .ZN(
        n7619) );
  AOI221_X1 U6411 ( .B1(\registers[48][8] ), .B2(n17637), .C1(
        \registers[4][8] ), .C2(n17634), .A(n7528), .ZN(n7521) );
  OAI22_X1 U6412 ( .A1(n17631), .A2(n15502), .B1(n17628), .B2(n14684), .ZN(
        n7528) );
  AOI221_X1 U6413 ( .B1(\registers[23][8] ), .B2(n17781), .C1(
        \registers[22][8] ), .C2(n17778), .A(n7504), .ZN(n7497) );
  OAI22_X1 U6414 ( .A1(n17775), .A2(n12212), .B1(n17772), .B2(n14838), .ZN(
        n7504) );
  AOI221_X1 U6415 ( .B1(\registers[48][9] ), .B2(n17637), .C1(
        \registers[4][9] ), .C2(n17634), .A(n7419), .ZN(n7412) );
  OAI22_X1 U6416 ( .A1(n17631), .A2(n15503), .B1(n17628), .B2(n14685), .ZN(
        n7419) );
  AOI221_X1 U6417 ( .B1(\registers[23][9] ), .B2(n17781), .C1(
        \registers[22][9] ), .C2(n17778), .A(n7395), .ZN(n7388) );
  OAI22_X1 U6418 ( .A1(n17775), .A2(n12213), .B1(n17772), .B2(n14839), .ZN(
        n7395) );
  AOI221_X1 U6419 ( .B1(\registers[48][10] ), .B2(n17637), .C1(
        \registers[4][10] ), .C2(n17634), .A(n7310), .ZN(n7303) );
  OAI22_X1 U6420 ( .A1(n17631), .A2(n15504), .B1(n17628), .B2(n14686), .ZN(
        n7310) );
  AOI221_X1 U6421 ( .B1(\registers[23][10] ), .B2(n17781), .C1(
        \registers[22][10] ), .C2(n17778), .A(n7286), .ZN(n7279) );
  OAI22_X1 U6422 ( .A1(n17775), .A2(n12214), .B1(n17772), .B2(n14840), .ZN(
        n7286) );
  AOI221_X1 U6423 ( .B1(\registers[48][11] ), .B2(n17638), .C1(
        \registers[4][11] ), .C2(n17635), .A(n7196), .ZN(n7189) );
  OAI22_X1 U6424 ( .A1(n17632), .A2(n15505), .B1(n17629), .B2(n14687), .ZN(
        n7196) );
  AOI221_X1 U6425 ( .B1(\registers[23][11] ), .B2(n17782), .C1(
        \registers[22][11] ), .C2(n17779), .A(n7172), .ZN(n7165) );
  OAI22_X1 U6426 ( .A1(n17776), .A2(n12215), .B1(n17773), .B2(n14841), .ZN(
        n7172) );
  AOI221_X1 U6427 ( .B1(\registers[48][12] ), .B2(n17638), .C1(
        \registers[4][12] ), .C2(n17635), .A(n7087), .ZN(n7080) );
  OAI22_X1 U6428 ( .A1(n17632), .A2(n15506), .B1(n17629), .B2(n14688), .ZN(
        n7087) );
  AOI221_X1 U6429 ( .B1(\registers[23][12] ), .B2(n17782), .C1(
        \registers[22][12] ), .C2(n17779), .A(n7063), .ZN(n7056) );
  OAI22_X1 U6430 ( .A1(n17776), .A2(n12253), .B1(n17773), .B2(n14842), .ZN(
        n7063) );
  AOI221_X1 U6431 ( .B1(\registers[48][13] ), .B2(n17638), .C1(
        \registers[4][13] ), .C2(n17635), .A(n6978), .ZN(n6971) );
  OAI22_X1 U6432 ( .A1(n17632), .A2(n15507), .B1(n17629), .B2(n14689), .ZN(
        n6978) );
  AOI221_X1 U6433 ( .B1(\registers[23][13] ), .B2(n17782), .C1(
        \registers[22][13] ), .C2(n17779), .A(n6954), .ZN(n6947) );
  OAI22_X1 U6434 ( .A1(n17776), .A2(n12254), .B1(n17773), .B2(n14843), .ZN(
        n6954) );
  AOI221_X1 U6435 ( .B1(\registers[48][14] ), .B2(n17638), .C1(
        \registers[4][14] ), .C2(n17635), .A(n6869), .ZN(n6862) );
  OAI22_X1 U6436 ( .A1(n17632), .A2(n15508), .B1(n17629), .B2(n14690), .ZN(
        n6869) );
  AOI221_X1 U6437 ( .B1(\registers[23][14] ), .B2(n17782), .C1(
        \registers[22][14] ), .C2(n17779), .A(n6845), .ZN(n6838) );
  OAI22_X1 U6438 ( .A1(n17776), .A2(n12255), .B1(n17773), .B2(n14844), .ZN(
        n6845) );
  AOI221_X1 U6439 ( .B1(\registers[48][15] ), .B2(n17638), .C1(
        \registers[4][15] ), .C2(n17635), .A(n6760), .ZN(n6753) );
  OAI22_X1 U6440 ( .A1(n17632), .A2(n15509), .B1(n17629), .B2(n14691), .ZN(
        n6760) );
  AOI221_X1 U6441 ( .B1(\registers[23][15] ), .B2(n17782), .C1(
        \registers[22][15] ), .C2(n17779), .A(n6736), .ZN(n6729) );
  OAI22_X1 U6442 ( .A1(n17776), .A2(n12256), .B1(n17773), .B2(n14845), .ZN(
        n6736) );
  AOI221_X1 U6443 ( .B1(\registers[48][16] ), .B2(n17638), .C1(
        \registers[4][16] ), .C2(n17635), .A(n6622), .ZN(n6612) );
  OAI22_X1 U6444 ( .A1(n17632), .A2(n15510), .B1(n17629), .B2(n14692), .ZN(
        n6622) );
  AOI221_X1 U6445 ( .B1(\registers[23][16] ), .B2(n17782), .C1(
        \registers[22][16] ), .C2(n17779), .A(n6576), .ZN(n6566) );
  OAI22_X1 U6446 ( .A1(n17776), .A2(n12257), .B1(n17773), .B2(n14846), .ZN(
        n6576) );
  AOI221_X1 U6447 ( .B1(\registers[48][17] ), .B2(n17638), .C1(
        \registers[4][17] ), .C2(n17635), .A(n6436), .ZN(n6426) );
  OAI22_X1 U6448 ( .A1(n17632), .A2(n15511), .B1(n17629), .B2(n14693), .ZN(
        n6436) );
  AOI221_X1 U6449 ( .B1(\registers[23][17] ), .B2(n17782), .C1(
        \registers[22][17] ), .C2(n17779), .A(n6391), .ZN(n6381) );
  OAI22_X1 U6450 ( .A1(n17776), .A2(n12258), .B1(n17773), .B2(n14847), .ZN(
        n6391) );
  AOI221_X1 U6451 ( .B1(\registers[48][18] ), .B2(n17638), .C1(
        \registers[4][18] ), .C2(n17635), .A(n6249), .ZN(n6239) );
  OAI22_X1 U6452 ( .A1(n17632), .A2(n15512), .B1(n17629), .B2(n14694), .ZN(
        n6249) );
  AOI221_X1 U6453 ( .B1(\registers[23][18] ), .B2(n17782), .C1(
        \registers[22][18] ), .C2(n17779), .A(n6204), .ZN(n6195) );
  OAI22_X1 U6454 ( .A1(n17776), .A2(n12301), .B1(n17773), .B2(n14848), .ZN(
        n6204) );
  AOI221_X1 U6455 ( .B1(\registers[48][19] ), .B2(n17638), .C1(
        \registers[4][19] ), .C2(n17635), .A(n6062), .ZN(n6052) );
  OAI22_X1 U6456 ( .A1(n17632), .A2(n15513), .B1(n17629), .B2(n14695), .ZN(
        n6062) );
  AOI221_X1 U6457 ( .B1(\registers[23][19] ), .B2(n17782), .C1(
        \registers[22][19] ), .C2(n17779), .A(n6032), .ZN(n6008) );
  OAI22_X1 U6458 ( .A1(n17776), .A2(n12303), .B1(n17773), .B2(n14849), .ZN(
        n6032) );
  AOI221_X1 U6459 ( .B1(\registers[48][20] ), .B2(n17638), .C1(
        \registers[4][20] ), .C2(n17635), .A(n5877), .ZN(n5867) );
  OAI22_X1 U6460 ( .A1(n17632), .A2(n15514), .B1(n17629), .B2(n14696), .ZN(
        n5877) );
  AOI221_X1 U6461 ( .B1(\registers[23][20] ), .B2(n17782), .C1(
        \registers[22][20] ), .C2(n17779), .A(n5845), .ZN(n5821) );
  OAI22_X1 U6462 ( .A1(n17776), .A2(n12304), .B1(n17773), .B2(n14850), .ZN(
        n5845) );
  AOI221_X1 U6463 ( .B1(\registers[48][21] ), .B2(n17638), .C1(
        \registers[4][21] ), .C2(n17635), .A(n5691), .ZN(n5681) );
  OAI22_X1 U6464 ( .A1(n17632), .A2(n15515), .B1(n17629), .B2(n14697), .ZN(
        n5691) );
  AOI221_X1 U6465 ( .B1(\registers[23][21] ), .B2(n17782), .C1(
        \registers[22][21] ), .C2(n17779), .A(n5658), .ZN(n5636) );
  OAI22_X1 U6466 ( .A1(n17776), .A2(n12305), .B1(n17773), .B2(n14851), .ZN(
        n5658) );
  AOI221_X1 U6467 ( .B1(\registers[48][22] ), .B2(n17638), .C1(
        \registers[4][22] ), .C2(n17635), .A(n5504), .ZN(n5494) );
  OAI22_X1 U6468 ( .A1(n17632), .A2(n15516), .B1(n17629), .B2(n14698), .ZN(
        n5504) );
  AOI221_X1 U6469 ( .B1(\registers[23][22] ), .B2(n17782), .C1(
        \registers[22][22] ), .C2(n17779), .A(n5471), .ZN(n5464) );
  OAI22_X1 U6470 ( .A1(n17776), .A2(n12306), .B1(n17773), .B2(n14852), .ZN(
        n5471) );
  AOI221_X1 U6471 ( .B1(\registers[48][31] ), .B2(n17637), .C1(
        \registers[4][31] ), .C2(n17634), .A(n14210), .ZN(n14187) );
  OAI22_X1 U6472 ( .A1(n17631), .A2(n15517), .B1(n17628), .B2(n14699), .ZN(
        n14210) );
  AOI221_X1 U6473 ( .B1(\registers[23][31] ), .B2(n17781), .C1(
        \registers[22][31] ), .C2(n17778), .A(n14106), .ZN(n14080) );
  OAI22_X1 U6474 ( .A1(n17775), .A2(n12307), .B1(n17772), .B2(n14853), .ZN(
        n14106) );
  NOR2_X1 U6475 ( .A1(n14097), .A2(call), .ZN(n14092) );
  NOR2_X1 U6476 ( .A1(n14003), .A2(\r590/carry[5] ), .ZN(n14196) );
  NOR2_X1 U6477 ( .A1(N9909), .A2(n10190), .ZN(n14129) );
  AOI21_X1 U6478 ( .B1(n14103), .B2(n14095), .A(n14192), .ZN(n4223) );
  AND3_X1 U6479 ( .A1(n14193), .A2(call), .A3(n14194), .ZN(n14192) );
  AOI22_X1 U6480 ( .A1(net226843), .A2(n16466), .B1(\registers[68][0] ), .B2(
        n16463), .ZN(n12416) );
  AOI221_X1 U6481 ( .B1(net226842), .B2(n16687), .C1(net226833), .C2(n16682), 
        .A(n12419), .ZN(n12418) );
  AOI221_X1 U6482 ( .B1(net226835), .B2(n16675), .C1(net226834), .C2(n16670), 
        .A(n12425), .ZN(n12417) );
  AOI22_X1 U6483 ( .A1(net227456), .A2(n16466), .B1(\registers[68][31] ), .B2(
        n16463), .ZN(n10513) );
  AOI221_X1 U6484 ( .B1(net227454), .B2(n16687), .C1(net227453), .C2(n16682), 
        .A(n10518), .ZN(n10515) );
  AOI221_X1 U6485 ( .B1(net227457), .B2(n16675), .C1(net227455), .C2(n16670), 
        .A(n10524), .ZN(n10514) );
  AOI22_X1 U6486 ( .A1(n16216), .A2(net227330), .B1(n16211), .B2(
        \registers[68][24] ), .ZN(n12889) );
  AOI221_X1 U6487 ( .B1(n16435), .B2(net227328), .C1(n16432), .C2(net227327), 
        .A(n12892), .ZN(n12891) );
  AOI221_X1 U6488 ( .B1(n16423), .B2(net227331), .C1(n16420), .C2(net227329), 
        .A(n12893), .ZN(n12890) );
  AOI22_X1 U6489 ( .A1(n16216), .A2(net227348), .B1(n16211), .B2(
        \registers[68][25] ), .ZN(n12847) );
  AOI221_X1 U6490 ( .B1(n16435), .B2(net227346), .C1(n16432), .C2(net227345), 
        .A(n12850), .ZN(n12849) );
  AOI221_X1 U6491 ( .B1(n16423), .B2(net227349), .C1(n16420), .C2(net227347), 
        .A(n12851), .ZN(n12848) );
  AOI22_X1 U6492 ( .A1(n16216), .A2(net227366), .B1(n16211), .B2(
        \registers[68][26] ), .ZN(n12805) );
  AOI221_X1 U6493 ( .B1(n16435), .B2(net227364), .C1(n16432), .C2(net227363), 
        .A(n12808), .ZN(n12807) );
  AOI221_X1 U6494 ( .B1(n16423), .B2(net227367), .C1(n16420), .C2(net227365), 
        .A(n12809), .ZN(n12806) );
  AOI22_X1 U6495 ( .A1(n16216), .A2(net227384), .B1(n16211), .B2(
        \registers[68][27] ), .ZN(n12763) );
  AOI221_X1 U6496 ( .B1(n16435), .B2(net227382), .C1(n16432), .C2(net227381), 
        .A(n12766), .ZN(n12765) );
  AOI221_X1 U6497 ( .B1(n16423), .B2(net227385), .C1(n16420), .C2(net227383), 
        .A(n12767), .ZN(n12764) );
  AOI22_X1 U6498 ( .A1(n16216), .A2(net227402), .B1(n16211), .B2(
        \registers[68][28] ), .ZN(n12721) );
  AOI221_X1 U6499 ( .B1(n16435), .B2(net227400), .C1(n16432), .C2(net227399), 
        .A(n12724), .ZN(n12723) );
  AOI221_X1 U6500 ( .B1(n16423), .B2(net227403), .C1(n16420), .C2(net227401), 
        .A(n12725), .ZN(n12722) );
  AOI22_X1 U6501 ( .A1(n16216), .A2(net227420), .B1(n16211), .B2(
        \registers[68][29] ), .ZN(n12679) );
  AOI221_X1 U6502 ( .B1(n16435), .B2(net227418), .C1(n16432), .C2(net227417), 
        .A(n12682), .ZN(n12681) );
  AOI221_X1 U6503 ( .B1(n16423), .B2(net227421), .C1(n16420), .C2(net227419), 
        .A(n12683), .ZN(n12680) );
  AOI22_X1 U6504 ( .A1(n16216), .A2(net227438), .B1(n16211), .B2(
        \registers[68][30] ), .ZN(n12635) );
  AOI221_X1 U6505 ( .B1(n16435), .B2(net227436), .C1(n16432), .C2(net227435), 
        .A(n12638), .ZN(n12637) );
  AOI221_X1 U6506 ( .B1(n16423), .B2(net227439), .C1(n16420), .C2(net227437), 
        .A(n12639), .ZN(n12636) );
  AOI22_X1 U6507 ( .A1(n16216), .A2(net227456), .B1(n16211), .B2(
        \registers[68][31] ), .ZN(n12516) );
  AOI221_X1 U6508 ( .B1(n16435), .B2(net227454), .C1(n16432), .C2(net227453), 
        .A(n12521), .ZN(n12518) );
  AOI221_X1 U6509 ( .B1(n16423), .B2(net227457), .C1(n16420), .C2(net227455), 
        .A(n12526), .ZN(n12517) );
  AOI22_X1 U6510 ( .A1(n16468), .A2(net226988), .B1(n16465), .B2(
        \registers[68][5] ), .ZN(n11757) );
  AOI221_X1 U6511 ( .B1(n16687), .B2(net226986), .C1(n16684), .C2(net226985), 
        .A(n11760), .ZN(n11759) );
  AOI221_X1 U6512 ( .B1(n16675), .B2(net226989), .C1(n16672), .C2(net226987), 
        .A(n11761), .ZN(n11758) );
  AOI22_X1 U6513 ( .A1(n16468), .A2(net227006), .B1(n16465), .B2(
        \registers[68][6] ), .ZN(n11714) );
  AOI221_X1 U6514 ( .B1(n16687), .B2(net227004), .C1(n16684), .C2(net227003), 
        .A(n11717), .ZN(n11716) );
  AOI221_X1 U6515 ( .B1(n16675), .B2(net227007), .C1(n16672), .C2(net227005), 
        .A(n11718), .ZN(n11715) );
  NOR2_X1 U6516 ( .A1(n14201), .A2(call), .ZN(n14152) );
  AOI21_X1 U6517 ( .B1(n14151), .B2(n14092), .A(n14169), .ZN(n4202) );
  AND3_X1 U6518 ( .A1(n14140), .A2(call), .A3(n14170), .ZN(n14169) );
  NOR2_X1 U6519 ( .A1(n10189), .A2(n10187), .ZN(n14128) );
  NOR2_X1 U6520 ( .A1(N9908), .A2(n10187), .ZN(n14146) );
  OAI21_X1 U6521 ( .B1(n14090), .B2(n14201), .A(n14211), .ZN(n4240) );
  NOR2_X1 U6522 ( .A1(n14089), .A2(call), .ZN(n14149) );
  NOR2_X1 U6523 ( .A1(n14098), .A2(call), .ZN(n14150) );
  AOI221_X1 U6524 ( .B1(\registers[56][23] ), .B2(n17675), .C1(
        \registers[55][23] ), .C2(n17672), .A(n5314), .ZN(n5313) );
  OAI22_X1 U6525 ( .A1(n17669), .A2(n15518), .B1(n17666), .B2(n14817), .ZN(
        n5314) );
  AOI221_X1 U6526 ( .B1(\registers[56][24] ), .B2(n17675), .C1(
        \registers[55][24] ), .C2(n17672), .A(n5142), .ZN(n5141) );
  OAI22_X1 U6527 ( .A1(n17669), .A2(n15519), .B1(n17666), .B2(n14818), .ZN(
        n5142) );
  AOI221_X1 U6528 ( .B1(\registers[56][25] ), .B2(n17675), .C1(
        \registers[55][25] ), .C2(n17672), .A(n5028), .ZN(n5027) );
  OAI22_X1 U6529 ( .A1(n17669), .A2(n15520), .B1(n17666), .B2(n14819), .ZN(
        n5028) );
  AOI221_X1 U6530 ( .B1(\registers[56][30] ), .B2(n17675), .C1(
        \registers[55][30] ), .C2(n17672), .A(n4221), .ZN(n4218) );
  OAI22_X1 U6531 ( .A1(n17669), .A2(n15315), .B1(n17666), .B2(n14632), .ZN(
        n4221) );
  AOI221_X1 U6532 ( .B1(net227344), .B2(n16315), .C1(\registers[44][24] ), 
        .C2(n16312), .A(n12919), .ZN(n12918) );
  OAI22_X1 U6533 ( .A1(n16309), .A2(n15144), .B1(n16306), .B2(n14527), .ZN(
        n12919) );
  AOI221_X1 U6534 ( .B1(\registers[7][24] ), .B2(n16228), .C1(
        \registers[42][24] ), .C2(n16225), .A(n12930), .ZN(n12923) );
  OAI22_X1 U6535 ( .A1(n16222), .A2(n15233), .B1(n16219), .B2(n14352), .ZN(
        n12930) );
  AOI221_X1 U6536 ( .B1(net227362), .B2(n16315), .C1(\registers[44][25] ), 
        .C2(n16312), .A(n12877), .ZN(n12876) );
  OAI22_X1 U6537 ( .A1(n16309), .A2(n15145), .B1(n16306), .B2(n14528), .ZN(
        n12877) );
  AOI221_X1 U6538 ( .B1(\registers[7][25] ), .B2(n16228), .C1(
        \registers[42][25] ), .C2(n16225), .A(n12888), .ZN(n12881) );
  OAI22_X1 U6539 ( .A1(n16222), .A2(n15234), .B1(n16219), .B2(n14353), .ZN(
        n12888) );
  AOI221_X1 U6540 ( .B1(net227380), .B2(n16315), .C1(\registers[44][26] ), 
        .C2(n16312), .A(n12835), .ZN(n12834) );
  OAI22_X1 U6541 ( .A1(n16309), .A2(n15146), .B1(n16306), .B2(n14529), .ZN(
        n12835) );
  AOI221_X1 U6542 ( .B1(\registers[7][26] ), .B2(n16228), .C1(
        \registers[42][26] ), .C2(n16225), .A(n12846), .ZN(n12839) );
  OAI22_X1 U6543 ( .A1(n16222), .A2(n15235), .B1(n16219), .B2(n14354), .ZN(
        n12846) );
  AOI221_X1 U6544 ( .B1(net227398), .B2(n16315), .C1(\registers[44][27] ), 
        .C2(n16312), .A(n12793), .ZN(n12792) );
  OAI22_X1 U6545 ( .A1(n16309), .A2(n15147), .B1(n16306), .B2(n14530), .ZN(
        n12793) );
  AOI221_X1 U6546 ( .B1(\registers[7][27] ), .B2(n16228), .C1(
        \registers[42][27] ), .C2(n16225), .A(n12804), .ZN(n12797) );
  OAI22_X1 U6547 ( .A1(n16222), .A2(n15236), .B1(n16219), .B2(n14355), .ZN(
        n12804) );
  AOI221_X1 U6548 ( .B1(net227416), .B2(n16315), .C1(\registers[44][28] ), 
        .C2(n16312), .A(n12751), .ZN(n12750) );
  OAI22_X1 U6549 ( .A1(n16309), .A2(n15148), .B1(n16306), .B2(n14531), .ZN(
        n12751) );
  AOI221_X1 U6550 ( .B1(\registers[7][28] ), .B2(n16228), .C1(
        \registers[42][28] ), .C2(n16225), .A(n12762), .ZN(n12755) );
  OAI22_X1 U6551 ( .A1(n16222), .A2(n15237), .B1(n16219), .B2(n14356), .ZN(
        n12762) );
  AOI221_X1 U6552 ( .B1(net227434), .B2(n16315), .C1(\registers[44][29] ), 
        .C2(n16312), .A(n12709), .ZN(n12708) );
  OAI22_X1 U6553 ( .A1(n16309), .A2(n15149), .B1(n16306), .B2(n14532), .ZN(
        n12709) );
  AOI221_X1 U6554 ( .B1(\registers[7][29] ), .B2(n16228), .C1(
        \registers[42][29] ), .C2(n16225), .A(n12720), .ZN(n12713) );
  OAI22_X1 U6555 ( .A1(n16222), .A2(n15238), .B1(n16219), .B2(n14357), .ZN(
        n12720) );
  AOI221_X1 U6556 ( .B1(net227452), .B2(n16315), .C1(\registers[44][30] ), 
        .C2(n16312), .A(n12666), .ZN(n12665) );
  OAI22_X1 U6557 ( .A1(n16309), .A2(n14871), .B1(n16306), .B2(n14069), .ZN(
        n12666) );
  AOI221_X1 U6558 ( .B1(\registers[7][30] ), .B2(n16228), .C1(
        \registers[42][30] ), .C2(n16225), .A(n12678), .ZN(n12671) );
  OAI22_X1 U6559 ( .A1(n16222), .A2(n14874), .B1(n16219), .B2(n14055), .ZN(
        n12678) );
  AOI221_X1 U6560 ( .B1(net227470), .B2(n16315), .C1(\registers[44][31] ), 
        .C2(n16312), .A(n12588), .ZN(n12585) );
  OAI22_X1 U6561 ( .A1(n16309), .A2(n15150), .B1(n16306), .B2(n14533), .ZN(
        n12588) );
  AOI221_X1 U6562 ( .B1(\registers[7][31] ), .B2(n16228), .C1(
        \registers[42][31] ), .C2(n16225), .A(n12630), .ZN(n12608) );
  OAI22_X1 U6563 ( .A1(n16222), .A2(n15239), .B1(n16219), .B2(n14358), .ZN(
        n12630) );
  AOI221_X1 U6564 ( .B1(\registers[50][0] ), .B2(n16277), .C1(net226846), .C2(
        n16274), .A(n13959), .ZN(n13948) );
  OAI22_X1 U6565 ( .A1(n16271), .A2(n12356), .B1(n16268), .B2(n14938), .ZN(
        n13959) );
  AOI221_X1 U6566 ( .B1(\registers[5][0] ), .B2(n16250), .C1(
        \registers[59][0] ), .C2(n16247), .A(n13971), .ZN(n13966) );
  OAI22_X1 U6567 ( .A1(n16244), .A2(n12357), .B1(n16241), .B2(n14910), .ZN(
        n13971) );
  AOI221_X1 U6568 ( .B1(\registers[50][1] ), .B2(n16277), .C1(net226859), .C2(
        n16274), .A(n13888), .ZN(n13881) );
  OAI22_X1 U6569 ( .A1(n16271), .A2(n12358), .B1(n16268), .B2(n14939), .ZN(
        n13888) );
  AOI221_X1 U6570 ( .B1(\registers[5][1] ), .B2(n16250), .C1(
        \registers[59][1] ), .C2(n16247), .A(n13894), .ZN(n13891) );
  OAI22_X1 U6571 ( .A1(n16244), .A2(n12359), .B1(n16241), .B2(n14911), .ZN(
        n13894) );
  AOI221_X1 U6572 ( .B1(\registers[50][2] ), .B2(n16277), .C1(net226885), .C2(
        n16274), .A(n13846), .ZN(n13839) );
  OAI22_X1 U6573 ( .A1(n16271), .A2(n12360), .B1(n16268), .B2(n14940), .ZN(
        n13846) );
  AOI221_X1 U6574 ( .B1(\registers[5][2] ), .B2(n16250), .C1(
        \registers[59][2] ), .C2(n16247), .A(n13852), .ZN(n13849) );
  OAI22_X1 U6575 ( .A1(n16244), .A2(n12361), .B1(n16241), .B2(n14912), .ZN(
        n13852) );
  AOI221_X1 U6576 ( .B1(\registers[50][3] ), .B2(n16277), .C1(net226898), .C2(
        n16274), .A(n13804), .ZN(n13797) );
  OAI22_X1 U6577 ( .A1(n16271), .A2(n12340), .B1(n16268), .B2(n14941), .ZN(
        n13804) );
  AOI221_X1 U6578 ( .B1(\registers[5][3] ), .B2(n16250), .C1(
        \registers[59][3] ), .C2(n16247), .A(n13810), .ZN(n13807) );
  OAI22_X1 U6579 ( .A1(n16244), .A2(n12362), .B1(n16241), .B2(n14863), .ZN(
        n13810) );
  AOI221_X1 U6580 ( .B1(\registers[50][4] ), .B2(n16277), .C1(net226980), .C2(
        n16274), .A(n13762), .ZN(n13755) );
  OAI22_X1 U6581 ( .A1(n16271), .A2(n12341), .B1(n16268), .B2(n14866), .ZN(
        n13762) );
  AOI221_X1 U6582 ( .B1(\registers[5][4] ), .B2(n16250), .C1(
        \registers[59][4] ), .C2(n16247), .A(n13768), .ZN(n13765) );
  OAI22_X1 U6583 ( .A1(n16244), .A2(n12363), .B1(n16241), .B2(n14864), .ZN(
        n13768) );
  AOI221_X1 U6584 ( .B1(\registers[50][5] ), .B2(n16277), .C1(net227000), .C2(
        n16274), .A(n13720), .ZN(n13713) );
  OAI22_X1 U6585 ( .A1(n16271), .A2(n12364), .B1(n16268), .B2(n14867), .ZN(
        n13720) );
  AOI221_X1 U6586 ( .B1(\registers[5][5] ), .B2(n16250), .C1(
        \registers[59][5] ), .C2(n16247), .A(n13726), .ZN(n13723) );
  OAI22_X1 U6587 ( .A1(n16244), .A2(n12365), .B1(n16241), .B2(n14865), .ZN(
        n13726) );
  AOI221_X1 U6588 ( .B1(\registers[50][6] ), .B2(n16277), .C1(net227011), .C2(
        n16274), .A(n13678), .ZN(n13671) );
  OAI22_X1 U6589 ( .A1(n16271), .A2(n12366), .B1(n16268), .B2(n14942), .ZN(
        n13678) );
  AOI221_X1 U6590 ( .B1(\registers[5][6] ), .B2(n16250), .C1(
        \registers[59][6] ), .C2(n16247), .A(n13684), .ZN(n13681) );
  OAI22_X1 U6591 ( .A1(n16244), .A2(n12367), .B1(n16241), .B2(n14913), .ZN(
        n13684) );
  AOI221_X1 U6592 ( .B1(\registers[50][7] ), .B2(n16277), .C1(net227029), .C2(
        n16274), .A(n13636), .ZN(n13629) );
  OAI22_X1 U6593 ( .A1(n16271), .A2(n12368), .B1(n16268), .B2(n14943), .ZN(
        n13636) );
  AOI221_X1 U6594 ( .B1(\registers[5][7] ), .B2(n16250), .C1(
        \registers[59][7] ), .C2(n16247), .A(n13642), .ZN(n13639) );
  OAI22_X1 U6595 ( .A1(n16244), .A2(n12369), .B1(n16241), .B2(n14914), .ZN(
        n13642) );
  AOI221_X1 U6596 ( .B1(\registers[50][8] ), .B2(n16277), .C1(net227047), .C2(
        n16274), .A(n13594), .ZN(n13587) );
  OAI22_X1 U6597 ( .A1(n16271), .A2(n12407), .B1(n16268), .B2(n14944), .ZN(
        n13594) );
  AOI221_X1 U6598 ( .B1(\registers[5][8] ), .B2(n16250), .C1(
        \registers[59][8] ), .C2(n16247), .A(n13600), .ZN(n13597) );
  OAI22_X1 U6599 ( .A1(n16244), .A2(n12408), .B1(n16241), .B2(n14915), .ZN(
        n13600) );
  AOI221_X1 U6600 ( .B1(\registers[50][9] ), .B2(n16277), .C1(net227065), .C2(
        n16274), .A(n13552), .ZN(n13545) );
  OAI22_X1 U6601 ( .A1(n16271), .A2(n12409), .B1(n16268), .B2(n14945), .ZN(
        n13552) );
  AOI221_X1 U6602 ( .B1(\registers[5][9] ), .B2(n16250), .C1(
        \registers[59][9] ), .C2(n16247), .A(n13558), .ZN(n13555) );
  OAI22_X1 U6603 ( .A1(n16244), .A2(n12410), .B1(n16241), .B2(n14916), .ZN(
        n13558) );
  AOI221_X1 U6604 ( .B1(\registers[50][10] ), .B2(n16277), .C1(net227083), 
        .C2(n16274), .A(n13510), .ZN(n13503) );
  OAI22_X1 U6605 ( .A1(n16271), .A2(n12411), .B1(n16268), .B2(n14946), .ZN(
        n13510) );
  AOI221_X1 U6606 ( .B1(\registers[5][10] ), .B2(n16250), .C1(
        \registers[59][10] ), .C2(n16247), .A(n13516), .ZN(n13513) );
  OAI22_X1 U6607 ( .A1(n16244), .A2(n12551), .B1(n16241), .B2(n14917), .ZN(
        n13516) );
  AOI221_X1 U6608 ( .B1(\registers[50][11] ), .B2(n16277), .C1(net227101), 
        .C2(n16274), .A(n13468), .ZN(n13461) );
  OAI22_X1 U6609 ( .A1(n16271), .A2(n12600), .B1(n16268), .B2(n14947), .ZN(
        n13468) );
  AOI221_X1 U6610 ( .B1(\registers[5][11] ), .B2(n16250), .C1(
        \registers[59][11] ), .C2(n16247), .A(n13474), .ZN(n13471) );
  OAI22_X1 U6611 ( .A1(n16244), .A2(n12602), .B1(n16241), .B2(n14918), .ZN(
        n13474) );
  AOI221_X1 U6612 ( .B1(\registers[50][12] ), .B2(n16278), .C1(net227119), 
        .C2(n16275), .A(n13426), .ZN(n13419) );
  OAI22_X1 U6613 ( .A1(n16272), .A2(n12652), .B1(n16269), .B2(n14948), .ZN(
        n13426) );
  AOI221_X1 U6614 ( .B1(\registers[5][12] ), .B2(n16251), .C1(
        \registers[59][12] ), .C2(n16248), .A(n13432), .ZN(n13429) );
  OAI22_X1 U6615 ( .A1(n16245), .A2(n12669), .B1(n16242), .B2(n14919), .ZN(
        n13432) );
  AOI221_X1 U6616 ( .B1(\registers[50][13] ), .B2(n16278), .C1(net227137), 
        .C2(n16275), .A(n13384), .ZN(n13377) );
  OAI22_X1 U6617 ( .A1(n16272), .A2(n13996), .B1(n16269), .B2(n14949), .ZN(
        n13384) );
  AOI221_X1 U6618 ( .B1(\registers[5][13] ), .B2(n16251), .C1(
        \registers[59][13] ), .C2(n16248), .A(n13390), .ZN(n13387) );
  OAI22_X1 U6619 ( .A1(n16245), .A2(n13999), .B1(n16242), .B2(n14920), .ZN(
        n13390) );
  AOI221_X1 U6620 ( .B1(\registers[50][14] ), .B2(n16278), .C1(net227155), 
        .C2(n16275), .A(n13342), .ZN(n13335) );
  OAI22_X1 U6621 ( .A1(n16272), .A2(n14008), .B1(n16269), .B2(n14950), .ZN(
        n13342) );
  AOI221_X1 U6622 ( .B1(\registers[5][14] ), .B2(n16251), .C1(
        \registers[59][14] ), .C2(n16248), .A(n13348), .ZN(n13345) );
  OAI22_X1 U6623 ( .A1(n16245), .A2(n14014), .B1(n16242), .B2(n14921), .ZN(
        n13348) );
  AOI221_X1 U6624 ( .B1(\registers[50][15] ), .B2(n16278), .C1(net227173), 
        .C2(n16275), .A(n13300), .ZN(n13293) );
  OAI22_X1 U6625 ( .A1(n16272), .A2(n14015), .B1(n16269), .B2(n14951), .ZN(
        n13300) );
  AOI221_X1 U6626 ( .B1(\registers[5][15] ), .B2(n16251), .C1(
        \registers[59][15] ), .C2(n16248), .A(n13306), .ZN(n13303) );
  OAI22_X1 U6627 ( .A1(n16245), .A2(n14032), .B1(n16242), .B2(n14922), .ZN(
        n13306) );
  AOI221_X1 U6628 ( .B1(\registers[50][16] ), .B2(n16278), .C1(net227191), 
        .C2(n16275), .A(n13258), .ZN(n13251) );
  OAI22_X1 U6629 ( .A1(n16272), .A2(n14035), .B1(n16269), .B2(n14952), .ZN(
        n13258) );
  AOI221_X1 U6630 ( .B1(\registers[5][16] ), .B2(n16251), .C1(
        \registers[59][16] ), .C2(n16248), .A(n13264), .ZN(n13261) );
  OAI22_X1 U6631 ( .A1(n16245), .A2(n14036), .B1(n16242), .B2(n14923), .ZN(
        n13264) );
  AOI221_X1 U6632 ( .B1(\registers[50][17] ), .B2(n16278), .C1(net227209), 
        .C2(n16275), .A(n13216), .ZN(n13209) );
  OAI22_X1 U6633 ( .A1(n16272), .A2(n14037), .B1(n16269), .B2(n14953), .ZN(
        n13216) );
  AOI221_X1 U6634 ( .B1(\registers[5][17] ), .B2(n16251), .C1(
        \registers[59][17] ), .C2(n16248), .A(n13222), .ZN(n13219) );
  OAI22_X1 U6635 ( .A1(n16245), .A2(n14038), .B1(n16242), .B2(n14924), .ZN(
        n13222) );
  AOI221_X1 U6636 ( .B1(\registers[50][18] ), .B2(n16278), .C1(net227227), 
        .C2(n16275), .A(n13174), .ZN(n13167) );
  OAI22_X1 U6637 ( .A1(n16272), .A2(n14039), .B1(n16269), .B2(n14954), .ZN(
        n13174) );
  AOI221_X1 U6638 ( .B1(\registers[5][18] ), .B2(n16251), .C1(
        \registers[59][18] ), .C2(n16248), .A(n13180), .ZN(n13177) );
  OAI22_X1 U6639 ( .A1(n16245), .A2(n14040), .B1(n16242), .B2(n14925), .ZN(
        n13180) );
  AOI221_X1 U6640 ( .B1(\registers[50][19] ), .B2(n16278), .C1(net227245), 
        .C2(n16275), .A(n13132), .ZN(n13125) );
  OAI22_X1 U6641 ( .A1(n16272), .A2(n14041), .B1(n16269), .B2(n14955), .ZN(
        n13132) );
  AOI221_X1 U6642 ( .B1(\registers[5][19] ), .B2(n16251), .C1(
        \registers[59][19] ), .C2(n16248), .A(n13138), .ZN(n13135) );
  OAI22_X1 U6643 ( .A1(n16245), .A2(n14042), .B1(n16242), .B2(n14926), .ZN(
        n13138) );
  AOI221_X1 U6644 ( .B1(\registers[50][20] ), .B2(n16278), .C1(net227263), 
        .C2(n16275), .A(n13090), .ZN(n13083) );
  OAI22_X1 U6645 ( .A1(n16272), .A2(n14043), .B1(n16269), .B2(n14956), .ZN(
        n13090) );
  AOI221_X1 U6646 ( .B1(\registers[5][20] ), .B2(n16251), .C1(
        \registers[59][20] ), .C2(n16248), .A(n13096), .ZN(n13093) );
  OAI22_X1 U6647 ( .A1(n16245), .A2(n14044), .B1(n16242), .B2(n14927), .ZN(
        n13096) );
  AOI221_X1 U6648 ( .B1(\registers[50][21] ), .B2(n16278), .C1(net227281), 
        .C2(n16275), .A(n13048), .ZN(n13041) );
  OAI22_X1 U6649 ( .A1(n16272), .A2(n14045), .B1(n16269), .B2(n14957), .ZN(
        n13048) );
  AOI221_X1 U6650 ( .B1(\registers[5][21] ), .B2(n16251), .C1(
        \registers[59][21] ), .C2(n16248), .A(n13054), .ZN(n13051) );
  OAI22_X1 U6651 ( .A1(n16245), .A2(n14046), .B1(n16242), .B2(n14928), .ZN(
        n13054) );
  AOI221_X1 U6652 ( .B1(\registers[50][22] ), .B2(n16278), .C1(net227299), 
        .C2(n16275), .A(n13006), .ZN(n12999) );
  OAI22_X1 U6653 ( .A1(n16272), .A2(n14047), .B1(n16269), .B2(n14958), .ZN(
        n13006) );
  AOI221_X1 U6654 ( .B1(\registers[5][22] ), .B2(n16251), .C1(
        \registers[59][22] ), .C2(n16248), .A(n13012), .ZN(n13009) );
  OAI22_X1 U6655 ( .A1(n16245), .A2(n14048), .B1(n16242), .B2(n14929), .ZN(
        n13012) );
  AOI221_X1 U6656 ( .B1(\registers[50][23] ), .B2(n16278), .C1(net227317), 
        .C2(n16275), .A(n12964), .ZN(n12957) );
  OAI22_X1 U6657 ( .A1(n16272), .A2(n14049), .B1(n16269), .B2(n14959), .ZN(
        n12964) );
  AOI221_X1 U6658 ( .B1(\registers[5][23] ), .B2(n16251), .C1(
        \registers[59][23] ), .C2(n16248), .A(n12970), .ZN(n12967) );
  OAI22_X1 U6659 ( .A1(n16245), .A2(n14050), .B1(n16242), .B2(n14930), .ZN(
        n12970) );
  AOI221_X1 U6660 ( .B1(\registers[49][0] ), .B2(n16541), .C1(
        \registers[51][0] ), .C2(n16538), .A(n12476), .ZN(n12468) );
  OAI22_X1 U6661 ( .A1(n16535), .A2(n15521), .B1(n16532), .B2(n14547), .ZN(
        n12476) );
  AOI221_X1 U6662 ( .B1(\registers[49][1] ), .B2(n16541), .C1(
        \registers[51][1] ), .C2(n16538), .A(n12291), .ZN(n12286) );
  OAI22_X1 U6663 ( .A1(n16535), .A2(n15522), .B1(n16532), .B2(n14548), .ZN(
        n12291) );
  AOI221_X1 U6664 ( .B1(\registers[49][2] ), .B2(n16541), .C1(
        \registers[51][2] ), .C2(n16538), .A(n12138), .ZN(n12133) );
  OAI22_X1 U6665 ( .A1(n16535), .A2(n15523), .B1(n16532), .B2(n14549), .ZN(
        n12138) );
  AOI221_X1 U6666 ( .B1(\registers[49][3] ), .B2(n16541), .C1(
        \registers[51][3] ), .C2(n16538), .A(n11985), .ZN(n11980) );
  OAI22_X1 U6667 ( .A1(n16535), .A2(n15524), .B1(n16532), .B2(n14536), .ZN(
        n11985) );
  AOI221_X1 U6668 ( .B1(\registers[49][4] ), .B2(n16541), .C1(
        \registers[51][4] ), .C2(n16538), .A(n11832), .ZN(n11827) );
  OAI22_X1 U6669 ( .A1(n16535), .A2(n15525), .B1(n16532), .B2(n14550), .ZN(
        n11832) );
  AOI221_X1 U6670 ( .B1(\registers[49][5] ), .B2(n16541), .C1(
        \registers[51][5] ), .C2(n16538), .A(n11789), .ZN(n11784) );
  OAI22_X1 U6671 ( .A1(n16535), .A2(n15526), .B1(n16532), .B2(n14537), .ZN(
        n11789) );
  AOI221_X1 U6672 ( .B1(\registers[49][6] ), .B2(n16541), .C1(
        \registers[51][6] ), .C2(n16538), .A(n11746), .ZN(n11741) );
  OAI22_X1 U6673 ( .A1(n16535), .A2(n15527), .B1(n16532), .B2(n14551), .ZN(
        n11746) );
  AOI221_X1 U6674 ( .B1(\registers[49][7] ), .B2(n16541), .C1(
        \registers[51][7] ), .C2(n16538), .A(n11703), .ZN(n11698) );
  OAI22_X1 U6675 ( .A1(n16535), .A2(n15528), .B1(n16532), .B2(n14552), .ZN(
        n11703) );
  AOI221_X1 U6676 ( .B1(\registers[49][8] ), .B2(n16541), .C1(
        \registers[51][8] ), .C2(n16538), .A(n11660), .ZN(n11655) );
  OAI22_X1 U6677 ( .A1(n16535), .A2(n15529), .B1(n16532), .B2(n14553), .ZN(
        n11660) );
  AOI221_X1 U6678 ( .B1(\registers[49][9] ), .B2(n16541), .C1(
        \registers[51][9] ), .C2(n16538), .A(n11617), .ZN(n11612) );
  OAI22_X1 U6679 ( .A1(n16535), .A2(n15530), .B1(n16532), .B2(n14554), .ZN(
        n11617) );
  AOI221_X1 U6680 ( .B1(\registers[49][10] ), .B2(n16541), .C1(
        \registers[51][10] ), .C2(n16538), .A(n11574), .ZN(n11569) );
  OAI22_X1 U6681 ( .A1(n16535), .A2(n15531), .B1(n16532), .B2(n14555), .ZN(
        n11574) );
  AOI221_X1 U6682 ( .B1(\registers[49][11] ), .B2(n16541), .C1(
        \registers[51][11] ), .C2(n16538), .A(n11531), .ZN(n11526) );
  OAI22_X1 U6683 ( .A1(n16535), .A2(n15532), .B1(n16532), .B2(n14556), .ZN(
        n11531) );
  AOI221_X1 U6684 ( .B1(\registers[49][12] ), .B2(n16542), .C1(
        \registers[51][12] ), .C2(n16539), .A(n11488), .ZN(n11483) );
  OAI22_X1 U6685 ( .A1(n16536), .A2(n15533), .B1(n16533), .B2(n14557), .ZN(
        n11488) );
  AOI221_X1 U6686 ( .B1(\registers[49][13] ), .B2(n16542), .C1(
        \registers[51][13] ), .C2(n16539), .A(n11444), .ZN(n11439) );
  OAI22_X1 U6687 ( .A1(n16536), .A2(n15534), .B1(n16533), .B2(n14558), .ZN(
        n11444) );
  AOI221_X1 U6688 ( .B1(\registers[49][14] ), .B2(n16542), .C1(
        \registers[51][14] ), .C2(n16539), .A(n11401), .ZN(n11396) );
  OAI22_X1 U6689 ( .A1(n16536), .A2(n15535), .B1(n16533), .B2(n14559), .ZN(
        n11401) );
  AOI221_X1 U6690 ( .B1(\registers[49][15] ), .B2(n16542), .C1(
        \registers[51][15] ), .C2(n16539), .A(n11358), .ZN(n11353) );
  OAI22_X1 U6691 ( .A1(n16536), .A2(n15536), .B1(n16533), .B2(n14560), .ZN(
        n11358) );
  AOI221_X1 U6692 ( .B1(\registers[49][16] ), .B2(n16542), .C1(
        \registers[51][16] ), .C2(n16539), .A(n11315), .ZN(n11310) );
  OAI22_X1 U6693 ( .A1(n16536), .A2(n15537), .B1(n16533), .B2(n14561), .ZN(
        n11315) );
  AOI221_X1 U6694 ( .B1(\registers[49][17] ), .B2(n16542), .C1(
        \registers[51][17] ), .C2(n16539), .A(n11272), .ZN(n11267) );
  OAI22_X1 U6695 ( .A1(n16536), .A2(n15538), .B1(n16533), .B2(n14562), .ZN(
        n11272) );
  AOI221_X1 U6696 ( .B1(\registers[49][18] ), .B2(n16542), .C1(
        \registers[51][18] ), .C2(n16539), .A(n11229), .ZN(n11224) );
  OAI22_X1 U6697 ( .A1(n16536), .A2(n15539), .B1(n16533), .B2(n14563), .ZN(
        n11229) );
  AOI221_X1 U6698 ( .B1(\registers[49][19] ), .B2(n16542), .C1(
        \registers[51][19] ), .C2(n16539), .A(n11186), .ZN(n11181) );
  OAI22_X1 U6699 ( .A1(n16536), .A2(n15540), .B1(n16533), .B2(n14564), .ZN(
        n11186) );
  AOI221_X1 U6700 ( .B1(\registers[49][20] ), .B2(n16542), .C1(
        \registers[51][20] ), .C2(n16539), .A(n11143), .ZN(n11138) );
  OAI22_X1 U6701 ( .A1(n16536), .A2(n15541), .B1(n16533), .B2(n14565), .ZN(
        n11143) );
  AOI221_X1 U6702 ( .B1(\registers[49][21] ), .B2(n16542), .C1(
        \registers[51][21] ), .C2(n16539), .A(n11100), .ZN(n11095) );
  OAI22_X1 U6703 ( .A1(n16536), .A2(n15542), .B1(n16533), .B2(n14566), .ZN(
        n11100) );
  AOI221_X1 U6704 ( .B1(\registers[49][22] ), .B2(n16542), .C1(
        \registers[51][22] ), .C2(n16539), .A(n11057), .ZN(n11052) );
  OAI22_X1 U6705 ( .A1(n16536), .A2(n15543), .B1(n16533), .B2(n14567), .ZN(
        n11057) );
  AOI221_X1 U6706 ( .B1(\registers[49][23] ), .B2(n16542), .C1(
        \registers[51][23] ), .C2(n16539), .A(n11014), .ZN(n11009) );
  OAI22_X1 U6707 ( .A1(n16536), .A2(n15544), .B1(n16533), .B2(n14568), .ZN(
        n11014) );
  AOI221_X1 U6708 ( .B1(net226841), .B2(n17697), .C1(\registers[9][0] ), .C2(
        n17694), .A(n12397), .ZN(n12392) );
  OAI22_X1 U6709 ( .A1(n17691), .A2(n15758), .B1(n17688), .B2(n12171), .ZN(
        n12397) );
  AOI221_X1 U6710 ( .B1(net226864), .B2(n17697), .C1(\registers[9][1] ), .C2(
        n17694), .A(n12243), .ZN(n12238) );
  OAI22_X1 U6711 ( .A1(n17691), .A2(n15759), .B1(n17688), .B2(n12172), .ZN(
        n12243) );
  AOI221_X1 U6712 ( .B1(net226882), .B2(n17697), .C1(\registers[9][2] ), .C2(
        n17694), .A(n12088), .ZN(n12083) );
  OAI22_X1 U6713 ( .A1(n17691), .A2(n15760), .B1(n17688), .B2(n12173), .ZN(
        n12088) );
  AOI221_X1 U6714 ( .B1(net226902), .B2(n17697), .C1(\registers[9][3] ), .C2(
        n17694), .A(n11935), .ZN(n11930) );
  OAI22_X1 U6715 ( .A1(n17691), .A2(n15761), .B1(n17688), .B2(n12174), .ZN(
        n11935) );
  AOI221_X1 U6716 ( .B1(net226975), .B2(n17697), .C1(\registers[9][4] ), .C2(
        n17694), .A(n10492), .ZN(n10487) );
  OAI22_X1 U6717 ( .A1(n17691), .A2(n15762), .B1(n17688), .B2(n12175), .ZN(
        n10492) );
  AOI221_X1 U6718 ( .B1(net226995), .B2(n17697), .C1(\registers[9][5] ), .C2(
        n17694), .A(n10382), .ZN(n10377) );
  OAI22_X1 U6719 ( .A1(n17691), .A2(n15763), .B1(n17688), .B2(n12162), .ZN(
        n10382) );
  AOI221_X1 U6720 ( .B1(net227019), .B2(n17697), .C1(\registers[9][6] ), .C2(
        n17694), .A(n10270), .ZN(n10265) );
  OAI22_X1 U6721 ( .A1(n17691), .A2(n15764), .B1(n17688), .B2(n12176), .ZN(
        n10270) );
  AOI221_X1 U6722 ( .B1(net227037), .B2(n17697), .C1(\registers[9][7] ), .C2(
        n17694), .A(n7634), .ZN(n7629) );
  OAI22_X1 U6723 ( .A1(n17691), .A2(n15765), .B1(n17688), .B2(n12177), .ZN(
        n7634) );
  AOI221_X1 U6724 ( .B1(net227055), .B2(n17697), .C1(\registers[9][8] ), .C2(
        n17694), .A(n7519), .ZN(n7514) );
  OAI22_X1 U6725 ( .A1(n17691), .A2(n15766), .B1(n17688), .B2(n12178), .ZN(
        n7519) );
  AOI221_X1 U6726 ( .B1(net227073), .B2(n17697), .C1(\registers[9][9] ), .C2(
        n17694), .A(n7410), .ZN(n7405) );
  OAI22_X1 U6727 ( .A1(n17691), .A2(n15767), .B1(n17688), .B2(n12179), .ZN(
        n7410) );
  AOI221_X1 U6728 ( .B1(net227091), .B2(n17697), .C1(\registers[9][10] ), .C2(
        n17694), .A(n7301), .ZN(n7296) );
  OAI22_X1 U6729 ( .A1(n17691), .A2(n15768), .B1(n17688), .B2(n12180), .ZN(
        n7301) );
  AOI221_X1 U6730 ( .B1(net227109), .B2(n17698), .C1(\registers[9][11] ), .C2(
        n17695), .A(n7187), .ZN(n7182) );
  OAI22_X1 U6731 ( .A1(n17692), .A2(n15769), .B1(n17689), .B2(n12181), .ZN(
        n7187) );
  AOI221_X1 U6732 ( .B1(net227127), .B2(n17698), .C1(\registers[9][12] ), .C2(
        n17695), .A(n7078), .ZN(n7073) );
  OAI22_X1 U6733 ( .A1(n17692), .A2(n15770), .B1(n17689), .B2(n12182), .ZN(
        n7078) );
  AOI221_X1 U6734 ( .B1(net227145), .B2(n17698), .C1(\registers[9][13] ), .C2(
        n17695), .A(n6969), .ZN(n6964) );
  OAI22_X1 U6735 ( .A1(n17692), .A2(n15771), .B1(n17689), .B2(n12183), .ZN(
        n6969) );
  AOI221_X1 U6736 ( .B1(net227163), .B2(n17698), .C1(\registers[9][14] ), .C2(
        n17695), .A(n6860), .ZN(n6855) );
  OAI22_X1 U6737 ( .A1(n17692), .A2(n15772), .B1(n17689), .B2(n12185), .ZN(
        n6860) );
  AOI221_X1 U6738 ( .B1(net227181), .B2(n17698), .C1(\registers[9][15] ), .C2(
        n17695), .A(n6751), .ZN(n6746) );
  OAI22_X1 U6739 ( .A1(n17692), .A2(n15773), .B1(n17689), .B2(n12186), .ZN(
        n6751) );
  AOI221_X1 U6740 ( .B1(net227199), .B2(n17698), .C1(\registers[9][16] ), .C2(
        n17695), .A(n6609), .ZN(n6603) );
  OAI22_X1 U6741 ( .A1(n17692), .A2(n15774), .B1(n17689), .B2(n12187), .ZN(
        n6609) );
  AOI221_X1 U6742 ( .B1(net227217), .B2(n17698), .C1(\registers[9][17] ), .C2(
        n17695), .A(n6423), .ZN(n6416) );
  OAI22_X1 U6743 ( .A1(n17692), .A2(n15775), .B1(n17689), .B2(n12188), .ZN(
        n6423) );
  AOI221_X1 U6744 ( .B1(net227235), .B2(n17698), .C1(\registers[9][18] ), .C2(
        n17695), .A(n6237), .ZN(n6229) );
  OAI22_X1 U6745 ( .A1(n17692), .A2(n15776), .B1(n17689), .B2(n12189), .ZN(
        n6237) );
  AOI221_X1 U6746 ( .B1(net227253), .B2(n17698), .C1(\registers[9][19] ), .C2(
        n17695), .A(n6050), .ZN(n6043) );
  OAI22_X1 U6747 ( .A1(n17692), .A2(n15777), .B1(n17689), .B2(n12190), .ZN(
        n6050) );
  AOI221_X1 U6748 ( .B1(net227271), .B2(n17698), .C1(\registers[9][20] ), .C2(
        n17695), .A(n5863), .ZN(n5858) );
  OAI22_X1 U6749 ( .A1(n17692), .A2(n15778), .B1(n17689), .B2(n12191), .ZN(
        n5863) );
  AOI221_X1 U6750 ( .B1(net227289), .B2(n17698), .C1(\registers[9][21] ), .C2(
        n17695), .A(n5678), .ZN(n5671) );
  OAI22_X1 U6751 ( .A1(n17692), .A2(n15779), .B1(n17689), .B2(n12192), .ZN(
        n5678) );
  AOI221_X1 U6752 ( .B1(net227307), .B2(n17698), .C1(\registers[9][22] ), .C2(
        n17695), .A(n5492), .ZN(n5484) );
  OAI22_X1 U6753 ( .A1(n17692), .A2(n15780), .B1(n17689), .B2(n12193), .ZN(
        n5492) );
  AOI221_X1 U6754 ( .B1(net227469), .B2(n17697), .C1(\registers[9][31] ), .C2(
        n17694), .A(n14168), .ZN(n14154) );
  OAI22_X1 U6755 ( .A1(n17691), .A2(n15781), .B1(n17688), .B2(n12194), .ZN(
        n14168) );
  NOR3_X1 U6756 ( .A1(n13994), .A2(n12514), .A3(n13995), .ZN(n13993) );
  XNOR2_X1 U6757 ( .A(n13984), .B(N192), .ZN(n13994) );
  NOR3_X1 U6758 ( .A1(n12513), .A2(n12514), .A3(n12515), .ZN(n12512) );
  XNOR2_X1 U6759 ( .A(n12503), .B(N192), .ZN(n12513) );
  NOR3_X1 U6760 ( .A1(n14030), .A2(n14031), .A3(n17824), .ZN(n14029) );
  XNOR2_X1 U6761 ( .A(swp[1]), .B(n10189), .ZN(n14031) );
  XNOR2_X1 U6762 ( .A(swp[4]), .B(n14820), .ZN(n14030) );
  NOR2_X1 U6763 ( .A1(n10190), .A2(n10188), .ZN(n14016) );
  NOR2_X1 U6764 ( .A1(n13986), .A2(N46056), .ZN(n13904) );
  INV_X1 U6765 ( .A(n13987), .ZN(n13986) );
  NOR2_X1 U6766 ( .A1(n12505), .A2(N45542), .ZN(n12423) );
  INV_X1 U6767 ( .A(n12506), .ZN(n12505) );
  NOR2_X1 U6768 ( .A1(N46058), .A2(N46057), .ZN(n13985) );
  NOR2_X1 U6769 ( .A1(N45544), .A2(N45543), .ZN(n12504) );
  OAI22_X1 U6770 ( .A1(n17557), .A2(n16199), .B1(n16439), .B2(n17548), .ZN(
        n7797) );
  OAI22_X1 U6771 ( .A1(n17612), .A2(n16111), .B1(n16439), .B2(n17603), .ZN(
        n7799) );
  OAI22_X1 U6772 ( .A1(n16875), .A2(n15911), .B1(n16439), .B2(n16866), .ZN(
        n7805) );
  OAI22_X1 U6773 ( .A1(n17159), .A2(n15791), .B1(n16440), .B2(n17150), .ZN(
        n7817) );
  OAI22_X1 U6774 ( .A1(n17225), .A2(n15881), .B1(n16441), .B2(n17216), .ZN(
        n7820) );
  OAI22_X1 U6775 ( .A1(n17277), .A2(n15792), .B1(n16441), .B2(n17268), .ZN(
        n7822) );
  OAI22_X1 U6776 ( .A1(n17543), .A2(n16115), .B1(n16445), .B2(n17534), .ZN(
        n7834) );
  OAI22_X1 U6777 ( .A1(n17598), .A2(n16116), .B1(n16445), .B2(n17589), .ZN(
        n7873) );
  OAI22_X1 U6778 ( .A1(n16909), .A2(n15969), .B1(n16445), .B2(n16900), .ZN(
        n7881) );
  OAI22_X1 U6779 ( .A1(n16998), .A2(n15912), .B1(n16446), .B2(n16989), .ZN(
        n7885) );
  OAI22_X1 U6780 ( .A1(n17225), .A2(n15882), .B1(n16447), .B2(n17216), .ZN(
        n7894) );
  OAI22_X1 U6781 ( .A1(n17277), .A2(n15793), .B1(n16447), .B2(n17268), .ZN(
        n7896) );
  OAI22_X1 U6782 ( .A1(n17543), .A2(n16117), .B1(n16451), .B2(n17534), .ZN(
        n7908) );
  OAI22_X1 U6783 ( .A1(n17557), .A2(n16200), .B1(n16451), .B2(n17548), .ZN(
        n7909) );
  OAI22_X1 U6784 ( .A1(n17571), .A2(n16207), .B1(n16451), .B2(n17562), .ZN(
        n7910) );
  OAI22_X1 U6785 ( .A1(n16875), .A2(n15913), .B1(n16451), .B2(n16866), .ZN(
        n7954) );
  OAI22_X1 U6786 ( .A1(n17159), .A2(n15794), .B1(n16452), .B2(n17150), .ZN(
        n7966) );
  OAI22_X1 U6787 ( .A1(n17225), .A2(n15883), .B1(n16453), .B2(n17216), .ZN(
        n7968) );
  OAI22_X1 U6788 ( .A1(n17530), .A2(n15795), .B1(n17522), .B2(n16438), .ZN(
        n7796) );
  OAI22_X1 U6789 ( .A1(n17530), .A2(n15796), .B1(n17522), .B2(n16444), .ZN(
        n7871) );
  OAI22_X1 U6790 ( .A1(n17530), .A2(n15797), .B1(n17521), .B2(n16450), .ZN(
        n7947) );
  OAI22_X1 U6791 ( .A1(n17529), .A2(n15798), .B1(n17521), .B2(n16459), .ZN(
        n8029) );
  OAI22_X1 U6792 ( .A1(n17529), .A2(n15799), .B1(n17522), .B2(n16712), .ZN(
        n8157) );
  OAI22_X1 U6793 ( .A1(n17529), .A2(n15800), .B1(n17522), .B2(n16721), .ZN(
        n8229) );
  OAI22_X1 U6794 ( .A1(n17530), .A2(n15801), .B1(n17521), .B2(n16702), .ZN(
        n10125) );
  OAI22_X1 U6795 ( .A1(n17626), .A2(n16201), .B1(n17618), .B2(n16436), .ZN(
        n7763) );
  OAI22_X1 U6796 ( .A1(n17998), .A2(n15998), .B1(n17990), .B2(n16436), .ZN(
        n7768) );
  OAI22_X1 U6797 ( .A1(n17626), .A2(n16202), .B1(n17618), .B2(n16442), .ZN(
        n7838) );
  OAI22_X1 U6798 ( .A1(n17998), .A2(n15999), .B1(n17990), .B2(n16442), .ZN(
        n7843) );
  OAI22_X1 U6799 ( .A1(n17626), .A2(n16203), .B1(n17618), .B2(n16448), .ZN(
        n7914) );
  OAI22_X1 U6800 ( .A1(n17998), .A2(n16000), .B1(n17990), .B2(n16448), .ZN(
        n7919) );
  OAI22_X1 U6801 ( .A1(n17626), .A2(n16204), .B1(n17618), .B2(n16456), .ZN(
        n7988) );
  OAI22_X1 U6802 ( .A1(n17625), .A2(n16124), .B1(n17618), .B2(n16709), .ZN(
        n8116) );
  OAI22_X1 U6803 ( .A1(n17625), .A2(n16125), .B1(n17618), .B2(n16718), .ZN(
        n8188) );
  OAI22_X1 U6804 ( .A1(n17998), .A2(n16001), .B1(n17990), .B2(n16725), .ZN(
        n8269) );
  OAI22_X1 U6805 ( .A1(n17997), .A2(n16002), .B1(n17990), .B2(n16732), .ZN(
        n8341) );
  OAI22_X1 U6806 ( .A1(n17997), .A2(n16003), .B1(n17990), .B2(n16744), .ZN(
        n8485) );
  OAI22_X1 U6807 ( .A1(n17529), .A2(n15802), .B1(n17522), .B2(n16730), .ZN(
        n8325) );
  OAI22_X1 U6808 ( .A1(n16875), .A2(n15914), .B1(n16867), .B2(n16442), .ZN(
        n7844) );
  OAI22_X1 U6809 ( .A1(n16874), .A2(n15915), .B1(n16867), .B2(n16456), .ZN(
        n7992) );
  OAI22_X1 U6810 ( .A1(n16874), .A2(n15916), .B1(n16867), .B2(n16725), .ZN(
        n8272) );
  OAI22_X1 U6811 ( .A1(n16874), .A2(n15917), .B1(n16867), .B2(n16732), .ZN(
        n8344) );
  OAI22_X1 U6812 ( .A1(n16874), .A2(n15918), .B1(n16867), .B2(n16738), .ZN(
        n8416) );
  OAI22_X1 U6813 ( .A1(n16873), .A2(n15919), .B1(n16867), .B2(n16744), .ZN(
        n8488) );
  OAI22_X1 U6814 ( .A1(n16875), .A2(n15920), .B1(n16867), .B2(n16706), .ZN(
        n10072) );
  OAI22_X1 U6815 ( .A1(n16909), .A2(n15970), .B1(n16901), .B2(n16436), .ZN(
        n7771) );
  OAI22_X1 U6816 ( .A1(n16998), .A2(n15921), .B1(n16990), .B2(n16437), .ZN(
        n7775) );
  OAI22_X1 U6817 ( .A1(n17159), .A2(n15803), .B1(n17151), .B2(n16443), .ZN(
        n7856) );
  OAI22_X1 U6818 ( .A1(n16909), .A2(n15971), .B1(n16901), .B2(n16448), .ZN(
        n7921) );
  OAI22_X1 U6819 ( .A1(n16998), .A2(n15922), .B1(n16990), .B2(n16449), .ZN(
        n7925) );
  OAI22_X1 U6820 ( .A1(n17277), .A2(n15804), .B1(n17269), .B2(n16450), .ZN(
        n7936) );
  OAI22_X1 U6821 ( .A1(n16908), .A2(n15972), .B1(n16901), .B2(n16457), .ZN(
        n7995) );
  OAI22_X1 U6822 ( .A1(n17224), .A2(n15884), .B1(n17217), .B2(n16458), .ZN(
        n8006) );
  OAI22_X1 U6823 ( .A1(n17276), .A2(n15805), .B1(n17269), .B2(n16458), .ZN(
        n8010) );
  OAI22_X1 U6824 ( .A1(n16997), .A2(n15923), .B1(n16990), .B2(n16710), .ZN(
        n8123) );
  OAI22_X1 U6825 ( .A1(n17158), .A2(n15806), .B1(n17151), .B2(n16718), .ZN(
        n8200) );
  OAI22_X1 U6826 ( .A1(n17224), .A2(n15885), .B1(n17217), .B2(n16719), .ZN(
        n8206) );
  OAI22_X1 U6827 ( .A1(n17276), .A2(n15807), .B1(n17269), .B2(n16719), .ZN(
        n8210) );
  OAI22_X1 U6828 ( .A1(n16908), .A2(n15973), .B1(n16901), .B2(n16726), .ZN(
        n8275) );
  OAI22_X1 U6829 ( .A1(n16997), .A2(n15924), .B1(n16990), .B2(n16726), .ZN(
        n8283) );
  OAI22_X1 U6830 ( .A1(n17158), .A2(n15808), .B1(n17151), .B2(n16727), .ZN(
        n8296) );
  OAI22_X1 U6831 ( .A1(n17224), .A2(n15886), .B1(n17217), .B2(n16728), .ZN(
        n8302) );
  OAI22_X1 U6832 ( .A1(n17276), .A2(n15809), .B1(n17269), .B2(n16728), .ZN(
        n8306) );
  OAI22_X1 U6833 ( .A1(n16908), .A2(n15974), .B1(n16901), .B2(n16732), .ZN(
        n8347) );
  OAI22_X1 U6834 ( .A1(n16997), .A2(n15925), .B1(n16990), .B2(n16733), .ZN(
        n8355) );
  OAI22_X1 U6835 ( .A1(n17158), .A2(n15810), .B1(n17151), .B2(n16734), .ZN(
        n8368) );
  OAI22_X1 U6836 ( .A1(n17224), .A2(n15887), .B1(n17217), .B2(n16735), .ZN(
        n8374) );
  OAI22_X1 U6837 ( .A1(n17276), .A2(n15811), .B1(n17269), .B2(n16735), .ZN(
        n8378) );
  OAI22_X1 U6838 ( .A1(n17158), .A2(n15812), .B1(n17151), .B2(n16740), .ZN(
        n8440) );
  OAI22_X1 U6839 ( .A1(n17223), .A2(n15888), .B1(n17217), .B2(n16741), .ZN(
        n8446) );
  OAI22_X1 U6840 ( .A1(n16909), .A2(n15975), .B1(n16901), .B2(n16706), .ZN(
        n10075) );
  OAI22_X1 U6841 ( .A1(n16998), .A2(n15926), .B1(n16990), .B2(n16706), .ZN(
        n10083) );
  OAI22_X1 U6842 ( .A1(n17159), .A2(n15813), .B1(n17151), .B2(n16704), .ZN(
        n10096) );
  OAI22_X1 U6843 ( .A1(n17225), .A2(n15889), .B1(n17217), .B2(n16704), .ZN(
        n10102) );
  OAI22_X1 U6844 ( .A1(n17277), .A2(n15814), .B1(n17269), .B2(n16704), .ZN(
        n10106) );
  OAI22_X1 U6845 ( .A1(n17543), .A2(n16118), .B1(n17535), .B2(n16436), .ZN(
        n7760) );
  OAI22_X1 U6846 ( .A1(n17542), .A2(n16119), .B1(n17535), .B2(n16456), .ZN(
        n7982) );
  OAI22_X1 U6847 ( .A1(n17542), .A2(n16036), .B1(n17535), .B2(n16709), .ZN(
        n8110) );
  OAI22_X1 U6848 ( .A1(n17542), .A2(n16037), .B1(n17535), .B2(n16718), .ZN(
        n8182) );
  OAI22_X1 U6849 ( .A1(n17542), .A2(n16038), .B1(n17535), .B2(n16731), .ZN(
        n8326) );
  OAI22_X1 U6850 ( .A1(n17541), .A2(n16039), .B1(n17535), .B2(n16737), .ZN(
        n8398) );
  OAI22_X1 U6851 ( .A1(n17571), .A2(n16208), .B1(n17563), .B2(n16436), .ZN(
        n7761) );
  OAI22_X1 U6852 ( .A1(n17598), .A2(n16120), .B1(n17590), .B2(n16436), .ZN(
        n7762) );
  OAI22_X1 U6853 ( .A1(n17557), .A2(n16205), .B1(n17549), .B2(n16442), .ZN(
        n7835) );
  OAI22_X1 U6854 ( .A1(n17571), .A2(n16209), .B1(n17563), .B2(n16442), .ZN(
        n7836) );
  OAI22_X1 U6855 ( .A1(n17612), .A2(n16112), .B1(n17604), .B2(n16442), .ZN(
        n7837) );
  OAI22_X1 U6856 ( .A1(n17598), .A2(n16121), .B1(n17590), .B2(n16448), .ZN(
        n7912) );
  OAI22_X1 U6857 ( .A1(n17612), .A2(n16113), .B1(n17604), .B2(n16448), .ZN(
        n7913) );
  OAI22_X1 U6858 ( .A1(n17557), .A2(n16206), .B1(n17549), .B2(n16456), .ZN(
        n7983) );
  OAI22_X1 U6859 ( .A1(n17571), .A2(n16210), .B1(n17563), .B2(n16456), .ZN(
        n7984) );
  OAI22_X1 U6860 ( .A1(n17598), .A2(n16122), .B1(n17590), .B2(n16456), .ZN(
        n7986) );
  OAI22_X1 U6861 ( .A1(n17612), .A2(n16114), .B1(n17604), .B2(n16456), .ZN(
        n7987) );
  OAI22_X1 U6862 ( .A1(n17556), .A2(n16126), .B1(n17549), .B2(n16709), .ZN(
        n8111) );
  OAI22_X1 U6863 ( .A1(n17570), .A2(n16174), .B1(n17563), .B2(n16709), .ZN(
        n8112) );
  OAI22_X1 U6864 ( .A1(n17597), .A2(n16040), .B1(n17590), .B2(n16709), .ZN(
        n8114) );
  OAI22_X1 U6865 ( .A1(n17611), .A2(n16086), .B1(n17604), .B2(n16709), .ZN(
        n8115) );
  OAI22_X1 U6866 ( .A1(n17556), .A2(n16127), .B1(n17549), .B2(n16718), .ZN(
        n8183) );
  OAI22_X1 U6867 ( .A1(n17570), .A2(n16175), .B1(n17563), .B2(n16718), .ZN(
        n8184) );
  OAI22_X1 U6868 ( .A1(n17597), .A2(n16041), .B1(n17590), .B2(n16718), .ZN(
        n8186) );
  OAI22_X1 U6869 ( .A1(n17611), .A2(n16087), .B1(n17604), .B2(n16718), .ZN(
        n8187) );
  OAI22_X1 U6870 ( .A1(n17556), .A2(n16128), .B1(n17549), .B2(n16731), .ZN(
        n8327) );
  OAI22_X1 U6871 ( .A1(n16908), .A2(n15976), .B1(n16901), .B2(n16738), .ZN(
        n8419) );
  OAI22_X1 U6872 ( .A1(n16997), .A2(n15927), .B1(n16990), .B2(n16739), .ZN(
        n8427) );
  OAI22_X1 U6873 ( .A1(n17275), .A2(n15815), .B1(n17269), .B2(n16741), .ZN(
        n8450) );
  OAI22_X1 U6874 ( .A1(n16907), .A2(n15977), .B1(n16901), .B2(n16744), .ZN(
        n8491) );
  OAI22_X1 U6875 ( .A1(n16996), .A2(n15928), .B1(n16990), .B2(n16745), .ZN(
        n8499) );
  OAI22_X1 U6876 ( .A1(n17157), .A2(n15816), .B1(n17151), .B2(n16746), .ZN(
        n8512) );
  OAI22_X1 U6877 ( .A1(n17223), .A2(n15890), .B1(n17217), .B2(n16747), .ZN(
        n8518) );
  OAI22_X1 U6878 ( .A1(n17275), .A2(n15817), .B1(n17269), .B2(n16747), .ZN(
        n8522) );
  OAI22_X1 U6879 ( .A1(n16907), .A2(n15978), .B1(n16901), .B2(n16750), .ZN(
        n8563) );
  OAI22_X1 U6880 ( .A1(n16996), .A2(n15929), .B1(n16990), .B2(n16751), .ZN(
        n8571) );
  OAI22_X1 U6881 ( .A1(n17157), .A2(n15818), .B1(n17151), .B2(n16752), .ZN(
        n8584) );
  OAI22_X1 U6882 ( .A1(n17223), .A2(n15891), .B1(n17217), .B2(n16753), .ZN(
        n8590) );
  OAI22_X1 U6883 ( .A1(n17275), .A2(n15819), .B1(n17269), .B2(n16753), .ZN(
        n8594) );
  OAI22_X1 U6884 ( .A1(n16907), .A2(n15979), .B1(n16901), .B2(n16756), .ZN(
        n8635) );
  OAI22_X1 U6885 ( .A1(n16996), .A2(n15930), .B1(n16990), .B2(n16757), .ZN(
        n8643) );
  OAI22_X1 U6886 ( .A1(n17157), .A2(n15820), .B1(n17151), .B2(n16758), .ZN(
        n8656) );
  OAI22_X1 U6887 ( .A1(n17223), .A2(n15892), .B1(n17217), .B2(n16759), .ZN(
        n8662) );
  OAI22_X1 U6888 ( .A1(n17275), .A2(n15821), .B1(n17269), .B2(n16759), .ZN(
        n8666) );
  OAI22_X1 U6889 ( .A1(n16907), .A2(n15980), .B1(n16901), .B2(n16762), .ZN(
        n8707) );
  OAI22_X1 U6890 ( .A1(n16996), .A2(n15931), .B1(n16990), .B2(n16763), .ZN(
        n8715) );
  OAI22_X1 U6891 ( .A1(n17157), .A2(n15822), .B1(n17151), .B2(n16764), .ZN(
        n8728) );
  OAI22_X1 U6892 ( .A1(n17222), .A2(n15893), .B1(n17217), .B2(n16765), .ZN(
        n8734) );
  OAI22_X1 U6893 ( .A1(n17274), .A2(n15823), .B1(n17269), .B2(n16765), .ZN(
        n8738) );
  OAI22_X1 U6894 ( .A1(n16906), .A2(n15981), .B1(n16901), .B2(n16768), .ZN(
        n8779) );
  OAI22_X1 U6895 ( .A1(n16995), .A2(n15932), .B1(n16990), .B2(n16769), .ZN(
        n8787) );
  OAI22_X1 U6896 ( .A1(n17156), .A2(n15824), .B1(n17151), .B2(n16770), .ZN(
        n8800) );
  OAI22_X1 U6897 ( .A1(n17222), .A2(n15894), .B1(n17217), .B2(n16771), .ZN(
        n8806) );
  OAI22_X1 U6898 ( .A1(n17274), .A2(n15825), .B1(n17269), .B2(n16771), .ZN(
        n8810) );
  OAI22_X1 U6899 ( .A1(n16906), .A2(n15982), .B1(n16901), .B2(n16774), .ZN(
        n8851) );
  OAI22_X1 U6900 ( .A1(n16995), .A2(n15933), .B1(n16990), .B2(n16775), .ZN(
        n8859) );
  OAI22_X1 U6901 ( .A1(n17156), .A2(n15826), .B1(n17151), .B2(n16776), .ZN(
        n8872) );
  OAI22_X1 U6902 ( .A1(n17222), .A2(n15895), .B1(n17217), .B2(n16777), .ZN(
        n8878) );
  OAI22_X1 U6903 ( .A1(n17274), .A2(n15827), .B1(n17269), .B2(n16777), .ZN(
        n8882) );
  OAI22_X1 U6904 ( .A1(n16906), .A2(n15983), .B1(n16901), .B2(n16780), .ZN(
        n8923) );
  OAI22_X1 U6905 ( .A1(n16995), .A2(n15934), .B1(n16990), .B2(n16781), .ZN(
        n8931) );
  OAI22_X1 U6906 ( .A1(n17156), .A2(n15828), .B1(n17151), .B2(n16782), .ZN(
        n8944) );
  OAI22_X1 U6907 ( .A1(n17221), .A2(n15896), .B1(n17217), .B2(n16783), .ZN(
        n8950) );
  OAI22_X1 U6908 ( .A1(n17273), .A2(n15829), .B1(n17269), .B2(n16783), .ZN(
        n8954) );
  OAI22_X1 U6909 ( .A1(n16905), .A2(n15984), .B1(n16901), .B2(n16786), .ZN(
        n8995) );
  OAI22_X1 U6910 ( .A1(n16994), .A2(n15935), .B1(n16990), .B2(n16787), .ZN(
        n9003) );
  OAI22_X1 U6911 ( .A1(n17155), .A2(n15830), .B1(n17151), .B2(n16788), .ZN(
        n9016) );
  OAI22_X1 U6912 ( .A1(n17221), .A2(n15897), .B1(n17217), .B2(n16789), .ZN(
        n9022) );
  OAI22_X1 U6913 ( .A1(n17273), .A2(n15831), .B1(n17269), .B2(n16789), .ZN(
        n9026) );
  OAI22_X1 U6914 ( .A1(n16905), .A2(n15985), .B1(n16901), .B2(n16792), .ZN(
        n9067) );
  OAI22_X1 U6915 ( .A1(n16994), .A2(n15936), .B1(n16990), .B2(n16793), .ZN(
        n9075) );
  OAI22_X1 U6916 ( .A1(n17155), .A2(n15832), .B1(n17151), .B2(n16794), .ZN(
        n9088) );
  OAI22_X1 U6917 ( .A1(n17221), .A2(n15898), .B1(n17217), .B2(n16795), .ZN(
        n9094) );
  OAI22_X1 U6918 ( .A1(n17273), .A2(n15833), .B1(n17269), .B2(n16795), .ZN(
        n9098) );
  OAI22_X1 U6919 ( .A1(n16905), .A2(n15986), .B1(n16901), .B2(n16798), .ZN(
        n9139) );
  OAI22_X1 U6920 ( .A1(n16994), .A2(n15937), .B1(n16990), .B2(n16799), .ZN(
        n9147) );
  OAI22_X1 U6921 ( .A1(n17155), .A2(n15834), .B1(n17151), .B2(n16800), .ZN(
        n9160) );
  OAI22_X1 U6922 ( .A1(n17221), .A2(n15899), .B1(n17217), .B2(n16801), .ZN(
        n9166) );
  OAI22_X1 U6923 ( .A1(n17273), .A2(n15835), .B1(n17269), .B2(n16801), .ZN(
        n9170) );
  OAI22_X1 U6924 ( .A1(n16905), .A2(n15987), .B1(n16901), .B2(n16804), .ZN(
        n9211) );
  OAI22_X1 U6925 ( .A1(n16994), .A2(n15938), .B1(n16990), .B2(n16805), .ZN(
        n9219) );
  OAI22_X1 U6926 ( .A1(n17155), .A2(n15836), .B1(n17151), .B2(n16806), .ZN(
        n9232) );
  OAI22_X1 U6927 ( .A1(n17220), .A2(n15900), .B1(n17217), .B2(n16807), .ZN(
        n9238) );
  OAI22_X1 U6928 ( .A1(n17272), .A2(n15837), .B1(n17269), .B2(n16807), .ZN(
        n9242) );
  OAI22_X1 U6929 ( .A1(n17154), .A2(n15838), .B1(n17151), .B2(n16812), .ZN(
        n9304) );
  OAI22_X1 U6930 ( .A1(n17220), .A2(n15901), .B1(n17217), .B2(n16813), .ZN(
        n9310) );
  OAI22_X1 U6931 ( .A1(n16906), .A2(n15988), .B1(n16901), .B2(n17513), .ZN(
        n9931) );
  OAI22_X1 U6932 ( .A1(n16995), .A2(n15939), .B1(n16990), .B2(n17514), .ZN(
        n9939) );
  OAI22_X1 U6933 ( .A1(n17156), .A2(n15839), .B1(n17151), .B2(n17515), .ZN(
        n9952) );
  OAI22_X1 U6934 ( .A1(n17222), .A2(n15902), .B1(n17217), .B2(n17516), .ZN(
        n9958) );
  OAI22_X1 U6935 ( .A1(n17274), .A2(n15840), .B1(n17269), .B2(n17516), .ZN(
        n9962) );
  NAND2_X1 U6936 ( .A1(N192), .A2(n14223), .ZN(n12413) );
  OAI22_X1 U6937 ( .A1(net227474), .A2(n14007), .B1(n14009), .B2(n14012), .ZN(
        n10136) );
  XNOR2_X1 U6938 ( .A(N9641), .B(n10189), .ZN(n14012) );
  OAI22_X1 U6939 ( .A1(net227475), .A2(n14007), .B1(n14009), .B2(n14010), .ZN(
        n10137) );
  OAI22_X1 U6940 ( .A1(n17220), .A2(n15903), .B1(n17216), .B2(n16819), .ZN(
        n9382) );
  OAI22_X1 U6941 ( .A1(n17220), .A2(n15904), .B1(n17216), .B2(n16825), .ZN(
        n9454) );
  OAI22_X1 U6942 ( .A1(n17219), .A2(n15905), .B1(n17216), .B2(n16831), .ZN(
        n9526) );
  OAI22_X1 U6943 ( .A1(n17219), .A2(n15906), .B1(n17216), .B2(n16837), .ZN(
        n9598) );
  OAI22_X1 U6944 ( .A1(n17219), .A2(n15907), .B1(n17216), .B2(n16843), .ZN(
        n9670) );
  OAI22_X1 U6945 ( .A1(n17219), .A2(n15908), .B1(n17216), .B2(n16849), .ZN(
        n9742) );
  OAI22_X1 U6946 ( .A1(n17218), .A2(n15909), .B1(n17216), .B2(n16855), .ZN(
        n9814) );
  OAI22_X1 U6947 ( .A1(n17218), .A2(n15910), .B1(n17216), .B2(n16861), .ZN(
        n9886) );
  OAI22_X1 U6948 ( .A1(n17154), .A2(n15841), .B1(n17150), .B2(n16818), .ZN(
        n9376) );
  OAI22_X1 U6949 ( .A1(n17154), .A2(n15842), .B1(n17150), .B2(n16824), .ZN(
        n9448) );
  OAI22_X1 U6950 ( .A1(n17153), .A2(n15843), .B1(n17150), .B2(n16830), .ZN(
        n9520) );
  OAI22_X1 U6951 ( .A1(n17154), .A2(n15844), .B1(n17150), .B2(n16836), .ZN(
        n9592) );
  OAI22_X1 U6952 ( .A1(n17153), .A2(n15845), .B1(n17150), .B2(n16842), .ZN(
        n9664) );
  OAI22_X1 U6953 ( .A1(n17153), .A2(n15846), .B1(n17150), .B2(n16848), .ZN(
        n9736) );
  OAI22_X1 U6954 ( .A1(n17153), .A2(n15847), .B1(n17150), .B2(n16854), .ZN(
        n9808) );
  OAI22_X1 U6955 ( .A1(n17152), .A2(n15848), .B1(n17150), .B2(n16860), .ZN(
        n9880) );
  OAI22_X1 U6956 ( .A1(n17272), .A2(n15849), .B1(n17268), .B2(n16813), .ZN(
        n9314) );
  OAI22_X1 U6957 ( .A1(n17272), .A2(n15850), .B1(n17268), .B2(n16819), .ZN(
        n9386) );
  OAI22_X1 U6958 ( .A1(n16870), .A2(n15940), .B1(n16866), .B2(n16822), .ZN(
        n9424) );
  OAI22_X1 U6959 ( .A1(n17272), .A2(n15851), .B1(n17268), .B2(n16825), .ZN(
        n9458) );
  OAI22_X1 U6960 ( .A1(n16870), .A2(n15941), .B1(n16866), .B2(n16828), .ZN(
        n9496) );
  OAI22_X1 U6961 ( .A1(n17271), .A2(n15852), .B1(n17268), .B2(n16831), .ZN(
        n9530) );
  OAI22_X1 U6962 ( .A1(n16869), .A2(n15942), .B1(n16866), .B2(n16834), .ZN(
        n9568) );
  OAI22_X1 U6963 ( .A1(n17271), .A2(n15853), .B1(n17268), .B2(n16837), .ZN(
        n9602) );
  OAI22_X1 U6964 ( .A1(n16869), .A2(n15943), .B1(n16866), .B2(n16840), .ZN(
        n9640) );
  OAI22_X1 U6965 ( .A1(n17271), .A2(n15854), .B1(n17268), .B2(n16843), .ZN(
        n9674) );
  OAI22_X1 U6966 ( .A1(n16869), .A2(n15944), .B1(n16866), .B2(n16846), .ZN(
        n9712) );
  OAI22_X1 U6967 ( .A1(n17271), .A2(n15855), .B1(n17268), .B2(n16849), .ZN(
        n9746) );
  OAI22_X1 U6968 ( .A1(n16869), .A2(n15945), .B1(n16866), .B2(n16852), .ZN(
        n9784) );
  OAI22_X1 U6969 ( .A1(n17270), .A2(n15856), .B1(n17268), .B2(n16855), .ZN(
        n9818) );
  OAI22_X1 U6970 ( .A1(n16868), .A2(n15946), .B1(n16866), .B2(n16858), .ZN(
        n9856) );
  OAI22_X1 U6971 ( .A1(n17270), .A2(n15857), .B1(n17268), .B2(n16861), .ZN(
        n9890) );
  OAI22_X1 U6972 ( .A1(n15782), .A2(n16868), .B1(n16866), .B2(n18031), .ZN(
        n10000) );
  OAI22_X1 U6973 ( .A1(n17552), .A2(n16129), .B1(n17548), .B2(n16809), .ZN(
        n9263) );
  OAI22_X1 U6974 ( .A1(n17538), .A2(n16042), .B1(n17534), .B2(n16815), .ZN(
        n9334) );
  OAI22_X1 U6975 ( .A1(n17552), .A2(n16130), .B1(n17548), .B2(n16815), .ZN(
        n9335) );
  OAI22_X1 U6976 ( .A1(n17537), .A2(n16043), .B1(n17534), .B2(n16827), .ZN(
        n9478) );
  OAI22_X1 U6977 ( .A1(n17552), .A2(n16131), .B1(n17548), .B2(n16827), .ZN(
        n9479) );
  OAI22_X1 U6978 ( .A1(n17537), .A2(n16044), .B1(n17534), .B2(n16833), .ZN(
        n9550) );
  OAI22_X1 U6979 ( .A1(n17551), .A2(n16132), .B1(n17548), .B2(n16833), .ZN(
        n9551) );
  OAI22_X1 U6980 ( .A1(n17538), .A2(n16045), .B1(n17534), .B2(n16839), .ZN(
        n9622) );
  OAI22_X1 U6981 ( .A1(n17552), .A2(n16133), .B1(n17548), .B2(n16839), .ZN(
        n9623) );
  OAI22_X1 U6982 ( .A1(n17537), .A2(n16046), .B1(n17534), .B2(n16845), .ZN(
        n9694) );
  OAI22_X1 U6983 ( .A1(n17551), .A2(n16134), .B1(n17548), .B2(n16845), .ZN(
        n9695) );
  OAI22_X1 U6984 ( .A1(n17536), .A2(n16047), .B1(n17534), .B2(n16851), .ZN(
        n9766) );
  OAI22_X1 U6985 ( .A1(n17551), .A2(n16135), .B1(n17548), .B2(n16851), .ZN(
        n9767) );
  OAI22_X1 U6986 ( .A1(n17537), .A2(n16048), .B1(n17534), .B2(n16857), .ZN(
        n9838) );
  OAI22_X1 U6987 ( .A1(n17551), .A2(n16136), .B1(n17548), .B2(n16857), .ZN(
        n9839) );
  OAI22_X1 U6988 ( .A1(n17536), .A2(n16049), .B1(n17534), .B2(n17512), .ZN(
        n9910) );
  OAI22_X1 U6989 ( .A1(n17550), .A2(n16137), .B1(n17548), .B2(n17512), .ZN(
        n9911) );
  OAI22_X1 U6990 ( .A1(n17543), .A2(n16123), .B1(n17534), .B2(n16702), .ZN(
        n10054) );
  OAI22_X1 U6991 ( .A1(n16904), .A2(n15989), .B1(n16900), .B2(n16810), .ZN(
        n9283) );
  OAI22_X1 U6992 ( .A1(n16993), .A2(n15947), .B1(n16989), .B2(n16811), .ZN(
        n9291) );
  OAI22_X1 U6993 ( .A1(n16904), .A2(n15990), .B1(n16900), .B2(n16816), .ZN(
        n9355) );
  OAI22_X1 U6994 ( .A1(n16993), .A2(n15948), .B1(n16989), .B2(n16817), .ZN(
        n9363) );
  OAI22_X1 U6995 ( .A1(n16904), .A2(n15991), .B1(n16900), .B2(n16822), .ZN(
        n9427) );
  OAI22_X1 U6996 ( .A1(n16993), .A2(n15949), .B1(n16989), .B2(n16823), .ZN(
        n9435) );
  OAI22_X1 U6997 ( .A1(n16904), .A2(n15992), .B1(n16900), .B2(n16828), .ZN(
        n9499) );
  OAI22_X1 U6998 ( .A1(n16992), .A2(n15950), .B1(n16989), .B2(n16829), .ZN(
        n9507) );
  OAI22_X1 U6999 ( .A1(n16903), .A2(n15993), .B1(n16900), .B2(n16834), .ZN(
        n9571) );
  OAI22_X1 U7000 ( .A1(n16993), .A2(n15951), .B1(n16989), .B2(n16835), .ZN(
        n9579) );
  OAI22_X1 U7001 ( .A1(n16903), .A2(n15994), .B1(n16900), .B2(n16840), .ZN(
        n9643) );
  OAI22_X1 U7002 ( .A1(n16992), .A2(n15952), .B1(n16989), .B2(n16841), .ZN(
        n9651) );
  OAI22_X1 U7003 ( .A1(n16903), .A2(n15995), .B1(n16900), .B2(n16846), .ZN(
        n9715) );
  OAI22_X1 U7004 ( .A1(n16992), .A2(n15953), .B1(n16989), .B2(n16847), .ZN(
        n9723) );
  OAI22_X1 U7005 ( .A1(n16903), .A2(n15996), .B1(n16900), .B2(n16852), .ZN(
        n9787) );
  OAI22_X1 U7006 ( .A1(n16992), .A2(n15954), .B1(n16989), .B2(n16853), .ZN(
        n9795) );
  OAI22_X1 U7007 ( .A1(n16902), .A2(n15997), .B1(n16900), .B2(n16858), .ZN(
        n9859) );
  OAI22_X1 U7008 ( .A1(n16991), .A2(n15955), .B1(n16989), .B2(n16859), .ZN(
        n9867) );
  OAI22_X1 U7009 ( .A1(n17567), .A2(n16176), .B1(n17562), .B2(n16803), .ZN(
        n9192) );
  OAI22_X1 U7010 ( .A1(n17594), .A2(n16050), .B1(n17589), .B2(n16803), .ZN(
        n9194) );
  OAI22_X1 U7011 ( .A1(n17608), .A2(n16088), .B1(n17603), .B2(n16803), .ZN(
        n9195) );
  OAI22_X1 U7012 ( .A1(n17566), .A2(n16177), .B1(n17562), .B2(n16809), .ZN(
        n9264) );
  OAI22_X1 U7013 ( .A1(n17593), .A2(n16051), .B1(n17589), .B2(n16809), .ZN(
        n9266) );
  OAI22_X1 U7014 ( .A1(n17607), .A2(n16089), .B1(n17603), .B2(n16809), .ZN(
        n9267) );
  OAI22_X1 U7015 ( .A1(n17566), .A2(n16178), .B1(n17562), .B2(n16815), .ZN(
        n9336) );
  OAI22_X1 U7016 ( .A1(n17593), .A2(n16052), .B1(n17589), .B2(n16815), .ZN(
        n9338) );
  OAI22_X1 U7017 ( .A1(n17607), .A2(n16090), .B1(n17603), .B2(n16815), .ZN(
        n9339) );
  OAI22_X1 U7018 ( .A1(n17566), .A2(n16179), .B1(n17562), .B2(n16827), .ZN(
        n9480) );
  OAI22_X1 U7019 ( .A1(n17593), .A2(n16053), .B1(n17589), .B2(n16827), .ZN(
        n9482) );
  OAI22_X1 U7020 ( .A1(n17607), .A2(n16091), .B1(n17603), .B2(n16827), .ZN(
        n9483) );
  OAI22_X1 U7021 ( .A1(n17565), .A2(n16180), .B1(n17562), .B2(n16833), .ZN(
        n9552) );
  OAI22_X1 U7022 ( .A1(n17592), .A2(n16054), .B1(n17589), .B2(n16833), .ZN(
        n9554) );
  OAI22_X1 U7023 ( .A1(n17606), .A2(n16092), .B1(n17603), .B2(n16833), .ZN(
        n9555) );
  OAI22_X1 U7024 ( .A1(n17566), .A2(n16181), .B1(n17562), .B2(n16839), .ZN(
        n9624) );
  OAI22_X1 U7025 ( .A1(n17593), .A2(n16055), .B1(n17589), .B2(n16839), .ZN(
        n9626) );
  OAI22_X1 U7026 ( .A1(n17607), .A2(n16093), .B1(n17603), .B2(n16839), .ZN(
        n9627) );
  OAI22_X1 U7027 ( .A1(n17565), .A2(n16182), .B1(n17562), .B2(n16845), .ZN(
        n9696) );
  OAI22_X1 U7028 ( .A1(n17592), .A2(n16056), .B1(n17589), .B2(n16845), .ZN(
        n9698) );
  OAI22_X1 U7029 ( .A1(n17606), .A2(n16094), .B1(n17603), .B2(n16845), .ZN(
        n9699) );
  OAI22_X1 U7030 ( .A1(n17565), .A2(n16183), .B1(n17562), .B2(n16851), .ZN(
        n9768) );
  OAI22_X1 U7031 ( .A1(n17592), .A2(n16057), .B1(n17589), .B2(n16851), .ZN(
        n9770) );
  OAI22_X1 U7032 ( .A1(n17606), .A2(n16095), .B1(n17603), .B2(n16851), .ZN(
        n9771) );
  OAI22_X1 U7033 ( .A1(n17565), .A2(n16184), .B1(n17562), .B2(n16857), .ZN(
        n9840) );
  OAI22_X1 U7034 ( .A1(n17592), .A2(n16058), .B1(n17589), .B2(n16857), .ZN(
        n9842) );
  OAI22_X1 U7035 ( .A1(n17606), .A2(n16096), .B1(n17603), .B2(n16857), .ZN(
        n9843) );
  OAI22_X1 U7036 ( .A1(n17564), .A2(n16185), .B1(n17562), .B2(n17512), .ZN(
        n9912) );
  OAI22_X1 U7037 ( .A1(n17591), .A2(n16059), .B1(n17589), .B2(n17512), .ZN(
        n9914) );
  OAI22_X1 U7038 ( .A1(n17605), .A2(n16097), .B1(n17603), .B2(n17512), .ZN(
        n9915) );
  OAI22_X1 U7039 ( .A1(n17994), .A2(n16004), .B1(n17989), .B2(n16810), .ZN(
        n9277) );
  OAI22_X1 U7040 ( .A1(n17994), .A2(n16005), .B1(n17989), .B2(n16816), .ZN(
        n9349) );
  OAI22_X1 U7041 ( .A1(n17993), .A2(n16006), .B1(n17989), .B2(n16828), .ZN(
        n9493) );
  OAI22_X1 U7042 ( .A1(n17993), .A2(n16007), .B1(n17989), .B2(n16834), .ZN(
        n9565) );
  OAI22_X1 U7043 ( .A1(n17993), .A2(n16008), .B1(n17989), .B2(n16840), .ZN(
        n9637) );
  OAI22_X1 U7044 ( .A1(n17992), .A2(n16009), .B1(n17989), .B2(n16846), .ZN(
        n9709) );
  OAI22_X1 U7045 ( .A1(n17992), .A2(n16010), .B1(n17989), .B2(n16852), .ZN(
        n9781) );
  OAI22_X1 U7046 ( .A1(n17992), .A2(n16011), .B1(n17989), .B2(n16858), .ZN(
        n9853) );
  OAI22_X1 U7047 ( .A1(n17993), .A2(n16012), .B1(n17989), .B2(n17513), .ZN(
        n9925) );
  OAI22_X1 U7048 ( .A1(n17528), .A2(n15858), .B1(n17522), .B2(n16736), .ZN(
        n8397) );
  OAI22_X1 U7049 ( .A1(n17528), .A2(n15859), .B1(n17522), .B2(n16742), .ZN(
        n8469) );
  OAI22_X1 U7050 ( .A1(n17528), .A2(n15860), .B1(n17522), .B2(n16748), .ZN(
        n8541) );
  OAI22_X1 U7051 ( .A1(n17528), .A2(n15861), .B1(n17522), .B2(n16754), .ZN(
        n8613) );
  OAI22_X1 U7052 ( .A1(n17527), .A2(n15862), .B1(n17522), .B2(n16760), .ZN(
        n8685) );
  OAI22_X1 U7053 ( .A1(n17527), .A2(n15863), .B1(n17522), .B2(n16766), .ZN(
        n8757) );
  OAI22_X1 U7054 ( .A1(n17527), .A2(n15864), .B1(n17522), .B2(n16772), .ZN(
        n8829) );
  OAI22_X1 U7055 ( .A1(n17526), .A2(n15865), .B1(n17522), .B2(n16778), .ZN(
        n8901) );
  OAI22_X1 U7056 ( .A1(n17526), .A2(n15866), .B1(n17522), .B2(n16784), .ZN(
        n8973) );
  OAI22_X1 U7057 ( .A1(n17526), .A2(n15867), .B1(n17522), .B2(n16790), .ZN(
        n9045) );
  OAI22_X1 U7058 ( .A1(n17526), .A2(n15868), .B1(n17522), .B2(n16796), .ZN(
        n9117) );
  OAI22_X1 U7059 ( .A1(n17525), .A2(n15869), .B1(n17521), .B2(n16802), .ZN(
        n9189) );
  OAI22_X1 U7060 ( .A1(n17525), .A2(n15870), .B1(n17521), .B2(n16808), .ZN(
        n9261) );
  OAI22_X1 U7061 ( .A1(n17525), .A2(n15871), .B1(n17521), .B2(n16814), .ZN(
        n9333) );
  OAI22_X1 U7062 ( .A1(n17525), .A2(n15872), .B1(n17521), .B2(n16820), .ZN(
        n9405) );
  OAI22_X1 U7063 ( .A1(n17524), .A2(n15873), .B1(n17521), .B2(n16826), .ZN(
        n9477) );
  OAI22_X1 U7064 ( .A1(n17524), .A2(n15874), .B1(n17521), .B2(n16832), .ZN(
        n9549) );
  OAI22_X1 U7065 ( .A1(n17524), .A2(n15875), .B1(n17521), .B2(n16838), .ZN(
        n9621) );
  OAI22_X1 U7066 ( .A1(n17524), .A2(n15876), .B1(n17521), .B2(n16844), .ZN(
        n9693) );
  OAI22_X1 U7067 ( .A1(n17523), .A2(n15877), .B1(n17521), .B2(n16850), .ZN(
        n9765) );
  OAI22_X1 U7068 ( .A1(n17523), .A2(n15878), .B1(n17521), .B2(n16856), .ZN(
        n9837) );
  OAI22_X1 U7069 ( .A1(n17523), .A2(n15879), .B1(n17521), .B2(n16862), .ZN(
        n9909) );
  OAI22_X1 U7070 ( .A1(n17527), .A2(n15880), .B1(n17521), .B2(n17517), .ZN(
        n9981) );
  OAI22_X1 U7071 ( .A1(n17622), .A2(n16138), .B1(n17617), .B2(n16797), .ZN(
        n9124) );
  OAI22_X1 U7072 ( .A1(n17622), .A2(n16139), .B1(n17617), .B2(n16803), .ZN(
        n9196) );
  OAI22_X1 U7073 ( .A1(n17621), .A2(n16140), .B1(n17617), .B2(n16809), .ZN(
        n9268) );
  OAI22_X1 U7074 ( .A1(n17621), .A2(n16141), .B1(n17617), .B2(n16815), .ZN(
        n9340) );
  OAI22_X1 U7075 ( .A1(n17621), .A2(n16142), .B1(n17617), .B2(n16827), .ZN(
        n9484) );
  OAI22_X1 U7076 ( .A1(n17620), .A2(n16143), .B1(n17617), .B2(n16833), .ZN(
        n9556) );
  OAI22_X1 U7077 ( .A1(n17621), .A2(n16144), .B1(n17617), .B2(n16839), .ZN(
        n9628) );
  OAI22_X1 U7078 ( .A1(n17620), .A2(n16145), .B1(n17617), .B2(n16845), .ZN(
        n9700) );
  OAI22_X1 U7079 ( .A1(n17620), .A2(n16146), .B1(n17617), .B2(n16851), .ZN(
        n9772) );
  OAI22_X1 U7080 ( .A1(n17620), .A2(n16147), .B1(n17617), .B2(n16857), .ZN(
        n9844) );
  OAI22_X1 U7081 ( .A1(n17619), .A2(n16148), .B1(n17617), .B2(n17512), .ZN(
        n9916) );
  OAI22_X1 U7082 ( .A1(n17625), .A2(n16149), .B1(n17618), .B2(n16731), .ZN(
        n8332) );
  OAI22_X1 U7083 ( .A1(n17625), .A2(n16150), .B1(n17618), .B2(n16737), .ZN(
        n8404) );
  OAI22_X1 U7084 ( .A1(n17997), .A2(n16013), .B1(n17990), .B2(n16738), .ZN(
        n8413) );
  OAI22_X1 U7085 ( .A1(n17624), .A2(n16151), .B1(n17618), .B2(n16743), .ZN(
        n8476) );
  OAI22_X1 U7086 ( .A1(n17624), .A2(n16152), .B1(n17618), .B2(n16749), .ZN(
        n8548) );
  OAI22_X1 U7087 ( .A1(n17997), .A2(n16014), .B1(n17990), .B2(n16750), .ZN(
        n8557) );
  OAI22_X1 U7088 ( .A1(n17624), .A2(n16153), .B1(n17618), .B2(n16755), .ZN(
        n8620) );
  OAI22_X1 U7089 ( .A1(n17996), .A2(n16015), .B1(n17990), .B2(n16756), .ZN(
        n8629) );
  OAI22_X1 U7090 ( .A1(n17624), .A2(n16154), .B1(n17618), .B2(n16761), .ZN(
        n8692) );
  OAI22_X1 U7091 ( .A1(n17996), .A2(n16016), .B1(n17990), .B2(n16762), .ZN(
        n8701) );
  OAI22_X1 U7092 ( .A1(n17623), .A2(n16155), .B1(n17618), .B2(n16767), .ZN(
        n8764) );
  OAI22_X1 U7093 ( .A1(n17996), .A2(n16017), .B1(n17990), .B2(n16768), .ZN(
        n8773) );
  OAI22_X1 U7094 ( .A1(n17623), .A2(n16156), .B1(n17618), .B2(n16773), .ZN(
        n8836) );
  OAI22_X1 U7095 ( .A1(n17996), .A2(n16018), .B1(n17990), .B2(n16774), .ZN(
        n8845) );
  OAI22_X1 U7096 ( .A1(n17623), .A2(n16157), .B1(n17618), .B2(n16779), .ZN(
        n8908) );
  OAI22_X1 U7097 ( .A1(n17995), .A2(n16019), .B1(n17990), .B2(n16780), .ZN(
        n8917) );
  OAI22_X1 U7098 ( .A1(n17622), .A2(n16158), .B1(n17618), .B2(n16785), .ZN(
        n8980) );
  OAI22_X1 U7099 ( .A1(n17995), .A2(n16020), .B1(n17990), .B2(n16786), .ZN(
        n8989) );
  OAI22_X1 U7100 ( .A1(n17622), .A2(n16159), .B1(n17618), .B2(n16791), .ZN(
        n9052) );
  OAI22_X1 U7101 ( .A1(n17995), .A2(n16021), .B1(n17990), .B2(n16792), .ZN(
        n9061) );
  OAI22_X1 U7102 ( .A1(n17994), .A2(n16022), .B1(n17990), .B2(n16798), .ZN(
        n9133) );
  OAI22_X1 U7103 ( .A1(n17994), .A2(n16023), .B1(n17990), .B2(n16804), .ZN(
        n9205) );
  OAI22_X1 U7104 ( .A1(n17623), .A2(n16160), .B1(n17618), .B2(n16821), .ZN(
        n9412) );
  OAI22_X1 U7105 ( .A1(n17995), .A2(n16024), .B1(n17990), .B2(n16822), .ZN(
        n9421) );
  OAI22_X1 U7106 ( .A1(n10189), .A2(n14033), .B1(n7588), .B2(n14034), .ZN(
        n10128) );
  OAI22_X1 U7107 ( .A1(n7725), .A2(n17833), .B1(n12370), .B2(n17824), .ZN(
        n7764) );
  NOR4_X1 U7108 ( .A1(n12371), .A2(n12372), .A3(n12373), .A4(n12374), .ZN(
        n12370) );
  NAND4_X1 U7109 ( .A1(n12375), .A2(n12376), .A3(n12377), .A4(n12378), .ZN(
        n12374) );
  NAND4_X1 U7110 ( .A1(n12399), .A2(n12400), .A3(n12401), .A4(n12402), .ZN(
        n12371) );
  OAI22_X1 U7111 ( .A1(n7724), .A2(n17833), .B1(n12216), .B2(n17824), .ZN(
        n7839) );
  NOR4_X1 U7112 ( .A1(n12217), .A2(n12218), .A3(n12219), .A4(n12220), .ZN(
        n12216) );
  NAND4_X1 U7113 ( .A1(n12221), .A2(n12222), .A3(n12223), .A4(n12224), .ZN(
        n12220) );
  NAND4_X1 U7114 ( .A1(n12245), .A2(n12246), .A3(n12247), .A4(n12248), .ZN(
        n12217) );
  OAI22_X1 U7115 ( .A1(n7695), .A2(n17826), .B1(n4091), .B2(n17824), .ZN(n9989) );
  NOR4_X1 U7116 ( .A1(n4095), .A2(n4098), .A3(n4099), .A4(n4100), .ZN(n4091)
         );
  NAND4_X1 U7117 ( .A1(n4101), .A2(n4102), .A3(n4103), .A4(n4106), .ZN(n4100)
         );
  NAND4_X1 U7118 ( .A1(n4213), .A2(n4214), .A3(n4217), .A4(n4218), .ZN(n4095)
         );
  OAI22_X1 U7119 ( .A1(net227471), .A2(n14007), .B1(n14019), .B2(n14009), .ZN(
        n10133) );
  AOI21_X1 U7120 ( .B1(n14021), .B2(\r590/carry[5] ), .A(n14011), .ZN(n14019)
         );
  OAI22_X1 U7121 ( .A1(net227472), .A2(n14007), .B1(n14018), .B2(n14009), .ZN(
        n10134) );
  XNOR2_X1 U7122 ( .A(n10187), .B(n14017), .ZN(n14018) );
  OAI22_X1 U7123 ( .A1(net227473), .A2(n14007), .B1(n14013), .B2(n14009), .ZN(
        n10135) );
  AOI211_X1 U7124 ( .C1(N9909), .C2(N9908), .A(n14016), .B(n14017), .ZN(n14013) );
  OAI22_X1 U7125 ( .A1(net227476), .A2(n14007), .B1(N9641), .B2(n14009), .ZN(
        n10138) );
  OAI22_X1 U7126 ( .A1(n7723), .A2(n17833), .B1(n12061), .B2(n17823), .ZN(
        n7915) );
  NOR4_X1 U7127 ( .A1(n12062), .A2(n12063), .A3(n12064), .A4(n12065), .ZN(
        n12061) );
  NAND4_X1 U7128 ( .A1(n12066), .A2(n12067), .A3(n12068), .A4(n12069), .ZN(
        n12065) );
  NAND4_X1 U7129 ( .A1(n12090), .A2(n12091), .A3(n12092), .A4(n12093), .ZN(
        n12062) );
  OAI22_X1 U7130 ( .A1(n7722), .A2(n17832), .B1(n11908), .B2(n17825), .ZN(
        n7989) );
  NOR4_X1 U7131 ( .A1(n11909), .A2(n11910), .A3(n11911), .A4(n11912), .ZN(
        n11908) );
  NAND4_X1 U7132 ( .A1(n11913), .A2(n11914), .A3(n11915), .A4(n11916), .ZN(
        n11912) );
  NAND4_X1 U7133 ( .A1(n11937), .A2(n11938), .A3(n11939), .A4(n11940), .ZN(
        n11909) );
  OAI22_X1 U7134 ( .A1(n7721), .A2(n17832), .B1(n10465), .B2(n17823), .ZN(
        n8117) );
  NOR4_X1 U7135 ( .A1(n10466), .A2(n10467), .A3(n10468), .A4(n10469), .ZN(
        n10465) );
  NAND4_X1 U7136 ( .A1(n10470), .A2(n10471), .A3(n10472), .A4(n10473), .ZN(
        n10469) );
  NAND4_X1 U7137 ( .A1(n10494), .A2(n10495), .A3(n10496), .A4(n10497), .ZN(
        n10466) );
  OAI22_X1 U7138 ( .A1(n7720), .A2(n17832), .B1(n10355), .B2(n17825), .ZN(
        n8189) );
  NOR4_X1 U7139 ( .A1(n10356), .A2(n10357), .A3(n10358), .A4(n10359), .ZN(
        n10355) );
  NAND4_X1 U7140 ( .A1(n10360), .A2(n10361), .A3(n10362), .A4(n10363), .ZN(
        n10359) );
  NAND4_X1 U7141 ( .A1(n10384), .A2(n10385), .A3(n10386), .A4(n10387), .ZN(
        n10356) );
  OAI22_X1 U7142 ( .A1(n7719), .A2(n17832), .B1(n10243), .B2(n17823), .ZN(
        n8261) );
  NOR4_X1 U7143 ( .A1(n10244), .A2(n10245), .A3(n10246), .A4(n10247), .ZN(
        n10243) );
  NAND4_X1 U7144 ( .A1(n10248), .A2(n10249), .A3(n10250), .A4(n10251), .ZN(
        n10247) );
  NAND4_X1 U7145 ( .A1(n10272), .A2(n10273), .A3(n10274), .A4(n10275), .ZN(
        n10244) );
  OAI22_X1 U7146 ( .A1(n7718), .A2(n17831), .B1(n7607), .B2(n17825), .ZN(n8333) );
  NOR4_X1 U7147 ( .A1(n7608), .A2(n7609), .A3(n7610), .A4(n7611), .ZN(n7607)
         );
  NAND4_X1 U7148 ( .A1(n7612), .A2(n7613), .A3(n7614), .A4(n7615), .ZN(n7611)
         );
  NAND4_X1 U7149 ( .A1(n7636), .A2(n7637), .A3(n7638), .A4(n7639), .ZN(n7608)
         );
  OAI22_X1 U7150 ( .A1(n7717), .A2(n17831), .B1(n7492), .B2(n17823), .ZN(n8405) );
  NOR4_X1 U7151 ( .A1(n7493), .A2(n7494), .A3(n7495), .A4(n7496), .ZN(n7492)
         );
  NAND4_X1 U7152 ( .A1(n7497), .A2(n7498), .A3(n7499), .A4(n7500), .ZN(n7496)
         );
  NAND4_X1 U7153 ( .A1(n7521), .A2(n7522), .A3(n7523), .A4(n7524), .ZN(n7493)
         );
  OAI22_X1 U7154 ( .A1(n7716), .A2(n17831), .B1(n7383), .B2(n17825), .ZN(n8477) );
  NOR4_X1 U7155 ( .A1(n7384), .A2(n7385), .A3(n7386), .A4(n7387), .ZN(n7383)
         );
  NAND4_X1 U7156 ( .A1(n7388), .A2(n7389), .A3(n7390), .A4(n7391), .ZN(n7387)
         );
  NAND4_X1 U7157 ( .A1(n7412), .A2(n7413), .A3(n7414), .A4(n7415), .ZN(n7384)
         );
  OAI22_X1 U7158 ( .A1(n7715), .A2(n17831), .B1(n7274), .B2(n17823), .ZN(n8549) );
  NOR4_X1 U7159 ( .A1(n7275), .A2(n7276), .A3(n7277), .A4(n7278), .ZN(n7274)
         );
  NAND4_X1 U7160 ( .A1(n7279), .A2(n7280), .A3(n7281), .A4(n7282), .ZN(n7278)
         );
  NAND4_X1 U7161 ( .A1(n7303), .A2(n7304), .A3(n7305), .A4(n7306), .ZN(n7275)
         );
  OAI22_X1 U7162 ( .A1(n7714), .A2(n17830), .B1(n7160), .B2(n17823), .ZN(n8621) );
  NOR4_X1 U7163 ( .A1(n7161), .A2(n7162), .A3(n7163), .A4(n7164), .ZN(n7160)
         );
  NAND4_X1 U7164 ( .A1(n7165), .A2(n7166), .A3(n7167), .A4(n7168), .ZN(n7164)
         );
  NAND4_X1 U7165 ( .A1(n7189), .A2(n7190), .A3(n7191), .A4(n7192), .ZN(n7161)
         );
  OAI22_X1 U7166 ( .A1(n7713), .A2(n17830), .B1(n7051), .B2(n17823), .ZN(n8693) );
  NOR4_X1 U7167 ( .A1(n7052), .A2(n7053), .A3(n7054), .A4(n7055), .ZN(n7051)
         );
  NAND4_X1 U7168 ( .A1(n7056), .A2(n7057), .A3(n7058), .A4(n7059), .ZN(n7055)
         );
  NAND4_X1 U7169 ( .A1(n7080), .A2(n7081), .A3(n7082), .A4(n7083), .ZN(n7052)
         );
  OAI22_X1 U7170 ( .A1(n7712), .A2(n17830), .B1(n6942), .B2(n17825), .ZN(n8765) );
  NOR4_X1 U7171 ( .A1(n6943), .A2(n6944), .A3(n6945), .A4(n6946), .ZN(n6942)
         );
  NAND4_X1 U7172 ( .A1(n6947), .A2(n6948), .A3(n6949), .A4(n6950), .ZN(n6946)
         );
  NAND4_X1 U7173 ( .A1(n6971), .A2(n6972), .A3(n6973), .A4(n6974), .ZN(n6943)
         );
  OAI22_X1 U7174 ( .A1(n7711), .A2(n17830), .B1(n6833), .B2(n17823), .ZN(n8837) );
  NOR4_X1 U7175 ( .A1(n6834), .A2(n6835), .A3(n6836), .A4(n6837), .ZN(n6833)
         );
  NAND4_X1 U7176 ( .A1(n6838), .A2(n6839), .A3(n6840), .A4(n6841), .ZN(n6837)
         );
  NAND4_X1 U7177 ( .A1(n6862), .A2(n6863), .A3(n6864), .A4(n6865), .ZN(n6834)
         );
  OAI22_X1 U7178 ( .A1(n7710), .A2(n17829), .B1(n6724), .B2(n17823), .ZN(n8909) );
  NOR4_X1 U7179 ( .A1(n6725), .A2(n6726), .A3(n6727), .A4(n6728), .ZN(n6724)
         );
  NAND4_X1 U7180 ( .A1(n6729), .A2(n6730), .A3(n6731), .A4(n6732), .ZN(n6728)
         );
  NAND4_X1 U7181 ( .A1(n6753), .A2(n6754), .A3(n6755), .A4(n6756), .ZN(n6725)
         );
  OAI22_X1 U7182 ( .A1(n7709), .A2(n17829), .B1(n6560), .B2(n17825), .ZN(n8981) );
  NOR4_X1 U7183 ( .A1(n6562), .A2(n6563), .A3(n6564), .A4(n6565), .ZN(n6560)
         );
  NAND4_X1 U7184 ( .A1(n6566), .A2(n6568), .A3(n6570), .A4(n6572), .ZN(n6565)
         );
  NAND4_X1 U7185 ( .A1(n6612), .A2(n6614), .A3(n6615), .A4(n6616), .ZN(n6562)
         );
  OAI22_X1 U7186 ( .A1(n7708), .A2(n17829), .B1(n6374), .B2(n17823), .ZN(n9053) );
  NOR4_X1 U7187 ( .A1(n6375), .A2(n6376), .A3(n6377), .A4(n6379), .ZN(n6374)
         );
  NAND4_X1 U7188 ( .A1(n6381), .A2(n6383), .A3(n6384), .A4(n6385), .ZN(n6379)
         );
  NAND4_X1 U7189 ( .A1(n6426), .A2(n6427), .A3(n6428), .A4(n6429), .ZN(n6375)
         );
  OAI22_X1 U7190 ( .A1(n7707), .A2(n17829), .B1(n6187), .B2(n17825), .ZN(n9125) );
  NOR4_X1 U7191 ( .A1(n6188), .A2(n6190), .A3(n6192), .A4(n6194), .ZN(n6187)
         );
  NAND4_X1 U7192 ( .A1(n6195), .A2(n6196), .A3(n6197), .A4(n6198), .ZN(n6194)
         );
  NAND4_X1 U7193 ( .A1(n6239), .A2(n6240), .A3(n6241), .A4(n6244), .ZN(n6188)
         );
  OAI22_X1 U7194 ( .A1(n7706), .A2(n17828), .B1(n6001), .B2(n17825), .ZN(n9197) );
  NOR4_X1 U7195 ( .A1(n6003), .A2(n6005), .A3(n6006), .A4(n6007), .ZN(n6001)
         );
  NAND4_X1 U7196 ( .A1(n6008), .A2(n6009), .A3(n6010), .A4(n6013), .ZN(n6007)
         );
  NAND4_X1 U7197 ( .A1(n6052), .A2(n6055), .A3(n6056), .A4(n6058), .ZN(n6003)
         );
  OAI22_X1 U7198 ( .A1(n7705), .A2(n17828), .B1(n5816), .B2(n17823), .ZN(n9269) );
  NOR4_X1 U7199 ( .A1(n5817), .A2(n5818), .A3(n5819), .A4(n5820), .ZN(n5816)
         );
  NAND4_X1 U7200 ( .A1(n5821), .A2(n5824), .A3(n5825), .A4(n5826), .ZN(n5820)
         );
  NAND4_X1 U7201 ( .A1(n5867), .A2(n5869), .A3(n5870), .A4(n5871), .ZN(n5817)
         );
  OAI22_X1 U7202 ( .A1(n7704), .A2(n17828), .B1(n5629), .B2(n17823), .ZN(n9341) );
  NOR4_X1 U7203 ( .A1(n5630), .A2(n5631), .A3(n5632), .A4(n5635), .ZN(n5629)
         );
  NAND4_X1 U7204 ( .A1(n5636), .A2(n5637), .A3(n5653), .A4(n5654), .ZN(n5635)
         );
  NAND4_X1 U7205 ( .A1(n5681), .A2(n5682), .A3(n5683), .A4(n5684), .ZN(n5630)
         );
  OAI22_X1 U7206 ( .A1(n7703), .A2(n17828), .B1(n5442), .B2(n17823), .ZN(n9413) );
  NOR4_X1 U7207 ( .A1(n5443), .A2(n5446), .A3(n5447), .A4(n5448), .ZN(n5442)
         );
  NAND4_X1 U7208 ( .A1(n5464), .A2(n5465), .A3(n5466), .A4(n5467), .ZN(n5448)
         );
  NAND4_X1 U7209 ( .A1(n5494), .A2(n5495), .A3(n5497), .A4(n5499), .ZN(n5443)
         );
  OAI22_X1 U7210 ( .A1(n7702), .A2(n17827), .B1(n5257), .B2(n17823), .ZN(n9485) );
  NOR4_X1 U7211 ( .A1(n5259), .A2(n5274), .A3(n5275), .A4(n5276), .ZN(n5257)
         );
  NAND4_X1 U7212 ( .A1(n5277), .A2(n5278), .A3(n5279), .A4(n5280), .ZN(n5276)
         );
  NAND4_X1 U7213 ( .A1(n5309), .A2(n5311), .A3(n5312), .A4(n5313), .ZN(n5259)
         );
  OAI22_X1 U7214 ( .A1(n7701), .A2(n17827), .B1(n5106), .B2(n17825), .ZN(n9557) );
  NOR4_X1 U7215 ( .A1(n5107), .A2(n5108), .A3(n5109), .A4(n5110), .ZN(n5106)
         );
  NAND4_X1 U7216 ( .A1(n5111), .A2(n5112), .A3(n5113), .A4(n5115), .ZN(n5110)
         );
  NAND4_X1 U7217 ( .A1(n5138), .A2(n5139), .A3(n5140), .A4(n5141), .ZN(n5107)
         );
  OAI22_X1 U7218 ( .A1(n7700), .A2(n17827), .B1(n4993), .B2(n17825), .ZN(n9629) );
  NOR4_X1 U7219 ( .A1(n4994), .A2(n4995), .A3(n4996), .A4(n4997), .ZN(n4993)
         );
  NAND4_X1 U7220 ( .A1(n4998), .A2(n4999), .A3(n5000), .A4(n5001), .ZN(n4997)
         );
  NAND4_X1 U7221 ( .A1(n5024), .A2(n5025), .A3(n5026), .A4(n5027), .ZN(n4994)
         );
  OAI22_X1 U7222 ( .A1(n3043), .A2(n14033), .B1(n7592), .B2(n14034), .ZN(
        n10132) );
  OAI22_X1 U7223 ( .A1(n10190), .A2(n14033), .B1(n7587), .B2(n14034), .ZN(
        n10127) );
  OAI22_X1 U7224 ( .A1(n10188), .A2(n14033), .B1(n7589), .B2(n14034), .ZN(
        n10129) );
  OAI22_X1 U7225 ( .A1(n10187), .A2(n14033), .B1(n7590), .B2(n14034), .ZN(
        n10130) );
  OAI22_X1 U7226 ( .A1(n14820), .A2(n14033), .B1(n7591), .B2(n14034), .ZN(
        n10131) );
  OAI22_X1 U7227 ( .A1(n17535), .A2(n18027), .B1(n17536), .B2(n16025), .ZN(
        n9982) );
  OAI22_X1 U7228 ( .A1(n17549), .A2(n18027), .B1(n17550), .B2(n16030), .ZN(
        n9983) );
  OAI22_X1 U7229 ( .A1(n17563), .A2(n18027), .B1(n17564), .B2(n16032), .ZN(
        n9984) );
  OAI22_X1 U7230 ( .A1(n17590), .A2(n18027), .B1(n17591), .B2(n16026), .ZN(
        n9986) );
  OAI22_X1 U7231 ( .A1(n17604), .A2(n18026), .B1(n17605), .B2(n16027), .ZN(
        n9987) );
  OAI22_X1 U7232 ( .A1(n17618), .A2(n18026), .B1(n17619), .B2(n16031), .ZN(
        n9988) );
  OAI22_X1 U7233 ( .A1(n17990), .A2(n18026), .B1(n17991), .B2(n15789), .ZN(
        n9997) );
  OAI22_X1 U7234 ( .A1(n16901), .A2(n18031), .B1(n15788), .B2(n16902), .ZN(
        n10003) );
  OAI22_X1 U7235 ( .A1(n16990), .A2(n18031), .B1(n15787), .B2(n16991), .ZN(
        n10011) );
  OAI22_X1 U7236 ( .A1(n17151), .A2(n18029), .B1(n15783), .B2(n17152), .ZN(
        n10024) );
  OAI22_X1 U7237 ( .A1(n17217), .A2(n18029), .B1(n15786), .B2(n17218), .ZN(
        n10030) );
  OAI22_X1 U7238 ( .A1(n17269), .A2(n18029), .B1(n15784), .B2(n17270), .ZN(
        n10034) );
  OAI22_X1 U7239 ( .A1(n17549), .A2(n16701), .B1(n17550), .B2(n16033), .ZN(
        n10055) );
  OAI22_X1 U7240 ( .A1(n17563), .A2(n16701), .B1(n17564), .B2(n16035), .ZN(
        n10056) );
  OAI22_X1 U7241 ( .A1(n17590), .A2(n16701), .B1(n17591), .B2(n16029), .ZN(
        n10058) );
  OAI22_X1 U7242 ( .A1(n17604), .A2(n16701), .B1(n17605), .B2(n16028), .ZN(
        n10059) );
  OAI22_X1 U7243 ( .A1(n17618), .A2(n16701), .B1(n17619), .B2(n16034), .ZN(
        n10060) );
  OAI22_X1 U7244 ( .A1(n17990), .A2(n16702), .B1(n17991), .B2(n15790), .ZN(
        n10069) );
  OAI22_X1 U7245 ( .A1(n17570), .A2(n16186), .B1(n17563), .B2(n16731), .ZN(
        n8328) );
  OAI22_X1 U7246 ( .A1(n17597), .A2(n16060), .B1(n17590), .B2(n16731), .ZN(
        n8330) );
  OAI22_X1 U7247 ( .A1(n17611), .A2(n16098), .B1(n17604), .B2(n16731), .ZN(
        n8331) );
  OAI22_X1 U7248 ( .A1(n17556), .A2(n16161), .B1(n17549), .B2(n16737), .ZN(
        n8399) );
  OAI22_X1 U7249 ( .A1(n17570), .A2(n16187), .B1(n17563), .B2(n16737), .ZN(
        n8400) );
  OAI22_X1 U7250 ( .A1(n17597), .A2(n16061), .B1(n17590), .B2(n16737), .ZN(
        n8402) );
  OAI22_X1 U7251 ( .A1(n17611), .A2(n16099), .B1(n17604), .B2(n16737), .ZN(
        n8403) );
  OAI22_X1 U7252 ( .A1(n17541), .A2(n16062), .B1(n17535), .B2(n16743), .ZN(
        n8470) );
  OAI22_X1 U7253 ( .A1(n17555), .A2(n16162), .B1(n17549), .B2(n16743), .ZN(
        n8471) );
  OAI22_X1 U7254 ( .A1(n17569), .A2(n16188), .B1(n17563), .B2(n16743), .ZN(
        n8472) );
  OAI22_X1 U7255 ( .A1(n17596), .A2(n16063), .B1(n17590), .B2(n16743), .ZN(
        n8474) );
  OAI22_X1 U7256 ( .A1(n17610), .A2(n16100), .B1(n17604), .B2(n16743), .ZN(
        n8475) );
  OAI22_X1 U7257 ( .A1(n17541), .A2(n16064), .B1(n17535), .B2(n16749), .ZN(
        n8542) );
  OAI22_X1 U7258 ( .A1(n17555), .A2(n16163), .B1(n17549), .B2(n16749), .ZN(
        n8543) );
  OAI22_X1 U7259 ( .A1(n17569), .A2(n16189), .B1(n17563), .B2(n16749), .ZN(
        n8544) );
  OAI22_X1 U7260 ( .A1(n17596), .A2(n16065), .B1(n17590), .B2(n16749), .ZN(
        n8546) );
  OAI22_X1 U7261 ( .A1(n17610), .A2(n16101), .B1(n17604), .B2(n16749), .ZN(
        n8547) );
  OAI22_X1 U7262 ( .A1(n16873), .A2(n15956), .B1(n16867), .B2(n16750), .ZN(
        n8560) );
  OAI22_X1 U7263 ( .A1(n17541), .A2(n16066), .B1(n17535), .B2(n16755), .ZN(
        n8614) );
  OAI22_X1 U7264 ( .A1(n17555), .A2(n16164), .B1(n17549), .B2(n16755), .ZN(
        n8615) );
  OAI22_X1 U7265 ( .A1(n17569), .A2(n16190), .B1(n17563), .B2(n16755), .ZN(
        n8616) );
  OAI22_X1 U7266 ( .A1(n17596), .A2(n16067), .B1(n17590), .B2(n16755), .ZN(
        n8618) );
  OAI22_X1 U7267 ( .A1(n17610), .A2(n16102), .B1(n17604), .B2(n16755), .ZN(
        n8619) );
  OAI22_X1 U7268 ( .A1(n16873), .A2(n15957), .B1(n16867), .B2(n16756), .ZN(
        n8632) );
  OAI22_X1 U7269 ( .A1(n17540), .A2(n16068), .B1(n17535), .B2(n16761), .ZN(
        n8686) );
  OAI22_X1 U7270 ( .A1(n17555), .A2(n16165), .B1(n17549), .B2(n16761), .ZN(
        n8687) );
  OAI22_X1 U7271 ( .A1(n17569), .A2(n16191), .B1(n17563), .B2(n16761), .ZN(
        n8688) );
  OAI22_X1 U7272 ( .A1(n17596), .A2(n16069), .B1(n17590), .B2(n16761), .ZN(
        n8690) );
  OAI22_X1 U7273 ( .A1(n17610), .A2(n16103), .B1(n17604), .B2(n16761), .ZN(
        n8691) );
  OAI22_X1 U7274 ( .A1(n16873), .A2(n15958), .B1(n16867), .B2(n16762), .ZN(
        n8704) );
  OAI22_X1 U7275 ( .A1(n17540), .A2(n16070), .B1(n17535), .B2(n16767), .ZN(
        n8758) );
  OAI22_X1 U7276 ( .A1(n17554), .A2(n16166), .B1(n17549), .B2(n16767), .ZN(
        n8759) );
  OAI22_X1 U7277 ( .A1(n17568), .A2(n16192), .B1(n17563), .B2(n16767), .ZN(
        n8760) );
  OAI22_X1 U7278 ( .A1(n17595), .A2(n16071), .B1(n17590), .B2(n16767), .ZN(
        n8762) );
  OAI22_X1 U7279 ( .A1(n17609), .A2(n16104), .B1(n17604), .B2(n16767), .ZN(
        n8763) );
  OAI22_X1 U7280 ( .A1(n16872), .A2(n15959), .B1(n16867), .B2(n16768), .ZN(
        n8776) );
  OAI22_X1 U7281 ( .A1(n17540), .A2(n16072), .B1(n17535), .B2(n16773), .ZN(
        n8830) );
  OAI22_X1 U7282 ( .A1(n17554), .A2(n16167), .B1(n17549), .B2(n16773), .ZN(
        n8831) );
  OAI22_X1 U7283 ( .A1(n17568), .A2(n16193), .B1(n17563), .B2(n16773), .ZN(
        n8832) );
  OAI22_X1 U7284 ( .A1(n17595), .A2(n16073), .B1(n17590), .B2(n16773), .ZN(
        n8834) );
  OAI22_X1 U7285 ( .A1(n17609), .A2(n16105), .B1(n17604), .B2(n16773), .ZN(
        n8835) );
  OAI22_X1 U7286 ( .A1(n16872), .A2(n15960), .B1(n16867), .B2(n16774), .ZN(
        n8848) );
  OAI22_X1 U7287 ( .A1(n17539), .A2(n16074), .B1(n17535), .B2(n16779), .ZN(
        n8902) );
  OAI22_X1 U7288 ( .A1(n17554), .A2(n16168), .B1(n17549), .B2(n16779), .ZN(
        n8903) );
  OAI22_X1 U7289 ( .A1(n17568), .A2(n16194), .B1(n17563), .B2(n16779), .ZN(
        n8904) );
  OAI22_X1 U7290 ( .A1(n17595), .A2(n16075), .B1(n17590), .B2(n16779), .ZN(
        n8906) );
  OAI22_X1 U7291 ( .A1(n17609), .A2(n16106), .B1(n17604), .B2(n16779), .ZN(
        n8907) );
  OAI22_X1 U7292 ( .A1(n16872), .A2(n15961), .B1(n16867), .B2(n16780), .ZN(
        n8920) );
  OAI22_X1 U7293 ( .A1(n17539), .A2(n16076), .B1(n17535), .B2(n16785), .ZN(
        n8974) );
  OAI22_X1 U7294 ( .A1(n17553), .A2(n16169), .B1(n17549), .B2(n16785), .ZN(
        n8975) );
  OAI22_X1 U7295 ( .A1(n17567), .A2(n16195), .B1(n17563), .B2(n16785), .ZN(
        n8976) );
  OAI22_X1 U7296 ( .A1(n17594), .A2(n16077), .B1(n17590), .B2(n16785), .ZN(
        n8978) );
  OAI22_X1 U7297 ( .A1(n17608), .A2(n16107), .B1(n17604), .B2(n16785), .ZN(
        n8979) );
  OAI22_X1 U7298 ( .A1(n16871), .A2(n15962), .B1(n16867), .B2(n16786), .ZN(
        n8992) );
  OAI22_X1 U7299 ( .A1(n17539), .A2(n16078), .B1(n17535), .B2(n16791), .ZN(
        n9046) );
  OAI22_X1 U7300 ( .A1(n17553), .A2(n16170), .B1(n17549), .B2(n16791), .ZN(
        n9047) );
  OAI22_X1 U7301 ( .A1(n17567), .A2(n16196), .B1(n17563), .B2(n16791), .ZN(
        n9048) );
  OAI22_X1 U7302 ( .A1(n17594), .A2(n16079), .B1(n17590), .B2(n16791), .ZN(
        n9050) );
  OAI22_X1 U7303 ( .A1(n17608), .A2(n16108), .B1(n17604), .B2(n16791), .ZN(
        n9051) );
  OAI22_X1 U7304 ( .A1(n16871), .A2(n15963), .B1(n16867), .B2(n16792), .ZN(
        n9064) );
  OAI22_X1 U7305 ( .A1(n17539), .A2(n16080), .B1(n17535), .B2(n16797), .ZN(
        n9118) );
  OAI22_X1 U7306 ( .A1(n17553), .A2(n16171), .B1(n17549), .B2(n16797), .ZN(
        n9119) );
  OAI22_X1 U7307 ( .A1(n17567), .A2(n16197), .B1(n17563), .B2(n16797), .ZN(
        n9120) );
  OAI22_X1 U7308 ( .A1(n17594), .A2(n16081), .B1(n17590), .B2(n16797), .ZN(
        n9122) );
  OAI22_X1 U7309 ( .A1(n17608), .A2(n16109), .B1(n17604), .B2(n16797), .ZN(
        n9123) );
  OAI22_X1 U7310 ( .A1(n16871), .A2(n15964), .B1(n16867), .B2(n16798), .ZN(
        n9136) );
  OAI22_X1 U7311 ( .A1(n17553), .A2(n16172), .B1(n17549), .B2(n16803), .ZN(
        n9191) );
  OAI22_X1 U7312 ( .A1(n16871), .A2(n15965), .B1(n16867), .B2(n16804), .ZN(
        n9208) );
  OAI22_X1 U7313 ( .A1(n17538), .A2(n16082), .B1(n17535), .B2(n16809), .ZN(
        n9262) );
  OAI22_X1 U7314 ( .A1(n16870), .A2(n15966), .B1(n16867), .B2(n16810), .ZN(
        n9280) );
  OAI22_X1 U7315 ( .A1(n16870), .A2(n15967), .B1(n16867), .B2(n16816), .ZN(
        n9352) );
  OAI22_X1 U7316 ( .A1(n17540), .A2(n16083), .B1(n17535), .B2(n16821), .ZN(
        n9406) );
  OAI22_X1 U7317 ( .A1(n17554), .A2(n16173), .B1(n17549), .B2(n16821), .ZN(
        n9407) );
  OAI22_X1 U7318 ( .A1(n17568), .A2(n16198), .B1(n17563), .B2(n16821), .ZN(
        n9408) );
  OAI22_X1 U7319 ( .A1(n17595), .A2(n16084), .B1(n17590), .B2(n16821), .ZN(
        n9410) );
  OAI22_X1 U7320 ( .A1(n17609), .A2(n16110), .B1(n17604), .B2(n16821), .ZN(
        n9411) );
  OAI22_X1 U7321 ( .A1(n16872), .A2(n15968), .B1(n16867), .B2(n17513), .ZN(
        n9928) );
  OAI22_X1 U7322 ( .A1(n17521), .A2(n18027), .B1(n15785), .B2(n17523), .ZN(
        n10053) );
  OAI22_X1 U7323 ( .A1(n17538), .A2(n16085), .B1(n17535), .B2(n16803), .ZN(
        n9190) );
  NAND2_X1 U7324 ( .A1(\sub_132/carry[4] ), .A2(add_rd1[4]), .ZN(n12502) );
  NOR2_X1 U7325 ( .A1(n14265), .A2(n7592), .ZN(n14231) );
  NAND4_X1 U7326 ( .A1(n12509), .A2(n12510), .A3(n12511), .A4(n12512), .ZN(
        n12492) );
  XNOR2_X1 U7327 ( .A(N45542), .B(N190), .ZN(n12510) );
  XNOR2_X1 U7328 ( .A(N45543), .B(N191), .ZN(n12511) );
  XNOR2_X1 U7329 ( .A(add_rd1[4]), .B(add_wr[4]), .ZN(n12509) );
  INV_X1 U7330 ( .A(n14023), .ZN(n14025) );
  NAND2_X1 U7331 ( .A1(\sub_146/carry[4] ), .A2(add_rd2[4]), .ZN(n13983) );
  NAND4_X1 U7332 ( .A1(n13990), .A2(n13991), .A3(n13992), .A4(n13993), .ZN(
        n13973) );
  XNOR2_X1 U7333 ( .A(add_rd2[4]), .B(add_wr[4]), .ZN(n13990) );
  XNOR2_X1 U7334 ( .A(N46056), .B(N190), .ZN(n13991) );
  XNOR2_X1 U7335 ( .A(N46057), .B(N191), .ZN(n13992) );
  NAND2_X1 U7336 ( .A1(n14223), .A2(n14224), .ZN(n14214) );
  INV_X1 U7337 ( .A(N192), .ZN(n14224) );
  NAND2_X1 U7338 ( .A1(n5522), .A2(n14821), .ZN(n14006) );
  AOI21_X1 U7339 ( .B1(n16414), .B2(net226799), .A(n13907), .ZN(n13906) );
  NOR4_X1 U7340 ( .A1(n13908), .A2(n13909), .A3(n13910), .A4(n13911), .ZN(
        n13907) );
  NAND4_X1 U7341 ( .A1(n13964), .A2(n13965), .A3(n13966), .A4(n13967), .ZN(
        n13908) );
  NAND4_X1 U7342 ( .A1(n13948), .A2(n13949), .A3(n13950), .A4(n13951), .ZN(
        n13909) );
  AOI21_X1 U7343 ( .B1(n16417), .B2(net226800), .A(n13860), .ZN(n13859) );
  NOR4_X1 U7344 ( .A1(n13861), .A2(n13862), .A3(n13863), .A4(n13864), .ZN(
        n13860) );
  NAND4_X1 U7345 ( .A1(n13889), .A2(n13890), .A3(n13891), .A4(n13892), .ZN(
        n13861) );
  NAND4_X1 U7346 ( .A1(n13881), .A2(n13882), .A3(n13883), .A4(n13884), .ZN(
        n13862) );
  AOI21_X1 U7347 ( .B1(n16417), .B2(net226801), .A(n13818), .ZN(n13817) );
  NOR4_X1 U7348 ( .A1(n13819), .A2(n13820), .A3(n13821), .A4(n13822), .ZN(
        n13818) );
  NAND4_X1 U7349 ( .A1(n13847), .A2(n13848), .A3(n13849), .A4(n13850), .ZN(
        n13819) );
  NAND4_X1 U7350 ( .A1(n13839), .A2(n13840), .A3(n13841), .A4(n13842), .ZN(
        n13820) );
  AOI21_X1 U7351 ( .B1(n16417), .B2(net226802), .A(n13776), .ZN(n13775) );
  NOR4_X1 U7352 ( .A1(n13777), .A2(n13778), .A3(n13779), .A4(n13780), .ZN(
        n13776) );
  NAND4_X1 U7353 ( .A1(n13805), .A2(n13806), .A3(n13807), .A4(n13808), .ZN(
        n13777) );
  NAND4_X1 U7354 ( .A1(n13797), .A2(n13798), .A3(n13799), .A4(n13800), .ZN(
        n13778) );
  AOI21_X1 U7355 ( .B1(n16416), .B2(net226803), .A(n13734), .ZN(n13733) );
  NOR4_X1 U7356 ( .A1(n13735), .A2(n13736), .A3(n13737), .A4(n13738), .ZN(
        n13734) );
  NAND4_X1 U7357 ( .A1(n13763), .A2(n13764), .A3(n13765), .A4(n13766), .ZN(
        n13735) );
  NAND4_X1 U7358 ( .A1(n13755), .A2(n13756), .A3(n13757), .A4(n13758), .ZN(
        n13736) );
  AOI21_X1 U7359 ( .B1(n16416), .B2(net226804), .A(n13692), .ZN(n13691) );
  NOR4_X1 U7360 ( .A1(n13693), .A2(n13694), .A3(n13695), .A4(n13696), .ZN(
        n13692) );
  NAND4_X1 U7361 ( .A1(n13721), .A2(n13722), .A3(n13723), .A4(n13724), .ZN(
        n13693) );
  NAND4_X1 U7362 ( .A1(n13713), .A2(n13714), .A3(n13715), .A4(n13716), .ZN(
        n13694) );
  AOI21_X1 U7363 ( .B1(n16416), .B2(net226805), .A(n13650), .ZN(n13649) );
  NOR4_X1 U7364 ( .A1(n13651), .A2(n13652), .A3(n13653), .A4(n13654), .ZN(
        n13650) );
  NAND4_X1 U7365 ( .A1(n13679), .A2(n13680), .A3(n13681), .A4(n13682), .ZN(
        n13651) );
  NAND4_X1 U7366 ( .A1(n13671), .A2(n13672), .A3(n13673), .A4(n13674), .ZN(
        n13652) );
  AOI21_X1 U7367 ( .B1(n16416), .B2(net226806), .A(n13608), .ZN(n13607) );
  NOR4_X1 U7368 ( .A1(n13609), .A2(n13610), .A3(n13611), .A4(n13612), .ZN(
        n13608) );
  NAND4_X1 U7369 ( .A1(n13637), .A2(n13638), .A3(n13639), .A4(n13640), .ZN(
        n13609) );
  NAND4_X1 U7370 ( .A1(n13629), .A2(n13630), .A3(n13631), .A4(n13632), .ZN(
        n13610) );
  AOI21_X1 U7371 ( .B1(n16416), .B2(net226807), .A(n13566), .ZN(n13565) );
  NOR4_X1 U7372 ( .A1(n13567), .A2(n13568), .A3(n13569), .A4(n13570), .ZN(
        n13566) );
  NAND4_X1 U7373 ( .A1(n13595), .A2(n13596), .A3(n13597), .A4(n13598), .ZN(
        n13567) );
  NAND4_X1 U7374 ( .A1(n13587), .A2(n13588), .A3(n13589), .A4(n13590), .ZN(
        n13568) );
  AOI21_X1 U7375 ( .B1(n16416), .B2(net226808), .A(n13524), .ZN(n13523) );
  NOR4_X1 U7376 ( .A1(n13525), .A2(n13526), .A3(n13527), .A4(n13528), .ZN(
        n13524) );
  NAND4_X1 U7377 ( .A1(n13553), .A2(n13554), .A3(n13555), .A4(n13556), .ZN(
        n13525) );
  NAND4_X1 U7378 ( .A1(n13545), .A2(n13546), .A3(n13547), .A4(n13548), .ZN(
        n13526) );
  AOI21_X1 U7379 ( .B1(n16416), .B2(net226809), .A(n13482), .ZN(n13481) );
  NOR4_X1 U7380 ( .A1(n13483), .A2(n13484), .A3(n13485), .A4(n13486), .ZN(
        n13482) );
  NAND4_X1 U7381 ( .A1(n13511), .A2(n13512), .A3(n13513), .A4(n13514), .ZN(
        n13483) );
  NAND4_X1 U7382 ( .A1(n13503), .A2(n13504), .A3(n13505), .A4(n13506), .ZN(
        n13484) );
  AOI21_X1 U7383 ( .B1(n16416), .B2(net226810), .A(n13440), .ZN(n13439) );
  NOR4_X1 U7384 ( .A1(n13441), .A2(n13442), .A3(n13443), .A4(n13444), .ZN(
        n13440) );
  NAND4_X1 U7385 ( .A1(n13469), .A2(n13470), .A3(n13471), .A4(n13472), .ZN(
        n13441) );
  NAND4_X1 U7386 ( .A1(n13461), .A2(n13462), .A3(n13463), .A4(n13464), .ZN(
        n13442) );
  AOI21_X1 U7387 ( .B1(n16416), .B2(net226811), .A(n13398), .ZN(n13397) );
  NOR4_X1 U7388 ( .A1(n13399), .A2(n13400), .A3(n13401), .A4(n13402), .ZN(
        n13398) );
  NAND4_X1 U7389 ( .A1(n13427), .A2(n13428), .A3(n13429), .A4(n13430), .ZN(
        n13399) );
  NAND4_X1 U7390 ( .A1(n13419), .A2(n13420), .A3(n13421), .A4(n13422), .ZN(
        n13400) );
  AOI21_X1 U7391 ( .B1(n16416), .B2(net226812), .A(n13356), .ZN(n13355) );
  NOR4_X1 U7392 ( .A1(n13357), .A2(n13358), .A3(n13359), .A4(n13360), .ZN(
        n13356) );
  NAND4_X1 U7393 ( .A1(n13385), .A2(n13386), .A3(n13387), .A4(n13388), .ZN(
        n13357) );
  NAND4_X1 U7394 ( .A1(n13377), .A2(n13378), .A3(n13379), .A4(n13380), .ZN(
        n13358) );
  AOI21_X1 U7395 ( .B1(n16416), .B2(net226813), .A(n13314), .ZN(n13313) );
  NOR4_X1 U7396 ( .A1(n13315), .A2(n13316), .A3(n13317), .A4(n13318), .ZN(
        n13314) );
  NAND4_X1 U7397 ( .A1(n13343), .A2(n13344), .A3(n13345), .A4(n13346), .ZN(
        n13315) );
  NAND4_X1 U7398 ( .A1(n13335), .A2(n13336), .A3(n13337), .A4(n13338), .ZN(
        n13316) );
  AOI21_X1 U7399 ( .B1(n16416), .B2(net226814), .A(n13272), .ZN(n13271) );
  NOR4_X1 U7400 ( .A1(n13273), .A2(n13274), .A3(n13275), .A4(n13276), .ZN(
        n13272) );
  NAND4_X1 U7401 ( .A1(n13301), .A2(n13302), .A3(n13303), .A4(n13304), .ZN(
        n13273) );
  NAND4_X1 U7402 ( .A1(n13293), .A2(n13294), .A3(n13295), .A4(n13296), .ZN(
        n13274) );
  AOI21_X1 U7403 ( .B1(n16416), .B2(net226815), .A(n13230), .ZN(n13229) );
  NOR4_X1 U7404 ( .A1(n13231), .A2(n13232), .A3(n13233), .A4(n13234), .ZN(
        n13230) );
  NAND4_X1 U7405 ( .A1(n13259), .A2(n13260), .A3(n13261), .A4(n13262), .ZN(
        n13231) );
  NAND4_X1 U7406 ( .A1(n13251), .A2(n13252), .A3(n13253), .A4(n13254), .ZN(
        n13232) );
  AOI21_X1 U7407 ( .B1(n16415), .B2(net226816), .A(n13188), .ZN(n13187) );
  NOR4_X1 U7408 ( .A1(n13189), .A2(n13190), .A3(n13191), .A4(n13192), .ZN(
        n13188) );
  NAND4_X1 U7409 ( .A1(n13217), .A2(n13218), .A3(n13219), .A4(n13220), .ZN(
        n13189) );
  NAND4_X1 U7410 ( .A1(n13209), .A2(n13210), .A3(n13211), .A4(n13212), .ZN(
        n13190) );
  AOI21_X1 U7411 ( .B1(n16415), .B2(net226817), .A(n13146), .ZN(n13145) );
  NOR4_X1 U7412 ( .A1(n13147), .A2(n13148), .A3(n13149), .A4(n13150), .ZN(
        n13146) );
  NAND4_X1 U7413 ( .A1(n13175), .A2(n13176), .A3(n13177), .A4(n13178), .ZN(
        n13147) );
  NAND4_X1 U7414 ( .A1(n13167), .A2(n13168), .A3(n13169), .A4(n13170), .ZN(
        n13148) );
  AOI21_X1 U7415 ( .B1(n16415), .B2(net226818), .A(n13104), .ZN(n13103) );
  NOR4_X1 U7416 ( .A1(n13105), .A2(n13106), .A3(n13107), .A4(n13108), .ZN(
        n13104) );
  NAND4_X1 U7417 ( .A1(n13133), .A2(n13134), .A3(n13135), .A4(n13136), .ZN(
        n13105) );
  NAND4_X1 U7418 ( .A1(n13125), .A2(n13126), .A3(n13127), .A4(n13128), .ZN(
        n13106) );
  AOI21_X1 U7419 ( .B1(n16415), .B2(net226819), .A(n13062), .ZN(n13061) );
  NOR4_X1 U7420 ( .A1(n13063), .A2(n13064), .A3(n13065), .A4(n13066), .ZN(
        n13062) );
  NAND4_X1 U7421 ( .A1(n13091), .A2(n13092), .A3(n13093), .A4(n13094), .ZN(
        n13063) );
  NAND4_X1 U7422 ( .A1(n13083), .A2(n13084), .A3(n13085), .A4(n13086), .ZN(
        n13064) );
  AOI21_X1 U7423 ( .B1(n16415), .B2(net226820), .A(n13020), .ZN(n13019) );
  NOR4_X1 U7424 ( .A1(n13021), .A2(n13022), .A3(n13023), .A4(n13024), .ZN(
        n13020) );
  NAND4_X1 U7425 ( .A1(n13049), .A2(n13050), .A3(n13051), .A4(n13052), .ZN(
        n13021) );
  NAND4_X1 U7426 ( .A1(n13041), .A2(n13042), .A3(n13043), .A4(n13044), .ZN(
        n13022) );
  AOI21_X1 U7427 ( .B1(n16415), .B2(net226821), .A(n12978), .ZN(n12977) );
  NOR4_X1 U7428 ( .A1(n12979), .A2(n12980), .A3(n12981), .A4(n12982), .ZN(
        n12978) );
  NAND4_X1 U7429 ( .A1(n13007), .A2(n13008), .A3(n13009), .A4(n13010), .ZN(
        n12979) );
  NAND4_X1 U7430 ( .A1(n12999), .A2(n13000), .A3(n13001), .A4(n13002), .ZN(
        n12980) );
  AOI21_X1 U7431 ( .B1(n16415), .B2(net226822), .A(n12936), .ZN(n12935) );
  NOR4_X1 U7432 ( .A1(n12937), .A2(n12938), .A3(n12939), .A4(n12940), .ZN(
        n12936) );
  NAND4_X1 U7433 ( .A1(n12965), .A2(n12966), .A3(n12967), .A4(n12968), .ZN(
        n12937) );
  NAND4_X1 U7434 ( .A1(n12957), .A2(n12958), .A3(n12959), .A4(n12960), .ZN(
        n12938) );
  AOI21_X1 U7435 ( .B1(n16415), .B2(net226823), .A(n12894), .ZN(n12893) );
  NOR4_X1 U7436 ( .A1(n12895), .A2(n12896), .A3(n12897), .A4(n12898), .ZN(
        n12894) );
  NAND4_X1 U7437 ( .A1(n12923), .A2(n12924), .A3(n12925), .A4(n12926), .ZN(
        n12895) );
  NAND4_X1 U7438 ( .A1(n12915), .A2(n12916), .A3(n12917), .A4(n12918), .ZN(
        n12896) );
  AOI21_X1 U7439 ( .B1(n16415), .B2(net226824), .A(n12852), .ZN(n12851) );
  NOR4_X1 U7440 ( .A1(n12853), .A2(n12854), .A3(n12855), .A4(n12856), .ZN(
        n12852) );
  NAND4_X1 U7441 ( .A1(n12881), .A2(n12882), .A3(n12883), .A4(n12884), .ZN(
        n12853) );
  NAND4_X1 U7442 ( .A1(n12873), .A2(n12874), .A3(n12875), .A4(n12876), .ZN(
        n12854) );
  AOI21_X1 U7443 ( .B1(n16415), .B2(net226825), .A(n12810), .ZN(n12809) );
  NOR4_X1 U7444 ( .A1(n12811), .A2(n12812), .A3(n12813), .A4(n12814), .ZN(
        n12810) );
  NAND4_X1 U7445 ( .A1(n12839), .A2(n12840), .A3(n12841), .A4(n12842), .ZN(
        n12811) );
  NAND4_X1 U7446 ( .A1(n12831), .A2(n12832), .A3(n12833), .A4(n12834), .ZN(
        n12812) );
  AOI21_X1 U7447 ( .B1(n16415), .B2(net226826), .A(n12768), .ZN(n12767) );
  NOR4_X1 U7448 ( .A1(n12769), .A2(n12770), .A3(n12771), .A4(n12772), .ZN(
        n12768) );
  NAND4_X1 U7449 ( .A1(n12797), .A2(n12798), .A3(n12799), .A4(n12800), .ZN(
        n12769) );
  NAND4_X1 U7450 ( .A1(n12789), .A2(n12790), .A3(n12791), .A4(n12792), .ZN(
        n12770) );
  AOI21_X1 U7451 ( .B1(n16414), .B2(net226827), .A(n12726), .ZN(n12725) );
  NOR4_X1 U7452 ( .A1(n12727), .A2(n12728), .A3(n12729), .A4(n12730), .ZN(
        n12726) );
  NAND4_X1 U7453 ( .A1(n12755), .A2(n12756), .A3(n12757), .A4(n12758), .ZN(
        n12727) );
  NAND4_X1 U7454 ( .A1(n12747), .A2(n12748), .A3(n12749), .A4(n12750), .ZN(
        n12728) );
  AOI21_X1 U7455 ( .B1(n16415), .B2(net226828), .A(n12684), .ZN(n12683) );
  NOR4_X1 U7456 ( .A1(n12685), .A2(n12686), .A3(n12687), .A4(n12688), .ZN(
        n12684) );
  NAND4_X1 U7457 ( .A1(n12713), .A2(n12714), .A3(n12715), .A4(n12716), .ZN(
        n12685) );
  NAND4_X1 U7458 ( .A1(n12705), .A2(n12706), .A3(n12707), .A4(n12708), .ZN(
        n12686) );
  AOI21_X1 U7459 ( .B1(n16414), .B2(net226829), .A(n12640), .ZN(n12639) );
  NOR4_X1 U7460 ( .A1(n12641), .A2(n12642), .A3(n12643), .A4(n12644), .ZN(
        n12640) );
  NAND4_X1 U7461 ( .A1(n12671), .A2(n12672), .A3(n12673), .A4(n12674), .ZN(
        n12641) );
  NAND4_X1 U7462 ( .A1(n12662), .A2(n12663), .A3(n12664), .A4(n12665), .ZN(
        n12642) );
  AOI21_X1 U7463 ( .B1(n16415), .B2(net226830), .A(n12528), .ZN(n12526) );
  NOR4_X1 U7464 ( .A1(n12529), .A2(n12530), .A3(n12531), .A4(n12532), .ZN(
        n12528) );
  NAND4_X1 U7465 ( .A1(n12608), .A2(n12609), .A3(n12610), .A4(n12611), .ZN(
        n12529) );
  NAND4_X1 U7466 ( .A1(n12582), .A2(n12583), .A3(n12584), .A4(n12585), .ZN(
        n12530) );
  AOI21_X1 U7467 ( .B1(n16666), .B2(net226831), .A(n12426), .ZN(n12425) );
  NOR4_X1 U7468 ( .A1(n12427), .A2(n12428), .A3(n12429), .A4(n12430), .ZN(
        n12426) );
  NAND4_X1 U7469 ( .A1(n12483), .A2(n12484), .A3(n12485), .A4(n12486), .ZN(
        n12427) );
  NAND4_X1 U7470 ( .A1(n12467), .A2(n12468), .A3(n12469), .A4(n12470), .ZN(
        n12428) );
  AOI21_X1 U7471 ( .B1(n16669), .B2(net226851), .A(n12264), .ZN(n12263) );
  NOR4_X1 U7472 ( .A1(n12265), .A2(n12266), .A3(n12267), .A4(n12268), .ZN(
        n12264) );
  NAND4_X1 U7473 ( .A1(n12293), .A2(n12294), .A3(n12295), .A4(n12296), .ZN(
        n12265) );
  NAND4_X1 U7474 ( .A1(n12285), .A2(n12286), .A3(n12287), .A4(n12288), .ZN(
        n12266) );
  AOI21_X1 U7475 ( .B1(n16669), .B2(net226871), .A(n12111), .ZN(n12110) );
  NOR4_X1 U7476 ( .A1(n12112), .A2(n12113), .A3(n12114), .A4(n12115), .ZN(
        n12111) );
  NAND4_X1 U7477 ( .A1(n12140), .A2(n12141), .A3(n12142), .A4(n12143), .ZN(
        n12112) );
  NAND4_X1 U7478 ( .A1(n12132), .A2(n12133), .A3(n12134), .A4(n12135), .ZN(
        n12113) );
  AOI21_X1 U7479 ( .B1(n16669), .B2(net226891), .A(n11958), .ZN(n11957) );
  NOR4_X1 U7480 ( .A1(n11959), .A2(n11960), .A3(n11961), .A4(n11962), .ZN(
        n11958) );
  NAND4_X1 U7481 ( .A1(n11987), .A2(n11988), .A3(n11989), .A4(n11990), .ZN(
        n11959) );
  NAND4_X1 U7482 ( .A1(n11979), .A2(n11980), .A3(n11981), .A4(n11982), .ZN(
        n11960) );
  AOI21_X1 U7483 ( .B1(n16668), .B2(net226911), .A(n11805), .ZN(n11804) );
  NOR4_X1 U7484 ( .A1(n11806), .A2(n11807), .A3(n11808), .A4(n11809), .ZN(
        n11805) );
  NAND4_X1 U7485 ( .A1(n11834), .A2(n11835), .A3(n11836), .A4(n11837), .ZN(
        n11806) );
  NAND4_X1 U7486 ( .A1(n11826), .A2(n11827), .A3(n11828), .A4(n11829), .ZN(
        n11807) );
  AOI21_X1 U7487 ( .B1(n16668), .B2(net226913), .A(n11762), .ZN(n11761) );
  NOR4_X1 U7488 ( .A1(n11763), .A2(n11764), .A3(n11765), .A4(n11766), .ZN(
        n11762) );
  NAND4_X1 U7489 ( .A1(n11791), .A2(n11792), .A3(n11793), .A4(n11794), .ZN(
        n11763) );
  NAND4_X1 U7490 ( .A1(n11783), .A2(n11784), .A3(n11785), .A4(n11786), .ZN(
        n11764) );
  AOI21_X1 U7491 ( .B1(n16668), .B2(net226915), .A(n11719), .ZN(n11718) );
  NOR4_X1 U7492 ( .A1(n11720), .A2(n11721), .A3(n11722), .A4(n11723), .ZN(
        n11719) );
  NAND4_X1 U7493 ( .A1(n11748), .A2(n11749), .A3(n11750), .A4(n11751), .ZN(
        n11720) );
  NAND4_X1 U7494 ( .A1(n11740), .A2(n11741), .A3(n11742), .A4(n11743), .ZN(
        n11721) );
  AOI21_X1 U7495 ( .B1(n16668), .B2(net226917), .A(n11676), .ZN(n11675) );
  NOR4_X1 U7496 ( .A1(n11677), .A2(n11678), .A3(n11679), .A4(n11680), .ZN(
        n11676) );
  NAND4_X1 U7497 ( .A1(n11705), .A2(n11706), .A3(n11707), .A4(n11708), .ZN(
        n11677) );
  NAND4_X1 U7498 ( .A1(n11697), .A2(n11698), .A3(n11699), .A4(n11700), .ZN(
        n11678) );
  AOI21_X1 U7499 ( .B1(n16668), .B2(net226919), .A(n11633), .ZN(n11632) );
  NOR4_X1 U7500 ( .A1(n11634), .A2(n11635), .A3(n11636), .A4(n11637), .ZN(
        n11633) );
  NAND4_X1 U7501 ( .A1(n11662), .A2(n11663), .A3(n11664), .A4(n11665), .ZN(
        n11634) );
  NAND4_X1 U7502 ( .A1(n11654), .A2(n11655), .A3(n11656), .A4(n11657), .ZN(
        n11635) );
  AOI21_X1 U7503 ( .B1(n16668), .B2(net226921), .A(n11590), .ZN(n11589) );
  NOR4_X1 U7504 ( .A1(n11591), .A2(n11592), .A3(n11593), .A4(n11594), .ZN(
        n11590) );
  NAND4_X1 U7505 ( .A1(n11619), .A2(n11620), .A3(n11621), .A4(n11622), .ZN(
        n11591) );
  NAND4_X1 U7506 ( .A1(n11611), .A2(n11612), .A3(n11613), .A4(n11614), .ZN(
        n11592) );
  AOI21_X1 U7507 ( .B1(n16668), .B2(net226923), .A(n11547), .ZN(n11546) );
  NOR4_X1 U7508 ( .A1(n11548), .A2(n11549), .A3(n11550), .A4(n11551), .ZN(
        n11547) );
  NAND4_X1 U7509 ( .A1(n11576), .A2(n11577), .A3(n11578), .A4(n11579), .ZN(
        n11548) );
  NAND4_X1 U7510 ( .A1(n11568), .A2(n11569), .A3(n11570), .A4(n11571), .ZN(
        n11549) );
  AOI21_X1 U7511 ( .B1(n16668), .B2(net226925), .A(n11504), .ZN(n11503) );
  NOR4_X1 U7512 ( .A1(n11505), .A2(n11506), .A3(n11507), .A4(n11508), .ZN(
        n11504) );
  NAND4_X1 U7513 ( .A1(n11533), .A2(n11534), .A3(n11535), .A4(n11536), .ZN(
        n11505) );
  NAND4_X1 U7514 ( .A1(n11525), .A2(n11526), .A3(n11527), .A4(n11528), .ZN(
        n11506) );
  AOI21_X1 U7515 ( .B1(n16668), .B2(net226927), .A(n11460), .ZN(n11459) );
  NOR4_X1 U7516 ( .A1(n11462), .A2(n11463), .A3(n11464), .A4(n11465), .ZN(
        n11460) );
  NAND4_X1 U7517 ( .A1(n11490), .A2(n11491), .A3(n11492), .A4(n11493), .ZN(
        n11462) );
  NAND4_X1 U7518 ( .A1(n11482), .A2(n11483), .A3(n11484), .A4(n11485), .ZN(
        n11463) );
  AOI21_X1 U7519 ( .B1(n16668), .B2(net226929), .A(n11417), .ZN(n11416) );
  NOR4_X1 U7520 ( .A1(n11418), .A2(n11419), .A3(n11420), .A4(n11421), .ZN(
        n11417) );
  NAND4_X1 U7521 ( .A1(n11446), .A2(n11447), .A3(n11448), .A4(n11449), .ZN(
        n11418) );
  NAND4_X1 U7522 ( .A1(n11438), .A2(n11439), .A3(n11440), .A4(n11441), .ZN(
        n11419) );
  AOI21_X1 U7523 ( .B1(n16668), .B2(net226931), .A(n11374), .ZN(n11373) );
  NOR4_X1 U7524 ( .A1(n11375), .A2(n11376), .A3(n11377), .A4(n11378), .ZN(
        n11374) );
  NAND4_X1 U7525 ( .A1(n11403), .A2(n11404), .A3(n11405), .A4(n11406), .ZN(
        n11375) );
  NAND4_X1 U7526 ( .A1(n11395), .A2(n11396), .A3(n11397), .A4(n11398), .ZN(
        n11376) );
  AOI21_X1 U7527 ( .B1(n16668), .B2(net226933), .A(n11331), .ZN(n11330) );
  NOR4_X1 U7528 ( .A1(n11332), .A2(n11333), .A3(n11334), .A4(n11335), .ZN(
        n11331) );
  NAND4_X1 U7529 ( .A1(n11360), .A2(n11361), .A3(n11362), .A4(n11363), .ZN(
        n11332) );
  NAND4_X1 U7530 ( .A1(n11352), .A2(n11353), .A3(n11354), .A4(n11355), .ZN(
        n11333) );
  AOI21_X1 U7531 ( .B1(n16668), .B2(net226935), .A(n11288), .ZN(n11287) );
  NOR4_X1 U7532 ( .A1(n11289), .A2(n11290), .A3(n11291), .A4(n11292), .ZN(
        n11288) );
  NAND4_X1 U7533 ( .A1(n11317), .A2(n11318), .A3(n11319), .A4(n11320), .ZN(
        n11289) );
  NAND4_X1 U7534 ( .A1(n11309), .A2(n11310), .A3(n11311), .A4(n11312), .ZN(
        n11290) );
  AOI21_X1 U7535 ( .B1(n16667), .B2(net226937), .A(n11245), .ZN(n11244) );
  NOR4_X1 U7536 ( .A1(n11246), .A2(n11247), .A3(n11248), .A4(n11249), .ZN(
        n11245) );
  NAND4_X1 U7537 ( .A1(n11274), .A2(n11275), .A3(n11276), .A4(n11277), .ZN(
        n11246) );
  NAND4_X1 U7538 ( .A1(n11266), .A2(n11267), .A3(n11268), .A4(n11269), .ZN(
        n11247) );
  AOI21_X1 U7539 ( .B1(n16667), .B2(net226939), .A(n11202), .ZN(n11201) );
  NOR4_X1 U7540 ( .A1(n11203), .A2(n11204), .A3(n11205), .A4(n11206), .ZN(
        n11202) );
  NAND4_X1 U7541 ( .A1(n11231), .A2(n11232), .A3(n11233), .A4(n11234), .ZN(
        n11203) );
  NAND4_X1 U7542 ( .A1(n11223), .A2(n11224), .A3(n11225), .A4(n11226), .ZN(
        n11204) );
  AOI21_X1 U7543 ( .B1(n16667), .B2(net226941), .A(n11159), .ZN(n11158) );
  NOR4_X1 U7544 ( .A1(n11160), .A2(n11161), .A3(n11162), .A4(n11163), .ZN(
        n11159) );
  NAND4_X1 U7545 ( .A1(n11188), .A2(n11189), .A3(n11190), .A4(n11191), .ZN(
        n11160) );
  NAND4_X1 U7546 ( .A1(n11180), .A2(n11181), .A3(n11182), .A4(n11183), .ZN(
        n11161) );
  AOI21_X1 U7547 ( .B1(n16667), .B2(net226943), .A(n11116), .ZN(n11115) );
  NOR4_X1 U7548 ( .A1(n11117), .A2(n11118), .A3(n11119), .A4(n11120), .ZN(
        n11116) );
  NAND4_X1 U7549 ( .A1(n11145), .A2(n11146), .A3(n11147), .A4(n11148), .ZN(
        n11117) );
  NAND4_X1 U7550 ( .A1(n11137), .A2(n11138), .A3(n11139), .A4(n11140), .ZN(
        n11118) );
  AOI21_X1 U7551 ( .B1(n16667), .B2(net226945), .A(n11073), .ZN(n11072) );
  NOR4_X1 U7552 ( .A1(n11074), .A2(n11075), .A3(n11076), .A4(n11077), .ZN(
        n11073) );
  NAND4_X1 U7553 ( .A1(n11102), .A2(n11103), .A3(n11104), .A4(n11105), .ZN(
        n11074) );
  NAND4_X1 U7554 ( .A1(n11094), .A2(n11095), .A3(n11096), .A4(n11097), .ZN(
        n11075) );
  AOI21_X1 U7555 ( .B1(n16667), .B2(net226947), .A(n11030), .ZN(n11029) );
  NOR4_X1 U7556 ( .A1(n11031), .A2(n11032), .A3(n11033), .A4(n11034), .ZN(
        n11030) );
  NAND4_X1 U7557 ( .A1(n11059), .A2(n11060), .A3(n11061), .A4(n11062), .ZN(
        n11031) );
  NAND4_X1 U7558 ( .A1(n11051), .A2(n11052), .A3(n11053), .A4(n11054), .ZN(
        n11032) );
  AOI21_X1 U7559 ( .B1(n16667), .B2(net226949), .A(n10987), .ZN(n10986) );
  NOR4_X1 U7560 ( .A1(n10988), .A2(n10989), .A3(n10990), .A4(n10991), .ZN(
        n10987) );
  NAND4_X1 U7561 ( .A1(n11016), .A2(n11017), .A3(n11018), .A4(n11019), .ZN(
        n10988) );
  NAND4_X1 U7562 ( .A1(n11008), .A2(n11009), .A3(n11010), .A4(n11011), .ZN(
        n10989) );
  AOI21_X1 U7563 ( .B1(n16667), .B2(net226951), .A(n10944), .ZN(n10943) );
  NOR4_X1 U7564 ( .A1(n10945), .A2(n10946), .A3(n10947), .A4(n10948), .ZN(
        n10944) );
  NAND4_X1 U7565 ( .A1(n10973), .A2(n10974), .A3(n10975), .A4(n10976), .ZN(
        n10945) );
  NAND4_X1 U7566 ( .A1(n10965), .A2(n10966), .A3(n10967), .A4(n10968), .ZN(
        n10946) );
  AOI21_X1 U7567 ( .B1(n16667), .B2(net226953), .A(n10901), .ZN(n10900) );
  NOR4_X1 U7568 ( .A1(n10902), .A2(n10903), .A3(n10904), .A4(n10905), .ZN(
        n10901) );
  NAND4_X1 U7569 ( .A1(n10930), .A2(n10931), .A3(n10932), .A4(n10933), .ZN(
        n10902) );
  NAND4_X1 U7570 ( .A1(n10922), .A2(n10923), .A3(n10924), .A4(n10925), .ZN(
        n10903) );
  AOI21_X1 U7571 ( .B1(n16667), .B2(net226955), .A(n10858), .ZN(n10857) );
  NOR4_X1 U7572 ( .A1(n10859), .A2(n10860), .A3(n10861), .A4(n10862), .ZN(
        n10858) );
  NAND4_X1 U7573 ( .A1(n10887), .A2(n10888), .A3(n10889), .A4(n10890), .ZN(
        n10859) );
  NAND4_X1 U7574 ( .A1(n10879), .A2(n10880), .A3(n10881), .A4(n10882), .ZN(
        n10860) );
  AOI21_X1 U7575 ( .B1(n16667), .B2(net226957), .A(n10815), .ZN(n10814) );
  NOR4_X1 U7576 ( .A1(n10816), .A2(n10817), .A3(n10818), .A4(n10819), .ZN(
        n10815) );
  NAND4_X1 U7577 ( .A1(n10844), .A2(n10845), .A3(n10846), .A4(n10847), .ZN(
        n10816) );
  NAND4_X1 U7578 ( .A1(n10836), .A2(n10837), .A3(n10838), .A4(n10839), .ZN(
        n10817) );
  AOI21_X1 U7579 ( .B1(n16666), .B2(net226959), .A(n10772), .ZN(n10771) );
  NOR4_X1 U7580 ( .A1(n10773), .A2(n10774), .A3(n10775), .A4(n10776), .ZN(
        n10772) );
  NAND4_X1 U7581 ( .A1(n10801), .A2(n10802), .A3(n10803), .A4(n10804), .ZN(
        n10773) );
  NAND4_X1 U7582 ( .A1(n10793), .A2(n10794), .A3(n10795), .A4(n10796), .ZN(
        n10774) );
  AOI21_X1 U7583 ( .B1(n16667), .B2(net226961), .A(n10729), .ZN(n10728) );
  NOR4_X1 U7584 ( .A1(n10730), .A2(n10731), .A3(n10732), .A4(n10733), .ZN(
        n10729) );
  NAND4_X1 U7585 ( .A1(n10758), .A2(n10759), .A3(n10760), .A4(n10761), .ZN(
        n10730) );
  NAND4_X1 U7586 ( .A1(n10750), .A2(n10751), .A3(n10752), .A4(n10753), .ZN(
        n10731) );
  AOI21_X1 U7587 ( .B1(n16666), .B2(net226963), .A(n10670), .ZN(n10669) );
  NOR4_X1 U7588 ( .A1(n10671), .A2(n10672), .A3(n10673), .A4(n10674), .ZN(
        n10670) );
  NAND4_X1 U7589 ( .A1(n10713), .A2(n10714), .A3(n10715), .A4(n10716), .ZN(
        n10671) );
  NAND4_X1 U7590 ( .A1(n10700), .A2(n10701), .A3(n10702), .A4(n10703), .ZN(
        n10672) );
  AOI21_X1 U7591 ( .B1(n16667), .B2(net226965), .A(n10526), .ZN(n10524) );
  NOR4_X1 U7592 ( .A1(n10527), .A2(n10528), .A3(n10529), .A4(n10530), .ZN(
        n10526) );
  NAND4_X1 U7593 ( .A1(n10628), .A2(n10629), .A3(n10630), .A4(n10631), .ZN(
        n10527) );
  NAND4_X1 U7594 ( .A1(n10596), .A2(n10597), .A3(n10598), .A4(n10599), .ZN(
        n10528) );
  NAND2_X1 U7595 ( .A1(call), .A2(n14133), .ZN(n14122) );
  NAND4_X1 U7596 ( .A1(n12907), .A2(n12908), .A3(n12909), .A4(n12910), .ZN(
        n12897) );
  AOI221_X1 U7597 ( .B1(net227339), .B2(n16351), .C1(\registers[30][24] ), 
        .C2(n16348), .A(n12912), .ZN(n12909) );
  AOI221_X1 U7598 ( .B1(\registers[10][24] ), .B2(n16327), .C1(
        \registers[0][24] ), .C2(n16324), .A(n12914), .ZN(n12907) );
  AOI221_X1 U7599 ( .B1(net227338), .B2(n16339), .C1(\registers[34][24] ), 
        .C2(n16336), .A(n12913), .ZN(n12908) );
  NAND4_X1 U7600 ( .A1(n12865), .A2(n12866), .A3(n12867), .A4(n12868), .ZN(
        n12855) );
  AOI221_X1 U7601 ( .B1(net227357), .B2(n16351), .C1(\registers[30][25] ), 
        .C2(n16348), .A(n12870), .ZN(n12867) );
  AOI221_X1 U7602 ( .B1(\registers[10][25] ), .B2(n16327), .C1(
        \registers[0][25] ), .C2(n16324), .A(n12872), .ZN(n12865) );
  AOI221_X1 U7603 ( .B1(net227356), .B2(n16339), .C1(\registers[34][25] ), 
        .C2(n16336), .A(n12871), .ZN(n12866) );
  NAND4_X1 U7604 ( .A1(n12823), .A2(n12824), .A3(n12825), .A4(n12826), .ZN(
        n12813) );
  AOI221_X1 U7605 ( .B1(net227375), .B2(n16351), .C1(\registers[30][26] ), 
        .C2(n16348), .A(n12828), .ZN(n12825) );
  AOI221_X1 U7606 ( .B1(\registers[10][26] ), .B2(n16327), .C1(
        \registers[0][26] ), .C2(n16324), .A(n12830), .ZN(n12823) );
  AOI221_X1 U7607 ( .B1(net227374), .B2(n16339), .C1(\registers[34][26] ), 
        .C2(n16336), .A(n12829), .ZN(n12824) );
  NAND4_X1 U7608 ( .A1(n12781), .A2(n12782), .A3(n12783), .A4(n12784), .ZN(
        n12771) );
  AOI221_X1 U7609 ( .B1(net227393), .B2(n16351), .C1(\registers[30][27] ), 
        .C2(n16348), .A(n12786), .ZN(n12783) );
  AOI221_X1 U7610 ( .B1(\registers[10][27] ), .B2(n16327), .C1(
        \registers[0][27] ), .C2(n16324), .A(n12788), .ZN(n12781) );
  AOI221_X1 U7611 ( .B1(net227392), .B2(n16339), .C1(\registers[34][27] ), 
        .C2(n16336), .A(n12787), .ZN(n12782) );
  NAND4_X1 U7612 ( .A1(n12739), .A2(n12740), .A3(n12741), .A4(n12742), .ZN(
        n12729) );
  AOI221_X1 U7613 ( .B1(net227411), .B2(n16351), .C1(\registers[30][28] ), 
        .C2(n16348), .A(n12744), .ZN(n12741) );
  AOI221_X1 U7614 ( .B1(\registers[10][28] ), .B2(n16327), .C1(
        \registers[0][28] ), .C2(n16324), .A(n12746), .ZN(n12739) );
  AOI221_X1 U7615 ( .B1(net227410), .B2(n16339), .C1(\registers[34][28] ), 
        .C2(n16336), .A(n12745), .ZN(n12740) );
  NAND4_X1 U7616 ( .A1(n12697), .A2(n12698), .A3(n12699), .A4(n12700), .ZN(
        n12687) );
  AOI221_X1 U7617 ( .B1(net227429), .B2(n16351), .C1(\registers[30][29] ), 
        .C2(n16348), .A(n12702), .ZN(n12699) );
  AOI221_X1 U7618 ( .B1(\registers[10][29] ), .B2(n16327), .C1(
        \registers[0][29] ), .C2(n16324), .A(n12704), .ZN(n12697) );
  AOI221_X1 U7619 ( .B1(net227428), .B2(n16339), .C1(\registers[34][29] ), 
        .C2(n16336), .A(n12703), .ZN(n12698) );
  NAND4_X1 U7620 ( .A1(n12654), .A2(n12655), .A3(n12656), .A4(n12657), .ZN(
        n12643) );
  AOI221_X1 U7621 ( .B1(net227447), .B2(n16351), .C1(\registers[30][30] ), 
        .C2(n16348), .A(n12659), .ZN(n12656) );
  AOI221_X1 U7622 ( .B1(\registers[10][30] ), .B2(n16327), .C1(
        \registers[0][30] ), .C2(n16324), .A(n12661), .ZN(n12654) );
  AOI221_X1 U7623 ( .B1(net227446), .B2(n16339), .C1(\registers[34][30] ), 
        .C2(n16336), .A(n12660), .ZN(n12655) );
  NAND4_X1 U7624 ( .A1(n12557), .A2(n12558), .A3(n12559), .A4(n12560), .ZN(
        n12531) );
  AOI221_X1 U7625 ( .B1(net227465), .B2(n16351), .C1(\registers[30][31] ), 
        .C2(n16348), .A(n12569), .ZN(n12559) );
  AOI221_X1 U7626 ( .B1(\registers[10][31] ), .B2(n16327), .C1(
        \registers[0][31] ), .C2(n16324), .A(n12579), .ZN(n12557) );
  AOI221_X1 U7627 ( .B1(net227464), .B2(n16339), .C1(\registers[34][31] ), 
        .C2(n16336), .A(n12574), .ZN(n12558) );
  NAND4_X1 U7628 ( .A1(n10957), .A2(n10958), .A3(n10959), .A4(n10960), .ZN(
        n10947) );
  AOI221_X1 U7629 ( .B1(net227339), .B2(n16603), .C1(\registers[30][24] ), 
        .C2(n16600), .A(n10962), .ZN(n10959) );
  AOI221_X1 U7630 ( .B1(\registers[10][24] ), .B2(n16579), .C1(
        \registers[0][24] ), .C2(n16576), .A(n10964), .ZN(n10957) );
  AOI221_X1 U7631 ( .B1(net227338), .B2(n16591), .C1(\registers[34][24] ), 
        .C2(n16588), .A(n10963), .ZN(n10958) );
  NAND4_X1 U7632 ( .A1(n10914), .A2(n10915), .A3(n10916), .A4(n10917), .ZN(
        n10904) );
  AOI221_X1 U7633 ( .B1(net227357), .B2(n16603), .C1(\registers[30][25] ), 
        .C2(n16600), .A(n10919), .ZN(n10916) );
  AOI221_X1 U7634 ( .B1(\registers[10][25] ), .B2(n16579), .C1(
        \registers[0][25] ), .C2(n16576), .A(n10921), .ZN(n10914) );
  AOI221_X1 U7635 ( .B1(net227356), .B2(n16591), .C1(\registers[34][25] ), 
        .C2(n16588), .A(n10920), .ZN(n10915) );
  NAND4_X1 U7636 ( .A1(n10871), .A2(n10872), .A3(n10873), .A4(n10874), .ZN(
        n10861) );
  AOI221_X1 U7637 ( .B1(net227375), .B2(n16603), .C1(\registers[30][26] ), 
        .C2(n16600), .A(n10876), .ZN(n10873) );
  AOI221_X1 U7638 ( .B1(\registers[10][26] ), .B2(n16579), .C1(
        \registers[0][26] ), .C2(n16576), .A(n10878), .ZN(n10871) );
  AOI221_X1 U7639 ( .B1(net227374), .B2(n16591), .C1(\registers[34][26] ), 
        .C2(n16588), .A(n10877), .ZN(n10872) );
  NAND4_X1 U7640 ( .A1(n10828), .A2(n10829), .A3(n10830), .A4(n10831), .ZN(
        n10818) );
  AOI221_X1 U7641 ( .B1(net227393), .B2(n16603), .C1(\registers[30][27] ), 
        .C2(n16600), .A(n10833), .ZN(n10830) );
  AOI221_X1 U7642 ( .B1(\registers[10][27] ), .B2(n16579), .C1(
        \registers[0][27] ), .C2(n16576), .A(n10835), .ZN(n10828) );
  AOI221_X1 U7643 ( .B1(net227392), .B2(n16591), .C1(\registers[34][27] ), 
        .C2(n16588), .A(n10834), .ZN(n10829) );
  NAND4_X1 U7644 ( .A1(n10785), .A2(n10786), .A3(n10787), .A4(n10788), .ZN(
        n10775) );
  AOI221_X1 U7645 ( .B1(net227411), .B2(n16603), .C1(\registers[30][28] ), 
        .C2(n16600), .A(n10790), .ZN(n10787) );
  AOI221_X1 U7646 ( .B1(\registers[10][28] ), .B2(n16579), .C1(
        \registers[0][28] ), .C2(n16576), .A(n10792), .ZN(n10785) );
  AOI221_X1 U7647 ( .B1(net227410), .B2(n16591), .C1(\registers[34][28] ), 
        .C2(n16588), .A(n10791), .ZN(n10786) );
  NAND4_X1 U7648 ( .A1(n10742), .A2(n10743), .A3(n10744), .A4(n10745), .ZN(
        n10732) );
  AOI221_X1 U7649 ( .B1(net227429), .B2(n16603), .C1(\registers[30][29] ), 
        .C2(n16600), .A(n10747), .ZN(n10744) );
  AOI221_X1 U7650 ( .B1(\registers[10][29] ), .B2(n16579), .C1(
        \registers[0][29] ), .C2(n16576), .A(n10749), .ZN(n10742) );
  AOI221_X1 U7651 ( .B1(net227428), .B2(n16591), .C1(\registers[34][29] ), 
        .C2(n16588), .A(n10748), .ZN(n10743) );
  NAND4_X1 U7652 ( .A1(n10687), .A2(n10688), .A3(n10689), .A4(n10690), .ZN(
        n10673) );
  AOI221_X1 U7653 ( .B1(net227447), .B2(n16603), .C1(\registers[30][30] ), 
        .C2(n16600), .A(n10694), .ZN(n10689) );
  AOI221_X1 U7654 ( .B1(\registers[10][30] ), .B2(n16579), .C1(
        \registers[0][30] ), .C2(n16576), .A(n10698), .ZN(n10687) );
  AOI221_X1 U7655 ( .B1(net227446), .B2(n16591), .C1(\registers[34][30] ), 
        .C2(n16588), .A(n10695), .ZN(n10688) );
  NAND4_X1 U7656 ( .A1(n10562), .A2(n10563), .A3(n10564), .A4(n10565), .ZN(
        n10529) );
  AOI221_X1 U7657 ( .B1(net227465), .B2(n16603), .C1(\registers[30][31] ), 
        .C2(n16600), .A(n10577), .ZN(n10564) );
  AOI221_X1 U7658 ( .B1(\registers[10][31] ), .B2(n16579), .C1(
        \registers[0][31] ), .C2(n16576), .A(n10591), .ZN(n10562) );
  AOI221_X1 U7659 ( .B1(net227464), .B2(n16591), .C1(\registers[34][31] ), 
        .C2(n16588), .A(n10584), .ZN(n10563) );
  NAND4_X1 U7660 ( .A1(n5286), .A2(n5288), .A3(n5290), .A4(n5291), .ZN(n5275)
         );
  AOI221_X1 U7661 ( .B1(net227323), .B2(n17759), .C1(\registers[25][23] ), 
        .C2(n17756), .A(n5293), .ZN(n5290) );
  AOI221_X1 U7662 ( .B1(\registers[36][23] ), .B2(n17735), .C1(
        \registers[38][23] ), .C2(n17732), .A(n5295), .ZN(n5286) );
  AOI221_X1 U7663 ( .B1(net227318), .B2(n17771), .C1(\registers[50][23] ), 
        .C2(n17768), .A(n5292), .ZN(n5291) );
  NAND4_X1 U7664 ( .A1(n5120), .A2(n5121), .A3(n5122), .A4(n5123), .ZN(n5109)
         );
  AOI221_X1 U7665 ( .B1(net227341), .B2(n17759), .C1(\registers[25][24] ), 
        .C2(n17756), .A(n5125), .ZN(n5122) );
  AOI221_X1 U7666 ( .B1(\registers[36][24] ), .B2(n17735), .C1(
        \registers[38][24] ), .C2(n17732), .A(n5129), .ZN(n5120) );
  AOI221_X1 U7667 ( .B1(net227336), .B2(n17771), .C1(\registers[50][24] ), 
        .C2(n17768), .A(n5124), .ZN(n5123) );
  NAND4_X1 U7668 ( .A1(n5006), .A2(n5007), .A3(n5008), .A4(n5009), .ZN(n4996)
         );
  AOI221_X1 U7669 ( .B1(net227359), .B2(n17759), .C1(\registers[25][25] ), 
        .C2(n17756), .A(n5011), .ZN(n5008) );
  AOI221_X1 U7670 ( .B1(\registers[36][25] ), .B2(n17735), .C1(
        \registers[38][25] ), .C2(n17732), .A(n5013), .ZN(n5006) );
  AOI221_X1 U7671 ( .B1(net227354), .B2(n17771), .C1(\registers[50][25] ), 
        .C2(n17768), .A(n5010), .ZN(n5009) );
  NAND4_X1 U7672 ( .A1(n4884), .A2(n4885), .A3(n4886), .A4(n4887), .ZN(n4874)
         );
  AOI221_X1 U7673 ( .B1(net227377), .B2(n17759), .C1(\registers[25][26] ), 
        .C2(n17756), .A(n4889), .ZN(n4886) );
  AOI221_X1 U7674 ( .B1(\registers[36][26] ), .B2(n17735), .C1(
        \registers[38][26] ), .C2(n17732), .A(n4891), .ZN(n4884) );
  AOI221_X1 U7675 ( .B1(net227372), .B2(n17771), .C1(\registers[50][26] ), 
        .C2(n17768), .A(n4888), .ZN(n4887) );
  NAND4_X1 U7676 ( .A1(n4757), .A2(n4758), .A3(n4759), .A4(n4760), .ZN(n4741)
         );
  AOI221_X1 U7677 ( .B1(net227395), .B2(n17759), .C1(\registers[25][27] ), 
        .C2(n17756), .A(n4762), .ZN(n4759) );
  AOI221_X1 U7678 ( .B1(\registers[36][27] ), .B2(n17735), .C1(
        \registers[38][27] ), .C2(n17732), .A(n4764), .ZN(n4757) );
  AOI221_X1 U7679 ( .B1(net227390), .B2(n17771), .C1(\registers[50][27] ), 
        .C2(n17768), .A(n4761), .ZN(n4760) );
  NAND4_X1 U7680 ( .A1(n4626), .A2(n4627), .A3(n4628), .A4(n4629), .ZN(n4614)
         );
  AOI221_X1 U7681 ( .B1(net227413), .B2(n17759), .C1(\registers[25][28] ), 
        .C2(n17756), .A(n4631), .ZN(n4628) );
  AOI221_X1 U7682 ( .B1(\registers[36][28] ), .B2(n17735), .C1(
        \registers[38][28] ), .C2(n17732), .A(n4633), .ZN(n4626) );
  AOI221_X1 U7683 ( .B1(net227408), .B2(n17771), .C1(\registers[50][28] ), 
        .C2(n17768), .A(n4630), .ZN(n4629) );
  NAND4_X1 U7684 ( .A1(n4495), .A2(n4498), .A3(n4499), .A4(n4500), .ZN(n4483)
         );
  AOI221_X1 U7685 ( .B1(net227431), .B2(n17759), .C1(\registers[25][29] ), 
        .C2(n17756), .A(n4502), .ZN(n4499) );
  AOI221_X1 U7686 ( .B1(\registers[36][29] ), .B2(n17735), .C1(
        \registers[38][29] ), .C2(n17732), .A(n4506), .ZN(n4495) );
  AOI221_X1 U7687 ( .B1(net227426), .B2(n17771), .C1(\registers[50][29] ), 
        .C2(n17768), .A(n4501), .ZN(n4500) );
  NAND4_X1 U7688 ( .A1(n4137), .A2(n4138), .A3(n4139), .A4(n4140), .ZN(n4099)
         );
  AOI221_X1 U7689 ( .B1(net227449), .B2(n17759), .C1(\registers[25][30] ), 
        .C2(n17756), .A(n4156), .ZN(n4139) );
  AOI221_X1 U7690 ( .B1(\registers[36][30] ), .B2(n17735), .C1(
        \registers[38][30] ), .C2(n17732), .A(n4172), .ZN(n4137) );
  AOI221_X1 U7691 ( .B1(net227444), .B2(n17771), .C1(\registers[50][30] ), 
        .C2(n17768), .A(n4145), .ZN(n4140) );
  NAND4_X1 U7692 ( .A1(n13938), .A2(n13939), .A3(n13940), .A4(n13941), .ZN(
        n13910) );
  AOI221_X1 U7693 ( .B1(net226848), .B2(n16349), .C1(\registers[30][0] ), .C2(
        n16346), .A(n13943), .ZN(n13940) );
  AOI221_X1 U7694 ( .B1(\registers[10][0] ), .B2(n16325), .C1(
        \registers[0][0] ), .C2(n16322), .A(n13947), .ZN(n13938) );
  AOI221_X1 U7695 ( .B1(net226847), .B2(n16337), .C1(\registers[34][0] ), .C2(
        n16334), .A(n13945), .ZN(n13939) );
  NAND4_X1 U7696 ( .A1(n13873), .A2(n13874), .A3(n13875), .A4(n13876), .ZN(
        n13863) );
  AOI221_X1 U7697 ( .B1(net226869), .B2(n16349), .C1(\registers[30][1] ), .C2(
        n16346), .A(n13878), .ZN(n13875) );
  AOI221_X1 U7698 ( .B1(\registers[10][1] ), .B2(n16325), .C1(
        \registers[0][1] ), .C2(n16322), .A(n13880), .ZN(n13873) );
  AOI221_X1 U7699 ( .B1(net226868), .B2(n16337), .C1(\registers[34][1] ), .C2(
        n16334), .A(n13879), .ZN(n13874) );
  NAND4_X1 U7700 ( .A1(n13831), .A2(n13832), .A3(n13833), .A4(n13834), .ZN(
        n13821) );
  AOI221_X1 U7701 ( .B1(net226888), .B2(n16349), .C1(\registers[30][2] ), .C2(
        n16346), .A(n13836), .ZN(n13833) );
  AOI221_X1 U7702 ( .B1(\registers[10][2] ), .B2(n16325), .C1(
        \registers[0][2] ), .C2(n16322), .A(n13838), .ZN(n13831) );
  AOI221_X1 U7703 ( .B1(net226880), .B2(n16337), .C1(\registers[34][2] ), .C2(
        n16334), .A(n13837), .ZN(n13832) );
  NAND4_X1 U7704 ( .A1(n13789), .A2(n13790), .A3(n13791), .A4(n13792), .ZN(
        n13779) );
  AOI221_X1 U7705 ( .B1(net226908), .B2(n16349), .C1(\registers[30][3] ), .C2(
        n16346), .A(n13794), .ZN(n13791) );
  AOI221_X1 U7706 ( .B1(\registers[10][3] ), .B2(n16325), .C1(
        \registers[0][3] ), .C2(n16322), .A(n13796), .ZN(n13789) );
  AOI221_X1 U7707 ( .B1(net226900), .B2(n16337), .C1(\registers[34][3] ), .C2(
        n16334), .A(n13795), .ZN(n13790) );
  NAND4_X1 U7708 ( .A1(n13747), .A2(n13748), .A3(n13749), .A4(n13750), .ZN(
        n13737) );
  AOI221_X1 U7709 ( .B1(net226982), .B2(n16349), .C1(\registers[30][4] ), .C2(
        n16346), .A(n13752), .ZN(n13749) );
  AOI221_X1 U7710 ( .B1(\registers[10][4] ), .B2(n16325), .C1(
        \registers[0][4] ), .C2(n16322), .A(n13754), .ZN(n13747) );
  AOI221_X1 U7711 ( .B1(net226973), .B2(n16337), .C1(\registers[34][4] ), .C2(
        n16334), .A(n13753), .ZN(n13748) );
  NAND4_X1 U7712 ( .A1(n13705), .A2(n13706), .A3(n13707), .A4(n13708), .ZN(
        n13695) );
  AOI221_X1 U7713 ( .B1(net226991), .B2(n16349), .C1(\registers[30][5] ), .C2(
        n16346), .A(n13710), .ZN(n13707) );
  AOI221_X1 U7714 ( .B1(\registers[10][5] ), .B2(n16325), .C1(
        \registers[0][5] ), .C2(n16322), .A(n13712), .ZN(n13705) );
  AOI221_X1 U7715 ( .B1(net226990), .B2(n16337), .C1(\registers[34][5] ), .C2(
        n16334), .A(n13711), .ZN(n13706) );
  NAND4_X1 U7716 ( .A1(n13663), .A2(n13664), .A3(n13665), .A4(n13666), .ZN(
        n13653) );
  AOI221_X1 U7717 ( .B1(net227015), .B2(n16349), .C1(\registers[30][6] ), .C2(
        n16346), .A(n13668), .ZN(n13665) );
  AOI221_X1 U7718 ( .B1(\registers[10][6] ), .B2(n16325), .C1(
        \registers[0][6] ), .C2(n16322), .A(n13670), .ZN(n13663) );
  AOI221_X1 U7719 ( .B1(net227014), .B2(n16337), .C1(\registers[34][6] ), .C2(
        n16334), .A(n13669), .ZN(n13664) );
  NAND4_X1 U7720 ( .A1(n13621), .A2(n13622), .A3(n13623), .A4(n13624), .ZN(
        n13611) );
  AOI221_X1 U7721 ( .B1(net227033), .B2(n16349), .C1(\registers[30][7] ), .C2(
        n16346), .A(n13626), .ZN(n13623) );
  AOI221_X1 U7722 ( .B1(\registers[10][7] ), .B2(n16325), .C1(
        \registers[0][7] ), .C2(n16322), .A(n13628), .ZN(n13621) );
  AOI221_X1 U7723 ( .B1(net227032), .B2(n16337), .C1(\registers[34][7] ), .C2(
        n16334), .A(n13627), .ZN(n13622) );
  NAND4_X1 U7724 ( .A1(n13579), .A2(n13580), .A3(n13581), .A4(n13582), .ZN(
        n13569) );
  AOI221_X1 U7725 ( .B1(net227051), .B2(n16349), .C1(\registers[30][8] ), .C2(
        n16346), .A(n13584), .ZN(n13581) );
  AOI221_X1 U7726 ( .B1(\registers[10][8] ), .B2(n16325), .C1(
        \registers[0][8] ), .C2(n16322), .A(n13586), .ZN(n13579) );
  AOI221_X1 U7727 ( .B1(net227050), .B2(n16337), .C1(\registers[34][8] ), .C2(
        n16334), .A(n13585), .ZN(n13580) );
  NAND4_X1 U7728 ( .A1(n13537), .A2(n13538), .A3(n13539), .A4(n13540), .ZN(
        n13527) );
  AOI221_X1 U7729 ( .B1(net227069), .B2(n16349), .C1(\registers[30][9] ), .C2(
        n16346), .A(n13542), .ZN(n13539) );
  AOI221_X1 U7730 ( .B1(\registers[10][9] ), .B2(n16325), .C1(
        \registers[0][9] ), .C2(n16322), .A(n13544), .ZN(n13537) );
  AOI221_X1 U7731 ( .B1(net227068), .B2(n16337), .C1(\registers[34][9] ), .C2(
        n16334), .A(n13543), .ZN(n13538) );
  NAND4_X1 U7732 ( .A1(n13495), .A2(n13496), .A3(n13497), .A4(n13498), .ZN(
        n13485) );
  AOI221_X1 U7733 ( .B1(net227087), .B2(n16349), .C1(\registers[30][10] ), 
        .C2(n16346), .A(n13500), .ZN(n13497) );
  AOI221_X1 U7734 ( .B1(\registers[10][10] ), .B2(n16325), .C1(
        \registers[0][10] ), .C2(n16322), .A(n13502), .ZN(n13495) );
  AOI221_X1 U7735 ( .B1(net227086), .B2(n16337), .C1(\registers[34][10] ), 
        .C2(n16334), .A(n13501), .ZN(n13496) );
  NAND4_X1 U7736 ( .A1(n13453), .A2(n13454), .A3(n13455), .A4(n13456), .ZN(
        n13443) );
  AOI221_X1 U7737 ( .B1(net227105), .B2(n16349), .C1(\registers[30][11] ), 
        .C2(n16346), .A(n13458), .ZN(n13455) );
  AOI221_X1 U7738 ( .B1(\registers[10][11] ), .B2(n16325), .C1(
        \registers[0][11] ), .C2(n16322), .A(n13460), .ZN(n13453) );
  AOI221_X1 U7739 ( .B1(net227104), .B2(n16337), .C1(\registers[34][11] ), 
        .C2(n16334), .A(n13459), .ZN(n13454) );
  NAND4_X1 U7740 ( .A1(n13411), .A2(n13412), .A3(n13413), .A4(n13414), .ZN(
        n13401) );
  AOI221_X1 U7741 ( .B1(net227123), .B2(n16350), .C1(\registers[30][12] ), 
        .C2(n16347), .A(n13416), .ZN(n13413) );
  AOI221_X1 U7742 ( .B1(\registers[10][12] ), .B2(n16326), .C1(
        \registers[0][12] ), .C2(n16323), .A(n13418), .ZN(n13411) );
  AOI221_X1 U7743 ( .B1(net227122), .B2(n16338), .C1(\registers[34][12] ), 
        .C2(n16335), .A(n13417), .ZN(n13412) );
  NAND4_X1 U7744 ( .A1(n13369), .A2(n13370), .A3(n13371), .A4(n13372), .ZN(
        n13359) );
  AOI221_X1 U7745 ( .B1(net227141), .B2(n16350), .C1(\registers[30][13] ), 
        .C2(n16347), .A(n13374), .ZN(n13371) );
  AOI221_X1 U7746 ( .B1(\registers[10][13] ), .B2(n16326), .C1(
        \registers[0][13] ), .C2(n16323), .A(n13376), .ZN(n13369) );
  AOI221_X1 U7747 ( .B1(net227140), .B2(n16338), .C1(\registers[34][13] ), 
        .C2(n16335), .A(n13375), .ZN(n13370) );
  NAND4_X1 U7748 ( .A1(n13327), .A2(n13328), .A3(n13329), .A4(n13330), .ZN(
        n13317) );
  AOI221_X1 U7749 ( .B1(net227159), .B2(n16350), .C1(\registers[30][14] ), 
        .C2(n16347), .A(n13332), .ZN(n13329) );
  AOI221_X1 U7750 ( .B1(\registers[10][14] ), .B2(n16326), .C1(
        \registers[0][14] ), .C2(n16323), .A(n13334), .ZN(n13327) );
  AOI221_X1 U7751 ( .B1(net227158), .B2(n16338), .C1(\registers[34][14] ), 
        .C2(n16335), .A(n13333), .ZN(n13328) );
  NAND4_X1 U7752 ( .A1(n13285), .A2(n13286), .A3(n13287), .A4(n13288), .ZN(
        n13275) );
  AOI221_X1 U7753 ( .B1(net227177), .B2(n16350), .C1(\registers[30][15] ), 
        .C2(n16347), .A(n13290), .ZN(n13287) );
  AOI221_X1 U7754 ( .B1(\registers[10][15] ), .B2(n16326), .C1(
        \registers[0][15] ), .C2(n16323), .A(n13292), .ZN(n13285) );
  AOI221_X1 U7755 ( .B1(net227176), .B2(n16338), .C1(\registers[34][15] ), 
        .C2(n16335), .A(n13291), .ZN(n13286) );
  NAND4_X1 U7756 ( .A1(n13243), .A2(n13244), .A3(n13245), .A4(n13246), .ZN(
        n13233) );
  AOI221_X1 U7757 ( .B1(net227195), .B2(n16350), .C1(\registers[30][16] ), 
        .C2(n16347), .A(n13248), .ZN(n13245) );
  AOI221_X1 U7758 ( .B1(\registers[10][16] ), .B2(n16326), .C1(
        \registers[0][16] ), .C2(n16323), .A(n13250), .ZN(n13243) );
  AOI221_X1 U7759 ( .B1(net227194), .B2(n16338), .C1(\registers[34][16] ), 
        .C2(n16335), .A(n13249), .ZN(n13244) );
  NAND4_X1 U7760 ( .A1(n13201), .A2(n13202), .A3(n13203), .A4(n13204), .ZN(
        n13191) );
  AOI221_X1 U7761 ( .B1(net227213), .B2(n16350), .C1(\registers[30][17] ), 
        .C2(n16347), .A(n13206), .ZN(n13203) );
  AOI221_X1 U7762 ( .B1(\registers[10][17] ), .B2(n16326), .C1(
        \registers[0][17] ), .C2(n16323), .A(n13208), .ZN(n13201) );
  AOI221_X1 U7763 ( .B1(net227212), .B2(n16338), .C1(\registers[34][17] ), 
        .C2(n16335), .A(n13207), .ZN(n13202) );
  NAND4_X1 U7764 ( .A1(n13159), .A2(n13160), .A3(n13161), .A4(n13162), .ZN(
        n13149) );
  AOI221_X1 U7765 ( .B1(net227231), .B2(n16350), .C1(\registers[30][18] ), 
        .C2(n16347), .A(n13164), .ZN(n13161) );
  AOI221_X1 U7766 ( .B1(\registers[10][18] ), .B2(n16326), .C1(
        \registers[0][18] ), .C2(n16323), .A(n13166), .ZN(n13159) );
  AOI221_X1 U7767 ( .B1(net227230), .B2(n16338), .C1(\registers[34][18] ), 
        .C2(n16335), .A(n13165), .ZN(n13160) );
  NAND4_X1 U7768 ( .A1(n13117), .A2(n13118), .A3(n13119), .A4(n13120), .ZN(
        n13107) );
  AOI221_X1 U7769 ( .B1(net227249), .B2(n16350), .C1(\registers[30][19] ), 
        .C2(n16347), .A(n13122), .ZN(n13119) );
  AOI221_X1 U7770 ( .B1(\registers[10][19] ), .B2(n16326), .C1(
        \registers[0][19] ), .C2(n16323), .A(n13124), .ZN(n13117) );
  AOI221_X1 U7771 ( .B1(net227248), .B2(n16338), .C1(\registers[34][19] ), 
        .C2(n16335), .A(n13123), .ZN(n13118) );
  NAND4_X1 U7772 ( .A1(n13075), .A2(n13076), .A3(n13077), .A4(n13078), .ZN(
        n13065) );
  AOI221_X1 U7773 ( .B1(net227267), .B2(n16350), .C1(\registers[30][20] ), 
        .C2(n16347), .A(n13080), .ZN(n13077) );
  AOI221_X1 U7774 ( .B1(\registers[10][20] ), .B2(n16326), .C1(
        \registers[0][20] ), .C2(n16323), .A(n13082), .ZN(n13075) );
  AOI221_X1 U7775 ( .B1(net227266), .B2(n16338), .C1(\registers[34][20] ), 
        .C2(n16335), .A(n13081), .ZN(n13076) );
  NAND4_X1 U7776 ( .A1(n13033), .A2(n13034), .A3(n13035), .A4(n13036), .ZN(
        n13023) );
  AOI221_X1 U7777 ( .B1(net227285), .B2(n16350), .C1(\registers[30][21] ), 
        .C2(n16347), .A(n13038), .ZN(n13035) );
  AOI221_X1 U7778 ( .B1(\registers[10][21] ), .B2(n16326), .C1(
        \registers[0][21] ), .C2(n16323), .A(n13040), .ZN(n13033) );
  AOI221_X1 U7779 ( .B1(net227284), .B2(n16338), .C1(\registers[34][21] ), 
        .C2(n16335), .A(n13039), .ZN(n13034) );
  NAND4_X1 U7780 ( .A1(n12991), .A2(n12992), .A3(n12993), .A4(n12994), .ZN(
        n12981) );
  AOI221_X1 U7781 ( .B1(net227303), .B2(n16350), .C1(\registers[30][22] ), 
        .C2(n16347), .A(n12996), .ZN(n12993) );
  AOI221_X1 U7782 ( .B1(\registers[10][22] ), .B2(n16326), .C1(
        \registers[0][22] ), .C2(n16323), .A(n12998), .ZN(n12991) );
  AOI221_X1 U7783 ( .B1(net227302), .B2(n16338), .C1(\registers[34][22] ), 
        .C2(n16335), .A(n12997), .ZN(n12992) );
  NAND4_X1 U7784 ( .A1(n12949), .A2(n12950), .A3(n12951), .A4(n12952), .ZN(
        n12939) );
  AOI221_X1 U7785 ( .B1(net227321), .B2(n16350), .C1(\registers[30][23] ), 
        .C2(n16347), .A(n12954), .ZN(n12951) );
  AOI221_X1 U7786 ( .B1(\registers[10][23] ), .B2(n16326), .C1(
        \registers[0][23] ), .C2(n16323), .A(n12956), .ZN(n12949) );
  AOI221_X1 U7787 ( .B1(net227320), .B2(n16338), .C1(\registers[34][23] ), 
        .C2(n16335), .A(n12955), .ZN(n12950) );
  NAND4_X1 U7788 ( .A1(n12457), .A2(n12458), .A3(n12459), .A4(n12460), .ZN(
        n12429) );
  AOI221_X1 U7789 ( .B1(net226848), .B2(n16601), .C1(\registers[30][0] ), .C2(
        n16598), .A(n12462), .ZN(n12459) );
  AOI221_X1 U7790 ( .B1(\registers[10][0] ), .B2(n16577), .C1(
        \registers[0][0] ), .C2(n16574), .A(n12466), .ZN(n12457) );
  AOI221_X1 U7791 ( .B1(net226847), .B2(n16589), .C1(\registers[34][0] ), .C2(
        n16586), .A(n12464), .ZN(n12458) );
  NAND4_X1 U7792 ( .A1(n12277), .A2(n12278), .A3(n12279), .A4(n12280), .ZN(
        n12267) );
  AOI221_X1 U7793 ( .B1(net226869), .B2(n16601), .C1(\registers[30][1] ), .C2(
        n16598), .A(n12282), .ZN(n12279) );
  AOI221_X1 U7794 ( .B1(\registers[10][1] ), .B2(n16577), .C1(
        \registers[0][1] ), .C2(n16574), .A(n12284), .ZN(n12277) );
  AOI221_X1 U7795 ( .B1(net226868), .B2(n16589), .C1(\registers[34][1] ), .C2(
        n16586), .A(n12283), .ZN(n12278) );
  NAND4_X1 U7796 ( .A1(n12124), .A2(n12125), .A3(n12126), .A4(n12127), .ZN(
        n12114) );
  AOI221_X1 U7797 ( .B1(net226888), .B2(n16601), .C1(\registers[30][2] ), .C2(
        n16598), .A(n12129), .ZN(n12126) );
  AOI221_X1 U7798 ( .B1(\registers[10][2] ), .B2(n16577), .C1(
        \registers[0][2] ), .C2(n16574), .A(n12131), .ZN(n12124) );
  AOI221_X1 U7799 ( .B1(net226880), .B2(n16589), .C1(\registers[34][2] ), .C2(
        n16586), .A(n12130), .ZN(n12125) );
  NAND4_X1 U7800 ( .A1(n11971), .A2(n11972), .A3(n11973), .A4(n11974), .ZN(
        n11961) );
  AOI221_X1 U7801 ( .B1(net226908), .B2(n16601), .C1(\registers[30][3] ), .C2(
        n16598), .A(n11976), .ZN(n11973) );
  AOI221_X1 U7802 ( .B1(\registers[10][3] ), .B2(n16577), .C1(
        \registers[0][3] ), .C2(n16574), .A(n11978), .ZN(n11971) );
  AOI221_X1 U7803 ( .B1(net226900), .B2(n16589), .C1(\registers[34][3] ), .C2(
        n16586), .A(n11977), .ZN(n11972) );
  NAND4_X1 U7804 ( .A1(n11818), .A2(n11819), .A3(n11820), .A4(n11821), .ZN(
        n11808) );
  AOI221_X1 U7805 ( .B1(net226982), .B2(n16601), .C1(\registers[30][4] ), .C2(
        n16598), .A(n11823), .ZN(n11820) );
  AOI221_X1 U7806 ( .B1(\registers[10][4] ), .B2(n16577), .C1(
        \registers[0][4] ), .C2(n16574), .A(n11825), .ZN(n11818) );
  AOI221_X1 U7807 ( .B1(net226973), .B2(n16589), .C1(\registers[34][4] ), .C2(
        n16586), .A(n11824), .ZN(n11819) );
  NAND4_X1 U7808 ( .A1(n11775), .A2(n11776), .A3(n11777), .A4(n11778), .ZN(
        n11765) );
  AOI221_X1 U7809 ( .B1(net226991), .B2(n16601), .C1(\registers[30][5] ), .C2(
        n16598), .A(n11780), .ZN(n11777) );
  AOI221_X1 U7810 ( .B1(\registers[10][5] ), .B2(n16577), .C1(
        \registers[0][5] ), .C2(n16574), .A(n11782), .ZN(n11775) );
  AOI221_X1 U7811 ( .B1(net226990), .B2(n16589), .C1(\registers[34][5] ), .C2(
        n16586), .A(n11781), .ZN(n11776) );
  NAND4_X1 U7812 ( .A1(n11732), .A2(n11733), .A3(n11734), .A4(n11735), .ZN(
        n11722) );
  AOI221_X1 U7813 ( .B1(net227015), .B2(n16601), .C1(\registers[30][6] ), .C2(
        n16598), .A(n11737), .ZN(n11734) );
  AOI221_X1 U7814 ( .B1(\registers[10][6] ), .B2(n16577), .C1(
        \registers[0][6] ), .C2(n16574), .A(n11739), .ZN(n11732) );
  AOI221_X1 U7815 ( .B1(net227014), .B2(n16589), .C1(\registers[34][6] ), .C2(
        n16586), .A(n11738), .ZN(n11733) );
  NAND4_X1 U7816 ( .A1(n11689), .A2(n11690), .A3(n11691), .A4(n11692), .ZN(
        n11679) );
  AOI221_X1 U7817 ( .B1(net227033), .B2(n16601), .C1(\registers[30][7] ), .C2(
        n16598), .A(n11694), .ZN(n11691) );
  AOI221_X1 U7818 ( .B1(\registers[10][7] ), .B2(n16577), .C1(
        \registers[0][7] ), .C2(n16574), .A(n11696), .ZN(n11689) );
  AOI221_X1 U7819 ( .B1(net227032), .B2(n16589), .C1(\registers[34][7] ), .C2(
        n16586), .A(n11695), .ZN(n11690) );
  NAND4_X1 U7820 ( .A1(n11646), .A2(n11647), .A3(n11648), .A4(n11649), .ZN(
        n11636) );
  AOI221_X1 U7821 ( .B1(net227051), .B2(n16601), .C1(\registers[30][8] ), .C2(
        n16598), .A(n11651), .ZN(n11648) );
  AOI221_X1 U7822 ( .B1(\registers[10][8] ), .B2(n16577), .C1(
        \registers[0][8] ), .C2(n16574), .A(n11653), .ZN(n11646) );
  AOI221_X1 U7823 ( .B1(net227050), .B2(n16589), .C1(\registers[34][8] ), .C2(
        n16586), .A(n11652), .ZN(n11647) );
  NAND4_X1 U7824 ( .A1(n11603), .A2(n11604), .A3(n11605), .A4(n11606), .ZN(
        n11593) );
  AOI221_X1 U7825 ( .B1(net227069), .B2(n16601), .C1(\registers[30][9] ), .C2(
        n16598), .A(n11608), .ZN(n11605) );
  AOI221_X1 U7826 ( .B1(\registers[10][9] ), .B2(n16577), .C1(
        \registers[0][9] ), .C2(n16574), .A(n11610), .ZN(n11603) );
  AOI221_X1 U7827 ( .B1(net227068), .B2(n16589), .C1(\registers[34][9] ), .C2(
        n16586), .A(n11609), .ZN(n11604) );
  NAND4_X1 U7828 ( .A1(n11560), .A2(n11561), .A3(n11562), .A4(n11563), .ZN(
        n11550) );
  AOI221_X1 U7829 ( .B1(net227087), .B2(n16601), .C1(\registers[30][10] ), 
        .C2(n16598), .A(n11565), .ZN(n11562) );
  AOI221_X1 U7830 ( .B1(\registers[10][10] ), .B2(n16577), .C1(
        \registers[0][10] ), .C2(n16574), .A(n11567), .ZN(n11560) );
  AOI221_X1 U7831 ( .B1(net227086), .B2(n16589), .C1(\registers[34][10] ), 
        .C2(n16586), .A(n11566), .ZN(n11561) );
  NAND4_X1 U7832 ( .A1(n11517), .A2(n11518), .A3(n11519), .A4(n11520), .ZN(
        n11507) );
  AOI221_X1 U7833 ( .B1(net227105), .B2(n16601), .C1(\registers[30][11] ), 
        .C2(n16598), .A(n11522), .ZN(n11519) );
  AOI221_X1 U7834 ( .B1(\registers[10][11] ), .B2(n16577), .C1(
        \registers[0][11] ), .C2(n16574), .A(n11524), .ZN(n11517) );
  AOI221_X1 U7835 ( .B1(net227104), .B2(n16589), .C1(\registers[34][11] ), 
        .C2(n16586), .A(n11523), .ZN(n11518) );
  NAND4_X1 U7836 ( .A1(n11474), .A2(n11475), .A3(n11476), .A4(n11477), .ZN(
        n11464) );
  AOI221_X1 U7837 ( .B1(net227123), .B2(n16602), .C1(\registers[30][12] ), 
        .C2(n16599), .A(n11479), .ZN(n11476) );
  AOI221_X1 U7838 ( .B1(\registers[10][12] ), .B2(n16578), .C1(
        \registers[0][12] ), .C2(n16575), .A(n11481), .ZN(n11474) );
  AOI221_X1 U7839 ( .B1(net227122), .B2(n16590), .C1(\registers[34][12] ), 
        .C2(n16587), .A(n11480), .ZN(n11475) );
  NAND4_X1 U7840 ( .A1(n11430), .A2(n11431), .A3(n11432), .A4(n11433), .ZN(
        n11420) );
  AOI221_X1 U7841 ( .B1(net227141), .B2(n16602), .C1(\registers[30][13] ), 
        .C2(n16599), .A(n11435), .ZN(n11432) );
  AOI221_X1 U7842 ( .B1(\registers[10][13] ), .B2(n16578), .C1(
        \registers[0][13] ), .C2(n16575), .A(n11437), .ZN(n11430) );
  AOI221_X1 U7843 ( .B1(net227140), .B2(n16590), .C1(\registers[34][13] ), 
        .C2(n16587), .A(n11436), .ZN(n11431) );
  NAND4_X1 U7844 ( .A1(n11387), .A2(n11388), .A3(n11389), .A4(n11390), .ZN(
        n11377) );
  AOI221_X1 U7845 ( .B1(net227159), .B2(n16602), .C1(\registers[30][14] ), 
        .C2(n16599), .A(n11392), .ZN(n11389) );
  AOI221_X1 U7846 ( .B1(\registers[10][14] ), .B2(n16578), .C1(
        \registers[0][14] ), .C2(n16575), .A(n11394), .ZN(n11387) );
  AOI221_X1 U7847 ( .B1(net227158), .B2(n16590), .C1(\registers[34][14] ), 
        .C2(n16587), .A(n11393), .ZN(n11388) );
  NAND4_X1 U7848 ( .A1(n11344), .A2(n11345), .A3(n11346), .A4(n11347), .ZN(
        n11334) );
  AOI221_X1 U7849 ( .B1(net227177), .B2(n16602), .C1(\registers[30][15] ), 
        .C2(n16599), .A(n11349), .ZN(n11346) );
  AOI221_X1 U7850 ( .B1(\registers[10][15] ), .B2(n16578), .C1(
        \registers[0][15] ), .C2(n16575), .A(n11351), .ZN(n11344) );
  AOI221_X1 U7851 ( .B1(net227176), .B2(n16590), .C1(\registers[34][15] ), 
        .C2(n16587), .A(n11350), .ZN(n11345) );
  NAND4_X1 U7852 ( .A1(n11301), .A2(n11302), .A3(n11303), .A4(n11304), .ZN(
        n11291) );
  AOI221_X1 U7853 ( .B1(net227195), .B2(n16602), .C1(\registers[30][16] ), 
        .C2(n16599), .A(n11306), .ZN(n11303) );
  AOI221_X1 U7854 ( .B1(\registers[10][16] ), .B2(n16578), .C1(
        \registers[0][16] ), .C2(n16575), .A(n11308), .ZN(n11301) );
  AOI221_X1 U7855 ( .B1(net227194), .B2(n16590), .C1(\registers[34][16] ), 
        .C2(n16587), .A(n11307), .ZN(n11302) );
  NAND4_X1 U7856 ( .A1(n11258), .A2(n11259), .A3(n11260), .A4(n11261), .ZN(
        n11248) );
  AOI221_X1 U7857 ( .B1(net227213), .B2(n16602), .C1(\registers[30][17] ), 
        .C2(n16599), .A(n11263), .ZN(n11260) );
  AOI221_X1 U7858 ( .B1(\registers[10][17] ), .B2(n16578), .C1(
        \registers[0][17] ), .C2(n16575), .A(n11265), .ZN(n11258) );
  AOI221_X1 U7859 ( .B1(net227212), .B2(n16590), .C1(\registers[34][17] ), 
        .C2(n16587), .A(n11264), .ZN(n11259) );
  NAND4_X1 U7860 ( .A1(n11215), .A2(n11216), .A3(n11217), .A4(n11218), .ZN(
        n11205) );
  AOI221_X1 U7861 ( .B1(net227231), .B2(n16602), .C1(\registers[30][18] ), 
        .C2(n16599), .A(n11220), .ZN(n11217) );
  AOI221_X1 U7862 ( .B1(\registers[10][18] ), .B2(n16578), .C1(
        \registers[0][18] ), .C2(n16575), .A(n11222), .ZN(n11215) );
  AOI221_X1 U7863 ( .B1(net227230), .B2(n16590), .C1(\registers[34][18] ), 
        .C2(n16587), .A(n11221), .ZN(n11216) );
  NAND4_X1 U7864 ( .A1(n11172), .A2(n11173), .A3(n11174), .A4(n11175), .ZN(
        n11162) );
  AOI221_X1 U7865 ( .B1(net227249), .B2(n16602), .C1(\registers[30][19] ), 
        .C2(n16599), .A(n11177), .ZN(n11174) );
  AOI221_X1 U7866 ( .B1(\registers[10][19] ), .B2(n16578), .C1(
        \registers[0][19] ), .C2(n16575), .A(n11179), .ZN(n11172) );
  AOI221_X1 U7867 ( .B1(net227248), .B2(n16590), .C1(\registers[34][19] ), 
        .C2(n16587), .A(n11178), .ZN(n11173) );
  NAND4_X1 U7868 ( .A1(n11129), .A2(n11130), .A3(n11131), .A4(n11132), .ZN(
        n11119) );
  AOI221_X1 U7869 ( .B1(net227267), .B2(n16602), .C1(\registers[30][20] ), 
        .C2(n16599), .A(n11134), .ZN(n11131) );
  AOI221_X1 U7870 ( .B1(\registers[10][20] ), .B2(n16578), .C1(
        \registers[0][20] ), .C2(n16575), .A(n11136), .ZN(n11129) );
  AOI221_X1 U7871 ( .B1(net227266), .B2(n16590), .C1(\registers[34][20] ), 
        .C2(n16587), .A(n11135), .ZN(n11130) );
  NAND4_X1 U7872 ( .A1(n11086), .A2(n11087), .A3(n11088), .A4(n11089), .ZN(
        n11076) );
  AOI221_X1 U7873 ( .B1(net227285), .B2(n16602), .C1(\registers[30][21] ), 
        .C2(n16599), .A(n11091), .ZN(n11088) );
  AOI221_X1 U7874 ( .B1(\registers[10][21] ), .B2(n16578), .C1(
        \registers[0][21] ), .C2(n16575), .A(n11093), .ZN(n11086) );
  AOI221_X1 U7875 ( .B1(net227284), .B2(n16590), .C1(\registers[34][21] ), 
        .C2(n16587), .A(n11092), .ZN(n11087) );
  NAND4_X1 U7876 ( .A1(n11043), .A2(n11044), .A3(n11045), .A4(n11046), .ZN(
        n11033) );
  AOI221_X1 U7877 ( .B1(net227303), .B2(n16602), .C1(\registers[30][22] ), 
        .C2(n16599), .A(n11048), .ZN(n11045) );
  AOI221_X1 U7878 ( .B1(\registers[10][22] ), .B2(n16578), .C1(
        \registers[0][22] ), .C2(n16575), .A(n11050), .ZN(n11043) );
  AOI221_X1 U7879 ( .B1(net227302), .B2(n16590), .C1(\registers[34][22] ), 
        .C2(n16587), .A(n11049), .ZN(n11044) );
  NAND4_X1 U7880 ( .A1(n11000), .A2(n11001), .A3(n11002), .A4(n11003), .ZN(
        n10990) );
  AOI221_X1 U7881 ( .B1(net227321), .B2(n16602), .C1(\registers[30][23] ), 
        .C2(n16599), .A(n11005), .ZN(n11002) );
  AOI221_X1 U7882 ( .B1(\registers[10][23] ), .B2(n16578), .C1(
        \registers[0][23] ), .C2(n16575), .A(n11007), .ZN(n11000) );
  AOI221_X1 U7883 ( .B1(net227320), .B2(n16590), .C1(\registers[34][23] ), 
        .C2(n16587), .A(n11006), .ZN(n11001) );
  NAND4_X1 U7884 ( .A1(n12383), .A2(n12384), .A3(n12385), .A4(n12386), .ZN(
        n12373) );
  AOI221_X1 U7885 ( .B1(net226840), .B2(n17757), .C1(\registers[25][0] ), .C2(
        n17754), .A(n12388), .ZN(n12385) );
  AOI221_X1 U7886 ( .B1(net226837), .B2(n17769), .C1(\registers[50][0] ), .C2(
        n17766), .A(n12387), .ZN(n12386) );
  AOI221_X1 U7887 ( .B1(\registers[36][0] ), .B2(n17733), .C1(
        \registers[38][0] ), .C2(n17730), .A(n12390), .ZN(n12383) );
  NAND4_X1 U7888 ( .A1(n12229), .A2(n12230), .A3(n12231), .A4(n12232), .ZN(
        n12219) );
  AOI221_X1 U7889 ( .B1(net226862), .B2(n17757), .C1(\registers[25][1] ), .C2(
        n17754), .A(n12234), .ZN(n12231) );
  AOI221_X1 U7890 ( .B1(net226860), .B2(n17769), .C1(\registers[50][1] ), .C2(
        n17766), .A(n12233), .ZN(n12232) );
  AOI221_X1 U7891 ( .B1(\registers[36][1] ), .B2(n17733), .C1(
        \registers[38][1] ), .C2(n17730), .A(n12236), .ZN(n12229) );
  NAND4_X1 U7892 ( .A1(n12074), .A2(n12075), .A3(n12076), .A4(n12077), .ZN(
        n12064) );
  AOI221_X1 U7893 ( .B1(net226881), .B2(n17757), .C1(\registers[25][2] ), .C2(
        n17754), .A(n12079), .ZN(n12076) );
  AOI221_X1 U7894 ( .B1(net226886), .B2(n17769), .C1(\registers[50][2] ), .C2(
        n17766), .A(n12078), .ZN(n12077) );
  AOI221_X1 U7895 ( .B1(\registers[36][2] ), .B2(n17733), .C1(
        \registers[38][2] ), .C2(n17730), .A(n12081), .ZN(n12074) );
  NAND4_X1 U7896 ( .A1(n11921), .A2(n11922), .A3(n11923), .A4(n11924), .ZN(
        n11911) );
  AOI221_X1 U7897 ( .B1(net226910), .B2(n17757), .C1(\registers[25][3] ), .C2(
        n17754), .A(n11926), .ZN(n11923) );
  AOI221_X1 U7898 ( .B1(net226899), .B2(n17769), .C1(\registers[50][3] ), .C2(
        n17766), .A(n11925), .ZN(n11924) );
  AOI221_X1 U7899 ( .B1(\registers[36][3] ), .B2(n17733), .C1(
        \registers[38][3] ), .C2(n17730), .A(n11928), .ZN(n11921) );
  NAND4_X1 U7900 ( .A1(n10478), .A2(n10479), .A3(n10480), .A4(n10481), .ZN(
        n10468) );
  AOI221_X1 U7901 ( .B1(net226984), .B2(n17757), .C1(\registers[25][4] ), .C2(
        n17754), .A(n10483), .ZN(n10480) );
  AOI221_X1 U7902 ( .B1(net226981), .B2(n17769), .C1(\registers[50][4] ), .C2(
        n17766), .A(n10482), .ZN(n10481) );
  AOI221_X1 U7903 ( .B1(\registers[36][4] ), .B2(n17733), .C1(
        \registers[38][4] ), .C2(n17730), .A(n10485), .ZN(n10478) );
  NAND4_X1 U7904 ( .A1(n10368), .A2(n10369), .A3(n10370), .A4(n10371), .ZN(
        n10358) );
  AOI221_X1 U7905 ( .B1(net226993), .B2(n17757), .C1(\registers[25][5] ), .C2(
        n17754), .A(n10373), .ZN(n10370) );
  AOI221_X1 U7906 ( .B1(net227001), .B2(n17769), .C1(\registers[50][5] ), .C2(
        n17766), .A(n10372), .ZN(n10371) );
  AOI221_X1 U7907 ( .B1(\registers[36][5] ), .B2(n17733), .C1(
        \registers[38][5] ), .C2(n17730), .A(n10375), .ZN(n10368) );
  NAND4_X1 U7908 ( .A1(n10256), .A2(n10257), .A3(n10258), .A4(n10259), .ZN(
        n10246) );
  AOI221_X1 U7909 ( .B1(net227017), .B2(n17757), .C1(\registers[25][6] ), .C2(
        n17754), .A(n10261), .ZN(n10258) );
  AOI221_X1 U7910 ( .B1(net227012), .B2(n17769), .C1(\registers[50][6] ), .C2(
        n17766), .A(n10260), .ZN(n10259) );
  AOI221_X1 U7911 ( .B1(\registers[36][6] ), .B2(n17733), .C1(
        \registers[38][6] ), .C2(n17730), .A(n10263), .ZN(n10256) );
  NAND4_X1 U7912 ( .A1(n7620), .A2(n7621), .A3(n7622), .A4(n7623), .ZN(n7610)
         );
  AOI221_X1 U7913 ( .B1(net227035), .B2(n17757), .C1(\registers[25][7] ), .C2(
        n17754), .A(n7625), .ZN(n7622) );
  AOI221_X1 U7914 ( .B1(net227030), .B2(n17769), .C1(\registers[50][7] ), .C2(
        n17766), .A(n7624), .ZN(n7623) );
  AOI221_X1 U7915 ( .B1(\registers[36][7] ), .B2(n17733), .C1(
        \registers[38][7] ), .C2(n17730), .A(n7627), .ZN(n7620) );
  NAND4_X1 U7916 ( .A1(n7505), .A2(n7506), .A3(n7507), .A4(n7508), .ZN(n7495)
         );
  AOI221_X1 U7917 ( .B1(net227053), .B2(n17757), .C1(\registers[25][8] ), .C2(
        n17754), .A(n7510), .ZN(n7507) );
  AOI221_X1 U7918 ( .B1(net227048), .B2(n17769), .C1(\registers[50][8] ), .C2(
        n17766), .A(n7509), .ZN(n7508) );
  AOI221_X1 U7919 ( .B1(\registers[36][8] ), .B2(n17733), .C1(
        \registers[38][8] ), .C2(n17730), .A(n7512), .ZN(n7505) );
  NAND4_X1 U7920 ( .A1(n7396), .A2(n7397), .A3(n7398), .A4(n7399), .ZN(n7386)
         );
  AOI221_X1 U7921 ( .B1(net227071), .B2(n17757), .C1(\registers[25][9] ), .C2(
        n17754), .A(n7401), .ZN(n7398) );
  AOI221_X1 U7922 ( .B1(net227066), .B2(n17769), .C1(\registers[50][9] ), .C2(
        n17766), .A(n7400), .ZN(n7399) );
  AOI221_X1 U7923 ( .B1(\registers[36][9] ), .B2(n17733), .C1(
        \registers[38][9] ), .C2(n17730), .A(n7403), .ZN(n7396) );
  NAND4_X1 U7924 ( .A1(n7287), .A2(n7288), .A3(n7289), .A4(n7290), .ZN(n7277)
         );
  AOI221_X1 U7925 ( .B1(net227089), .B2(n17757), .C1(\registers[25][10] ), 
        .C2(n17754), .A(n7292), .ZN(n7289) );
  AOI221_X1 U7926 ( .B1(net227084), .B2(n17769), .C1(\registers[50][10] ), 
        .C2(n17766), .A(n7291), .ZN(n7290) );
  AOI221_X1 U7927 ( .B1(\registers[36][10] ), .B2(n17733), .C1(
        \registers[38][10] ), .C2(n17730), .A(n7294), .ZN(n7287) );
  NAND4_X1 U7928 ( .A1(n7173), .A2(n7174), .A3(n7175), .A4(n7176), .ZN(n7163)
         );
  AOI221_X1 U7929 ( .B1(net227107), .B2(n17758), .C1(\registers[25][11] ), 
        .C2(n17755), .A(n7178), .ZN(n7175) );
  AOI221_X1 U7930 ( .B1(net227102), .B2(n17770), .C1(\registers[50][11] ), 
        .C2(n17767), .A(n7177), .ZN(n7176) );
  AOI221_X1 U7931 ( .B1(\registers[36][11] ), .B2(n17734), .C1(
        \registers[38][11] ), .C2(n17731), .A(n7180), .ZN(n7173) );
  NAND4_X1 U7932 ( .A1(n7064), .A2(n7065), .A3(n7066), .A4(n7067), .ZN(n7054)
         );
  AOI221_X1 U7933 ( .B1(net227125), .B2(n17758), .C1(\registers[25][12] ), 
        .C2(n17755), .A(n7069), .ZN(n7066) );
  AOI221_X1 U7934 ( .B1(net227120), .B2(n17770), .C1(\registers[50][12] ), 
        .C2(n17767), .A(n7068), .ZN(n7067) );
  AOI221_X1 U7935 ( .B1(\registers[36][12] ), .B2(n17734), .C1(
        \registers[38][12] ), .C2(n17731), .A(n7071), .ZN(n7064) );
  NAND4_X1 U7936 ( .A1(n6955), .A2(n6956), .A3(n6957), .A4(n6958), .ZN(n6945)
         );
  AOI221_X1 U7937 ( .B1(net227143), .B2(n17758), .C1(\registers[25][13] ), 
        .C2(n17755), .A(n6960), .ZN(n6957) );
  AOI221_X1 U7938 ( .B1(net227138), .B2(n17770), .C1(\registers[50][13] ), 
        .C2(n17767), .A(n6959), .ZN(n6958) );
  AOI221_X1 U7939 ( .B1(\registers[36][13] ), .B2(n17734), .C1(
        \registers[38][13] ), .C2(n17731), .A(n6962), .ZN(n6955) );
  NAND4_X1 U7940 ( .A1(n6846), .A2(n6847), .A3(n6848), .A4(n6849), .ZN(n6836)
         );
  AOI221_X1 U7941 ( .B1(net227161), .B2(n17758), .C1(\registers[25][14] ), 
        .C2(n17755), .A(n6851), .ZN(n6848) );
  AOI221_X1 U7942 ( .B1(net227156), .B2(n17770), .C1(\registers[50][14] ), 
        .C2(n17767), .A(n6850), .ZN(n6849) );
  AOI221_X1 U7943 ( .B1(\registers[36][14] ), .B2(n17734), .C1(
        \registers[38][14] ), .C2(n17731), .A(n6853), .ZN(n6846) );
  NAND4_X1 U7944 ( .A1(n6737), .A2(n6738), .A3(n6739), .A4(n6740), .ZN(n6727)
         );
  AOI221_X1 U7945 ( .B1(net227179), .B2(n17758), .C1(\registers[25][15] ), 
        .C2(n17755), .A(n6742), .ZN(n6739) );
  AOI221_X1 U7946 ( .B1(net227174), .B2(n17770), .C1(\registers[50][15] ), 
        .C2(n17767), .A(n6741), .ZN(n6740) );
  AOI221_X1 U7947 ( .B1(\registers[36][15] ), .B2(n17734), .C1(
        \registers[38][15] ), .C2(n17731), .A(n6744), .ZN(n6737) );
  NAND4_X1 U7948 ( .A1(n6577), .A2(n6580), .A3(n6581), .A4(n6582), .ZN(n6564)
         );
  AOI221_X1 U7949 ( .B1(net227197), .B2(n17758), .C1(\registers[25][16] ), 
        .C2(n17755), .A(n6599), .ZN(n6581) );
  AOI221_X1 U7950 ( .B1(net227192), .B2(n17770), .C1(\registers[50][16] ), 
        .C2(n17767), .A(n6598), .ZN(n6582) );
  AOI221_X1 U7951 ( .B1(\registers[36][16] ), .B2(n17734), .C1(
        \registers[38][16] ), .C2(n17731), .A(n6601), .ZN(n6577) );
  NAND4_X1 U7952 ( .A1(n6392), .A2(n6393), .A3(n6409), .A4(n6410), .ZN(n6377)
         );
  AOI221_X1 U7953 ( .B1(net227215), .B2(n17758), .C1(\registers[25][17] ), 
        .C2(n17755), .A(n6412), .ZN(n6409) );
  AOI221_X1 U7954 ( .B1(net227210), .B2(n17770), .C1(\registers[50][17] ), 
        .C2(n17767), .A(n6411), .ZN(n6410) );
  AOI221_X1 U7955 ( .B1(\registers[36][17] ), .B2(n17734), .C1(
        \registers[38][17] ), .C2(n17731), .A(n6414), .ZN(n6392) );
  NAND4_X1 U7956 ( .A1(n6220), .A2(n6221), .A3(n6222), .A4(n6223), .ZN(n6192)
         );
  AOI221_X1 U7957 ( .B1(net227233), .B2(n17758), .C1(\registers[25][18] ), 
        .C2(n17755), .A(n6225), .ZN(n6222) );
  AOI221_X1 U7958 ( .B1(net227228), .B2(n17770), .C1(\registers[50][18] ), 
        .C2(n17767), .A(n6224), .ZN(n6223) );
  AOI221_X1 U7959 ( .B1(\registers[36][18] ), .B2(n17734), .C1(
        \registers[38][18] ), .C2(n17731), .A(n6227), .ZN(n6220) );
  NAND4_X1 U7960 ( .A1(n6033), .A2(n6034), .A3(n6035), .A4(n6036), .ZN(n6006)
         );
  AOI221_X1 U7961 ( .B1(net227251), .B2(n17758), .C1(\registers[25][19] ), 
        .C2(n17755), .A(n6038), .ZN(n6035) );
  AOI221_X1 U7962 ( .B1(net227246), .B2(n17770), .C1(\registers[50][19] ), 
        .C2(n17767), .A(n6037), .ZN(n6036) );
  AOI221_X1 U7963 ( .B1(\registers[36][19] ), .B2(n17734), .C1(
        \registers[38][19] ), .C2(n17731), .A(n6040), .ZN(n6033) );
  NAND4_X1 U7964 ( .A1(n5846), .A2(n5847), .A3(n5848), .A4(n5849), .ZN(n5819)
         );
  AOI221_X1 U7965 ( .B1(net227269), .B2(n17758), .C1(\registers[25][20] ), 
        .C2(n17755), .A(n5851), .ZN(n5848) );
  AOI221_X1 U7966 ( .B1(net227264), .B2(n17770), .C1(\registers[50][20] ), 
        .C2(n17767), .A(n5850), .ZN(n5849) );
  AOI221_X1 U7967 ( .B1(\registers[36][20] ), .B2(n17734), .C1(
        \registers[38][20] ), .C2(n17731), .A(n5854), .ZN(n5846) );
  NAND4_X1 U7968 ( .A1(n5659), .A2(n5660), .A3(n5661), .A4(n5662), .ZN(n5632)
         );
  AOI221_X1 U7969 ( .B1(net227287), .B2(n17758), .C1(\registers[25][21] ), 
        .C2(n17755), .A(n5665), .ZN(n5661) );
  AOI221_X1 U7970 ( .B1(net227282), .B2(n17770), .C1(\registers[50][21] ), 
        .C2(n17767), .A(n5664), .ZN(n5662) );
  AOI221_X1 U7971 ( .B1(\registers[36][21] ), .B2(n17734), .C1(
        \registers[38][21] ), .C2(n17731), .A(n5669), .ZN(n5659) );
  NAND4_X1 U7972 ( .A1(n5472), .A2(n5473), .A3(n5475), .A4(n5476), .ZN(n5447)
         );
  AOI221_X1 U7973 ( .B1(net227305), .B2(n17758), .C1(\registers[25][22] ), 
        .C2(n17755), .A(n5480), .ZN(n5475) );
  AOI221_X1 U7974 ( .B1(net227300), .B2(n17770), .C1(\registers[50][22] ), 
        .C2(n17767), .A(n5478), .ZN(n5476) );
  AOI221_X1 U7975 ( .B1(\registers[36][22] ), .B2(n17734), .C1(
        \registers[38][22] ), .C2(n17731), .A(n5482), .ZN(n5472) );
  NAND4_X1 U7976 ( .A1(n14109), .A2(n14110), .A3(n14111), .A4(n14112), .ZN(
        n14078) );
  AOI221_X1 U7977 ( .B1(net227467), .B2(n17757), .C1(\registers[25][31] ), 
        .C2(n17754), .A(n14126), .ZN(n14111) );
  AOI221_X1 U7978 ( .B1(net227462), .B2(n17769), .C1(\registers[50][31] ), 
        .C2(n17766), .A(n14113), .ZN(n14112) );
  AOI221_X1 U7979 ( .B1(\registers[36][31] ), .B2(n17733), .C1(
        \registers[38][31] ), .C2(n17730), .A(n14148), .ZN(n14109) );
  NAND2_X1 U7980 ( .A1(n14129), .A2(call), .ZN(n14115) );
  NAND4_X1 U7981 ( .A1(n5298), .A2(n5299), .A3(n5301), .A4(n5302), .ZN(n5274)
         );
  AOI221_X1 U7982 ( .B1(net227316), .B2(n17711), .C1(net227315), .C2(n17708), 
        .A(n5304), .ZN(n5301) );
  AOI221_X1 U7983 ( .B1(net227317), .B2(n17723), .C1(\registers[54][23] ), 
        .C2(n17720), .A(n5303), .ZN(n5302) );
  AOI221_X1 U7984 ( .B1(\registers[42][23] ), .B2(n17687), .C1(
        \registers[43][23] ), .C2(n17684), .A(n5307), .ZN(n5298) );
  NAND4_X1 U7985 ( .A1(n5130), .A2(n5131), .A3(n5132), .A4(n5133), .ZN(n5108)
         );
  AOI221_X1 U7986 ( .B1(net227334), .B2(n17711), .C1(net227333), .C2(n17708), 
        .A(n5135), .ZN(n5132) );
  AOI221_X1 U7987 ( .B1(net227335), .B2(n17723), .C1(\registers[54][24] ), 
        .C2(n17720), .A(n5134), .ZN(n5133) );
  AOI221_X1 U7988 ( .B1(\registers[42][24] ), .B2(n17687), .C1(
        \registers[43][24] ), .C2(n17684), .A(n5137), .ZN(n5130) );
  NAND4_X1 U7989 ( .A1(n5014), .A2(n5015), .A3(n5016), .A4(n5017), .ZN(n4995)
         );
  AOI221_X1 U7990 ( .B1(net227352), .B2(n17711), .C1(net227351), .C2(n17708), 
        .A(n5021), .ZN(n5016) );
  AOI221_X1 U7991 ( .B1(net227353), .B2(n17723), .C1(\registers[54][25] ), 
        .C2(n17720), .A(n5020), .ZN(n5017) );
  AOI221_X1 U7992 ( .B1(\registers[42][25] ), .B2(n17687), .C1(
        \registers[43][25] ), .C2(n17684), .A(n5023), .ZN(n5014) );
  NAND4_X1 U7993 ( .A1(n4892), .A2(n4895), .A3(n4898), .A4(n4899), .ZN(n4873)
         );
  AOI221_X1 U7994 ( .B1(net227370), .B2(n17711), .C1(net227369), .C2(n17708), 
        .A(n4901), .ZN(n4898) );
  AOI221_X1 U7995 ( .B1(net227371), .B2(n17723), .C1(\registers[54][26] ), 
        .C2(n17720), .A(n4900), .ZN(n4899) );
  AOI221_X1 U7996 ( .B1(\registers[42][26] ), .B2(n17687), .C1(
        \registers[43][26] ), .C2(n17684), .A(n4903), .ZN(n4892) );
  NAND4_X1 U7997 ( .A1(n4767), .A2(n4768), .A3(n4769), .A4(n4770), .ZN(n4740)
         );
  AOI221_X1 U7998 ( .B1(net227388), .B2(n17711), .C1(net227387), .C2(n17708), 
        .A(n4772), .ZN(n4769) );
  AOI221_X1 U7999 ( .B1(net227389), .B2(n17723), .C1(\registers[54][27] ), 
        .C2(n17720), .A(n4771), .ZN(n4770) );
  AOI221_X1 U8000 ( .B1(\registers[42][27] ), .B2(n17687), .C1(
        \registers[43][27] ), .C2(n17684), .A(n4774), .ZN(n4767) );
  NAND4_X1 U8001 ( .A1(n4634), .A2(n4635), .A3(n4636), .A4(n4637), .ZN(n4613)
         );
  AOI221_X1 U8002 ( .B1(net227406), .B2(n17711), .C1(net227405), .C2(n17708), 
        .A(n4639), .ZN(n4636) );
  AOI221_X1 U8003 ( .B1(net227407), .B2(n17723), .C1(\registers[54][28] ), 
        .C2(n17720), .A(n4638), .ZN(n4637) );
  AOI221_X1 U8004 ( .B1(\registers[42][28] ), .B2(n17687), .C1(
        \registers[43][28] ), .C2(n17684), .A(n4641), .ZN(n4634) );
  NAND4_X1 U8005 ( .A1(n4507), .A2(n4508), .A3(n4509), .A4(n4510), .ZN(n4482)
         );
  AOI221_X1 U8006 ( .B1(net227424), .B2(n17711), .C1(net227423), .C2(n17708), 
        .A(n4512), .ZN(n4509) );
  AOI221_X1 U8007 ( .B1(net227425), .B2(n17723), .C1(\registers[54][29] ), 
        .C2(n17720), .A(n4511), .ZN(n4510) );
  AOI221_X1 U8008 ( .B1(\registers[42][29] ), .B2(n17687), .C1(
        \registers[43][29] ), .C2(n17684), .A(n4514), .ZN(n4507) );
  NAND4_X1 U8009 ( .A1(n4177), .A2(n4178), .A3(n4179), .A4(n4180), .ZN(n4098)
         );
  AOI221_X1 U8010 ( .B1(net227442), .B2(n17711), .C1(net227441), .C2(n17708), 
        .A(n4190), .ZN(n4179) );
  AOI221_X1 U8011 ( .B1(net227443), .B2(n17723), .C1(\registers[54][30] ), 
        .C2(n17720), .A(n4183), .ZN(n4180) );
  AOI221_X1 U8012 ( .B1(\registers[42][30] ), .B2(n17687), .C1(
        \registers[43][30] ), .C2(n17684), .A(n4208), .ZN(n4177) );
  NAND4_X1 U8013 ( .A1(n12391), .A2(n12392), .A3(n12393), .A4(n12394), .ZN(
        n12372) );
  AOI221_X1 U8014 ( .B1(net226845), .B2(n17709), .C1(net226836), .C2(n17706), 
        .A(n12396), .ZN(n12393) );
  AOI221_X1 U8015 ( .B1(net226846), .B2(n17721), .C1(\registers[54][0] ), .C2(
        n17718), .A(n12395), .ZN(n12394) );
  AOI221_X1 U8016 ( .B1(\registers[42][0] ), .B2(n17685), .C1(
        \registers[43][0] ), .C2(n17682), .A(n12398), .ZN(n12391) );
  NAND4_X1 U8017 ( .A1(n12237), .A2(n12238), .A3(n12239), .A4(n12240), .ZN(
        n12218) );
  AOI221_X1 U8018 ( .B1(net226858), .B2(n17709), .C1(net226866), .C2(n17706), 
        .A(n12242), .ZN(n12239) );
  AOI221_X1 U8019 ( .B1(net226859), .B2(n17721), .C1(\registers[54][1] ), .C2(
        n17718), .A(n12241), .ZN(n12240) );
  AOI221_X1 U8020 ( .B1(\registers[42][1] ), .B2(n17685), .C1(
        \registers[43][1] ), .C2(n17682), .A(n12244), .ZN(n12237) );
  NAND4_X1 U8021 ( .A1(n12082), .A2(n12083), .A3(n12084), .A4(n12085), .ZN(
        n12063) );
  AOI221_X1 U8022 ( .B1(net226879), .B2(n17709), .C1(net226878), .C2(n17706), 
        .A(n12087), .ZN(n12084) );
  AOI221_X1 U8023 ( .B1(net226885), .B2(n17721), .C1(\registers[54][2] ), .C2(
        n17718), .A(n12086), .ZN(n12085) );
  AOI221_X1 U8024 ( .B1(\registers[42][2] ), .B2(n17685), .C1(
        \registers[43][2] ), .C2(n17682), .A(n12089), .ZN(n12082) );
  NAND4_X1 U8025 ( .A1(n11929), .A2(n11930), .A3(n11931), .A4(n11932), .ZN(
        n11910) );
  AOI221_X1 U8026 ( .B1(net226906), .B2(n17709), .C1(net226905), .C2(n17706), 
        .A(n11934), .ZN(n11931) );
  AOI221_X1 U8027 ( .B1(net226898), .B2(n17721), .C1(\registers[54][3] ), .C2(
        n17718), .A(n11933), .ZN(n11932) );
  AOI221_X1 U8028 ( .B1(\registers[42][3] ), .B2(n17685), .C1(
        \registers[43][3] ), .C2(n17682), .A(n11936), .ZN(n11929) );
  NAND4_X1 U8029 ( .A1(n10486), .A2(n10487), .A3(n10488), .A4(n10489), .ZN(
        n10467) );
  AOI221_X1 U8030 ( .B1(net226979), .B2(n17709), .C1(net226978), .C2(n17706), 
        .A(n10491), .ZN(n10488) );
  AOI221_X1 U8031 ( .B1(net226980), .B2(n17721), .C1(\registers[54][4] ), .C2(
        n17718), .A(n10490), .ZN(n10489) );
  AOI221_X1 U8032 ( .B1(\registers[42][4] ), .B2(n17685), .C1(
        \registers[43][4] ), .C2(n17682), .A(n10493), .ZN(n10486) );
  NAND4_X1 U8033 ( .A1(n10376), .A2(n10377), .A3(n10378), .A4(n10379), .ZN(
        n10357) );
  AOI221_X1 U8034 ( .B1(net226999), .B2(n17709), .C1(net226998), .C2(n17706), 
        .A(n10381), .ZN(n10378) );
  AOI221_X1 U8035 ( .B1(net227000), .B2(n17721), .C1(\registers[54][5] ), .C2(
        n17718), .A(n10380), .ZN(n10379) );
  AOI221_X1 U8036 ( .B1(\registers[42][5] ), .B2(n17685), .C1(
        \registers[43][5] ), .C2(n17682), .A(n10383), .ZN(n10376) );
  NAND4_X1 U8037 ( .A1(n10264), .A2(n10265), .A3(n10266), .A4(n10267), .ZN(
        n10245) );
  AOI221_X1 U8038 ( .B1(net227010), .B2(n17709), .C1(net227009), .C2(n17706), 
        .A(n10269), .ZN(n10266) );
  AOI221_X1 U8039 ( .B1(net227011), .B2(n17721), .C1(\registers[54][6] ), .C2(
        n17718), .A(n10268), .ZN(n10267) );
  AOI221_X1 U8040 ( .B1(\registers[42][6] ), .B2(n17685), .C1(
        \registers[43][6] ), .C2(n17682), .A(n10271), .ZN(n10264) );
  NAND4_X1 U8041 ( .A1(n7628), .A2(n7629), .A3(n7630), .A4(n7631), .ZN(n7609)
         );
  AOI221_X1 U8042 ( .B1(net227028), .B2(n17709), .C1(net227027), .C2(n17706), 
        .A(n7633), .ZN(n7630) );
  AOI221_X1 U8043 ( .B1(net227029), .B2(n17721), .C1(\registers[54][7] ), .C2(
        n17718), .A(n7632), .ZN(n7631) );
  AOI221_X1 U8044 ( .B1(\registers[42][7] ), .B2(n17685), .C1(
        \registers[43][7] ), .C2(n17682), .A(n7635), .ZN(n7628) );
  NAND4_X1 U8045 ( .A1(n7513), .A2(n7514), .A3(n7515), .A4(n7516), .ZN(n7494)
         );
  AOI221_X1 U8046 ( .B1(net227046), .B2(n17709), .C1(net227045), .C2(n17706), 
        .A(n7518), .ZN(n7515) );
  AOI221_X1 U8047 ( .B1(net227047), .B2(n17721), .C1(\registers[54][8] ), .C2(
        n17718), .A(n7517), .ZN(n7516) );
  AOI221_X1 U8048 ( .B1(\registers[42][8] ), .B2(n17685), .C1(
        \registers[43][8] ), .C2(n17682), .A(n7520), .ZN(n7513) );
  NAND4_X1 U8049 ( .A1(n7404), .A2(n7405), .A3(n7406), .A4(n7407), .ZN(n7385)
         );
  AOI221_X1 U8050 ( .B1(net227064), .B2(n17709), .C1(net227063), .C2(n17706), 
        .A(n7409), .ZN(n7406) );
  AOI221_X1 U8051 ( .B1(net227065), .B2(n17721), .C1(\registers[54][9] ), .C2(
        n17718), .A(n7408), .ZN(n7407) );
  AOI221_X1 U8052 ( .B1(\registers[42][9] ), .B2(n17685), .C1(
        \registers[43][9] ), .C2(n17682), .A(n7411), .ZN(n7404) );
  NAND4_X1 U8053 ( .A1(n7295), .A2(n7296), .A3(n7297), .A4(n7298), .ZN(n7276)
         );
  AOI221_X1 U8054 ( .B1(net227082), .B2(n17709), .C1(net227081), .C2(n17706), 
        .A(n7300), .ZN(n7297) );
  AOI221_X1 U8055 ( .B1(net227083), .B2(n17721), .C1(\registers[54][10] ), 
        .C2(n17718), .A(n7299), .ZN(n7298) );
  AOI221_X1 U8056 ( .B1(\registers[42][10] ), .B2(n17685), .C1(
        \registers[43][10] ), .C2(n17682), .A(n7302), .ZN(n7295) );
  NAND4_X1 U8057 ( .A1(n7181), .A2(n7182), .A3(n7183), .A4(n7184), .ZN(n7162)
         );
  AOI221_X1 U8058 ( .B1(net227100), .B2(n17710), .C1(net227099), .C2(n17707), 
        .A(n7186), .ZN(n7183) );
  AOI221_X1 U8059 ( .B1(net227101), .B2(n17722), .C1(\registers[54][11] ), 
        .C2(n17719), .A(n7185), .ZN(n7184) );
  AOI221_X1 U8060 ( .B1(\registers[42][11] ), .B2(n17686), .C1(
        \registers[43][11] ), .C2(n17683), .A(n7188), .ZN(n7181) );
  NAND4_X1 U8061 ( .A1(n7072), .A2(n7073), .A3(n7074), .A4(n7075), .ZN(n7053)
         );
  AOI221_X1 U8062 ( .B1(net227118), .B2(n17710), .C1(net227117), .C2(n17707), 
        .A(n7077), .ZN(n7074) );
  AOI221_X1 U8063 ( .B1(net227119), .B2(n17722), .C1(\registers[54][12] ), 
        .C2(n17719), .A(n7076), .ZN(n7075) );
  AOI221_X1 U8064 ( .B1(\registers[42][12] ), .B2(n17686), .C1(
        \registers[43][12] ), .C2(n17683), .A(n7079), .ZN(n7072) );
  NAND4_X1 U8065 ( .A1(n6963), .A2(n6964), .A3(n6965), .A4(n6966), .ZN(n6944)
         );
  AOI221_X1 U8066 ( .B1(net227136), .B2(n17710), .C1(net227135), .C2(n17707), 
        .A(n6968), .ZN(n6965) );
  AOI221_X1 U8067 ( .B1(net227137), .B2(n17722), .C1(\registers[54][13] ), 
        .C2(n17719), .A(n6967), .ZN(n6966) );
  AOI221_X1 U8068 ( .B1(\registers[42][13] ), .B2(n17686), .C1(
        \registers[43][13] ), .C2(n17683), .A(n6970), .ZN(n6963) );
  NAND4_X1 U8069 ( .A1(n6854), .A2(n6855), .A3(n6856), .A4(n6857), .ZN(n6835)
         );
  AOI221_X1 U8070 ( .B1(net227154), .B2(n17710), .C1(net227153), .C2(n17707), 
        .A(n6859), .ZN(n6856) );
  AOI221_X1 U8071 ( .B1(net227155), .B2(n17722), .C1(\registers[54][14] ), 
        .C2(n17719), .A(n6858), .ZN(n6857) );
  AOI221_X1 U8072 ( .B1(\registers[42][14] ), .B2(n17686), .C1(
        \registers[43][14] ), .C2(n17683), .A(n6861), .ZN(n6854) );
  NAND4_X1 U8073 ( .A1(n6745), .A2(n6746), .A3(n6747), .A4(n6748), .ZN(n6726)
         );
  AOI221_X1 U8074 ( .B1(net227172), .B2(n17710), .C1(net227171), .C2(n17707), 
        .A(n6750), .ZN(n6747) );
  AOI221_X1 U8075 ( .B1(net227173), .B2(n17722), .C1(\registers[54][15] ), 
        .C2(n17719), .A(n6749), .ZN(n6748) );
  AOI221_X1 U8076 ( .B1(\registers[42][15] ), .B2(n17686), .C1(
        \registers[43][15] ), .C2(n17683), .A(n6752), .ZN(n6745) );
  NAND4_X1 U8077 ( .A1(n6602), .A2(n6603), .A3(n6604), .A4(n6605), .ZN(n6563)
         );
  AOI221_X1 U8078 ( .B1(net227190), .B2(n17710), .C1(net227189), .C2(n17707), 
        .A(n6607), .ZN(n6604) );
  AOI221_X1 U8079 ( .B1(net227191), .B2(n17722), .C1(\registers[54][16] ), 
        .C2(n17719), .A(n6606), .ZN(n6605) );
  AOI221_X1 U8080 ( .B1(\registers[42][16] ), .B2(n17686), .C1(
        \registers[43][16] ), .C2(n17683), .A(n6610), .ZN(n6602) );
  NAND4_X1 U8081 ( .A1(n6415), .A2(n6416), .A3(n6417), .A4(n6418), .ZN(n6376)
         );
  AOI221_X1 U8082 ( .B1(net227208), .B2(n17710), .C1(net227207), .C2(n17707), 
        .A(n6421), .ZN(n6417) );
  AOI221_X1 U8083 ( .B1(net227209), .B2(n17722), .C1(\registers[54][17] ), 
        .C2(n17719), .A(n6420), .ZN(n6418) );
  AOI221_X1 U8084 ( .B1(\registers[42][17] ), .B2(n17686), .C1(
        \registers[43][17] ), .C2(n17683), .A(n6425), .ZN(n6415) );
  NAND4_X1 U8085 ( .A1(n6228), .A2(n6229), .A3(n6231), .A4(n6232), .ZN(n6190)
         );
  AOI221_X1 U8086 ( .B1(net227226), .B2(n17710), .C1(net227225), .C2(n17707), 
        .A(n6236), .ZN(n6231) );
  AOI221_X1 U8087 ( .B1(net227227), .B2(n17722), .C1(\registers[54][18] ), 
        .C2(n17719), .A(n6234), .ZN(n6232) );
  AOI221_X1 U8088 ( .B1(\registers[42][18] ), .B2(n17686), .C1(
        \registers[43][18] ), .C2(n17683), .A(n6238), .ZN(n6228) );
  NAND4_X1 U8089 ( .A1(n6042), .A2(n6043), .A3(n6045), .A4(n6047), .ZN(n6005)
         );
  AOI221_X1 U8090 ( .B1(net227244), .B2(n17710), .C1(net227243), .C2(n17707), 
        .A(n6049), .ZN(n6045) );
  AOI221_X1 U8091 ( .B1(net227245), .B2(n17722), .C1(\registers[54][19] ), 
        .C2(n17719), .A(n6048), .ZN(n6047) );
  AOI221_X1 U8092 ( .B1(\registers[42][19] ), .B2(n17686), .C1(
        \registers[43][19] ), .C2(n17683), .A(n6051), .ZN(n6042) );
  NAND4_X1 U8093 ( .A1(n5856), .A2(n5858), .A3(n5859), .A4(n5860), .ZN(n5818)
         );
  AOI221_X1 U8094 ( .B1(net227262), .B2(n17710), .C1(net227261), .C2(n17707), 
        .A(n5862), .ZN(n5859) );
  AOI221_X1 U8095 ( .B1(net227263), .B2(n17722), .C1(\registers[54][20] ), 
        .C2(n17719), .A(n5861), .ZN(n5860) );
  AOI221_X1 U8096 ( .B1(\registers[42][20] ), .B2(n17686), .C1(
        \registers[43][20] ), .C2(n17683), .A(n5866), .ZN(n5856) );
  NAND4_X1 U8097 ( .A1(n5670), .A2(n5671), .A3(n5672), .A4(n5673), .ZN(n5631)
         );
  AOI221_X1 U8098 ( .B1(net227280), .B2(n17710), .C1(net227279), .C2(n17707), 
        .A(n5677), .ZN(n5672) );
  AOI221_X1 U8099 ( .B1(net227281), .B2(n17722), .C1(\registers[54][21] ), 
        .C2(n17719), .A(n5674), .ZN(n5673) );
  AOI221_X1 U8100 ( .B1(\registers[42][21] ), .B2(n17686), .C1(
        \registers[43][21] ), .C2(n17683), .A(n5680), .ZN(n5670) );
  NAND4_X1 U8101 ( .A1(n5483), .A2(n5484), .A3(n5485), .A4(n5488), .ZN(n5446)
         );
  AOI221_X1 U8102 ( .B1(net227298), .B2(n17710), .C1(net227297), .C2(n17707), 
        .A(n5491), .ZN(n5485) );
  AOI221_X1 U8103 ( .B1(net227299), .B2(n17722), .C1(\registers[54][22] ), 
        .C2(n17719), .A(n5489), .ZN(n5488) );
  AOI221_X1 U8104 ( .B1(\registers[42][22] ), .B2(n17686), .C1(
        \registers[43][22] ), .C2(n17683), .A(n5493), .ZN(n5483) );
  NAND4_X1 U8105 ( .A1(n14153), .A2(n14154), .A3(n14155), .A4(n14156), .ZN(
        n14077) );
  AOI221_X1 U8106 ( .B1(net227460), .B2(n17709), .C1(net227459), .C2(n17706), 
        .A(n14161), .ZN(n14155) );
  AOI221_X1 U8107 ( .B1(net227461), .B2(n17721), .C1(\registers[54][31] ), 
        .C2(n17718), .A(n14157), .ZN(n14156) );
  AOI221_X1 U8108 ( .B1(\registers[42][31] ), .B2(n17685), .C1(
        \registers[43][31] ), .C2(n17682), .A(n14175), .ZN(n14153) );
  NAND4_X1 U8109 ( .A1(n13912), .A2(n13913), .A3(n13914), .A4(n13915), .ZN(
        n13911) );
  AOI211_X1 U8110 ( .C1(\registers[23][0] ), .C2(n16373), .A(n13934), .B(
        n16412), .ZN(n13912) );
  AOI221_X1 U8111 ( .B1(\registers[1][0] ), .B2(n16385), .C1(
        \registers[19][0] ), .C2(n16382), .A(n13930), .ZN(n13913) );
  AOI221_X1 U8112 ( .B1(\registers[16][0] ), .B2(n16397), .C1(
        \registers[15][0] ), .C2(n16394), .A(n13924), .ZN(n13914) );
  NAND4_X1 U8113 ( .A1(n13865), .A2(n13866), .A3(n13867), .A4(n13868), .ZN(
        n13864) );
  AOI211_X1 U8114 ( .C1(\registers[23][1] ), .C2(n16373), .A(n13872), .B(
        n16412), .ZN(n13865) );
  AOI221_X1 U8115 ( .B1(\registers[1][1] ), .B2(n16385), .C1(
        \registers[19][1] ), .C2(n16382), .A(n13871), .ZN(n13866) );
  AOI221_X1 U8116 ( .B1(\registers[16][1] ), .B2(n16397), .C1(
        \registers[15][1] ), .C2(n16394), .A(n13870), .ZN(n13867) );
  NAND4_X1 U8117 ( .A1(n13823), .A2(n13824), .A3(n13825), .A4(n13826), .ZN(
        n13822) );
  AOI211_X1 U8118 ( .C1(\registers[23][2] ), .C2(n16373), .A(n13830), .B(
        n16412), .ZN(n13823) );
  AOI221_X1 U8119 ( .B1(\registers[1][2] ), .B2(n16385), .C1(
        \registers[19][2] ), .C2(n16382), .A(n13829), .ZN(n13824) );
  AOI221_X1 U8120 ( .B1(\registers[16][2] ), .B2(n16397), .C1(
        \registers[15][2] ), .C2(n16394), .A(n13828), .ZN(n13825) );
  NAND4_X1 U8121 ( .A1(n13781), .A2(n13782), .A3(n13783), .A4(n13784), .ZN(
        n13780) );
  AOI211_X1 U8122 ( .C1(\registers[23][3] ), .C2(n16373), .A(n13788), .B(
        n16412), .ZN(n13781) );
  AOI221_X1 U8123 ( .B1(\registers[1][3] ), .B2(n16385), .C1(
        \registers[19][3] ), .C2(n16382), .A(n13787), .ZN(n13782) );
  AOI221_X1 U8124 ( .B1(\registers[16][3] ), .B2(n16397), .C1(
        \registers[15][3] ), .C2(n16394), .A(n13786), .ZN(n13783) );
  NAND4_X1 U8125 ( .A1(n13739), .A2(n13740), .A3(n13741), .A4(n13742), .ZN(
        n13738) );
  AOI211_X1 U8126 ( .C1(\registers[23][4] ), .C2(n16373), .A(n13746), .B(
        n16412), .ZN(n13739) );
  AOI221_X1 U8127 ( .B1(\registers[1][4] ), .B2(n16385), .C1(
        \registers[19][4] ), .C2(n16382), .A(n13745), .ZN(n13740) );
  AOI221_X1 U8128 ( .B1(\registers[16][4] ), .B2(n16397), .C1(
        \registers[15][4] ), .C2(n16394), .A(n13744), .ZN(n13741) );
  NAND4_X1 U8129 ( .A1(n13697), .A2(n13698), .A3(n13699), .A4(n13700), .ZN(
        n13696) );
  AOI211_X1 U8130 ( .C1(\registers[23][5] ), .C2(n16373), .A(n13704), .B(
        n16412), .ZN(n13697) );
  AOI221_X1 U8131 ( .B1(\registers[1][5] ), .B2(n16385), .C1(
        \registers[19][5] ), .C2(n16382), .A(n13703), .ZN(n13698) );
  AOI221_X1 U8132 ( .B1(\registers[16][5] ), .B2(n16397), .C1(
        \registers[15][5] ), .C2(n16394), .A(n13702), .ZN(n13699) );
  NAND4_X1 U8133 ( .A1(n13655), .A2(n13656), .A3(n13657), .A4(n13658), .ZN(
        n13654) );
  AOI211_X1 U8134 ( .C1(\registers[23][6] ), .C2(n16373), .A(n13662), .B(
        n16412), .ZN(n13655) );
  AOI221_X1 U8135 ( .B1(\registers[1][6] ), .B2(n16385), .C1(
        \registers[19][6] ), .C2(n16382), .A(n13661), .ZN(n13656) );
  AOI221_X1 U8136 ( .B1(\registers[16][6] ), .B2(n16397), .C1(
        \registers[15][6] ), .C2(n16394), .A(n13660), .ZN(n13657) );
  NAND4_X1 U8137 ( .A1(n13613), .A2(n13614), .A3(n13615), .A4(n13616), .ZN(
        n13612) );
  AOI211_X1 U8138 ( .C1(\registers[23][7] ), .C2(n16373), .A(n13620), .B(
        n16412), .ZN(n13613) );
  AOI221_X1 U8139 ( .B1(\registers[1][7] ), .B2(n16385), .C1(
        \registers[19][7] ), .C2(n16382), .A(n13619), .ZN(n13614) );
  AOI221_X1 U8140 ( .B1(\registers[16][7] ), .B2(n16397), .C1(
        \registers[15][7] ), .C2(n16394), .A(n13618), .ZN(n13615) );
  NAND4_X1 U8141 ( .A1(n13571), .A2(n13572), .A3(n13573), .A4(n13574), .ZN(
        n13570) );
  AOI211_X1 U8142 ( .C1(\registers[23][8] ), .C2(n16373), .A(n13578), .B(
        n16413), .ZN(n13571) );
  AOI221_X1 U8143 ( .B1(\registers[1][8] ), .B2(n16385), .C1(
        \registers[19][8] ), .C2(n16382), .A(n13577), .ZN(n13572) );
  AOI221_X1 U8144 ( .B1(\registers[16][8] ), .B2(n16397), .C1(
        \registers[15][8] ), .C2(n16394), .A(n13576), .ZN(n13573) );
  NAND4_X1 U8145 ( .A1(n13529), .A2(n13530), .A3(n13531), .A4(n13532), .ZN(
        n13528) );
  AOI211_X1 U8146 ( .C1(\registers[23][9] ), .C2(n16373), .A(n13536), .B(
        n16413), .ZN(n13529) );
  AOI221_X1 U8147 ( .B1(\registers[1][9] ), .B2(n16385), .C1(
        \registers[19][9] ), .C2(n16382), .A(n13535), .ZN(n13530) );
  AOI221_X1 U8148 ( .B1(\registers[16][9] ), .B2(n16397), .C1(
        \registers[15][9] ), .C2(n16394), .A(n13534), .ZN(n13531) );
  NAND4_X1 U8149 ( .A1(n13487), .A2(n13488), .A3(n13489), .A4(n13490), .ZN(
        n13486) );
  AOI211_X1 U8150 ( .C1(\registers[23][10] ), .C2(n16373), .A(n13494), .B(
        n16413), .ZN(n13487) );
  AOI221_X1 U8151 ( .B1(\registers[1][10] ), .B2(n16385), .C1(
        \registers[19][10] ), .C2(n16382), .A(n13493), .ZN(n13488) );
  AOI221_X1 U8152 ( .B1(\registers[16][10] ), .B2(n16397), .C1(
        \registers[15][10] ), .C2(n16394), .A(n13492), .ZN(n13489) );
  NAND4_X1 U8153 ( .A1(n13445), .A2(n13446), .A3(n13447), .A4(n13448), .ZN(
        n13444) );
  AOI211_X1 U8154 ( .C1(\registers[23][11] ), .C2(n16373), .A(n13452), .B(
        n16413), .ZN(n13445) );
  AOI221_X1 U8155 ( .B1(\registers[1][11] ), .B2(n16385), .C1(
        \registers[19][11] ), .C2(n16382), .A(n13451), .ZN(n13446) );
  AOI221_X1 U8156 ( .B1(\registers[16][11] ), .B2(n16397), .C1(
        \registers[15][11] ), .C2(n16394), .A(n13450), .ZN(n13447) );
  NAND4_X1 U8157 ( .A1(n13403), .A2(n13404), .A3(n13405), .A4(n13406), .ZN(
        n13402) );
  AOI211_X1 U8158 ( .C1(\registers[23][12] ), .C2(n16374), .A(n13410), .B(
        n16413), .ZN(n13403) );
  AOI221_X1 U8159 ( .B1(\registers[1][12] ), .B2(n16386), .C1(
        \registers[19][12] ), .C2(n16383), .A(n13409), .ZN(n13404) );
  AOI221_X1 U8160 ( .B1(\registers[16][12] ), .B2(n16398), .C1(
        \registers[15][12] ), .C2(n16395), .A(n13408), .ZN(n13405) );
  NAND4_X1 U8161 ( .A1(n13361), .A2(n13362), .A3(n13363), .A4(n13364), .ZN(
        n13360) );
  AOI211_X1 U8162 ( .C1(\registers[23][13] ), .C2(n16374), .A(n13368), .B(
        n16413), .ZN(n13361) );
  AOI221_X1 U8163 ( .B1(\registers[1][13] ), .B2(n16386), .C1(
        \registers[19][13] ), .C2(n16383), .A(n13367), .ZN(n13362) );
  AOI221_X1 U8164 ( .B1(\registers[16][13] ), .B2(n16398), .C1(
        \registers[15][13] ), .C2(n16395), .A(n13366), .ZN(n13363) );
  NAND4_X1 U8165 ( .A1(n13319), .A2(n13320), .A3(n13321), .A4(n13322), .ZN(
        n13318) );
  AOI211_X1 U8166 ( .C1(\registers[23][14] ), .C2(n16374), .A(n13326), .B(
        n16413), .ZN(n13319) );
  AOI221_X1 U8167 ( .B1(\registers[1][14] ), .B2(n16386), .C1(
        \registers[19][14] ), .C2(n16383), .A(n13325), .ZN(n13320) );
  AOI221_X1 U8168 ( .B1(\registers[16][14] ), .B2(n16398), .C1(
        \registers[15][14] ), .C2(n16395), .A(n13324), .ZN(n13321) );
  NAND4_X1 U8169 ( .A1(n13277), .A2(n13278), .A3(n13279), .A4(n13280), .ZN(
        n13276) );
  AOI211_X1 U8170 ( .C1(\registers[23][15] ), .C2(n16374), .A(n13284), .B(
        n16413), .ZN(n13277) );
  AOI221_X1 U8171 ( .B1(\registers[1][15] ), .B2(n16386), .C1(
        \registers[19][15] ), .C2(n16383), .A(n13283), .ZN(n13278) );
  AOI221_X1 U8172 ( .B1(\registers[16][15] ), .B2(n16398), .C1(
        \registers[15][15] ), .C2(n16395), .A(n13282), .ZN(n13279) );
  NAND4_X1 U8173 ( .A1(n13151), .A2(n13152), .A3(n13153), .A4(n13154), .ZN(
        n13150) );
  AOI211_X1 U8174 ( .C1(\registers[23][18] ), .C2(n16374), .A(n13158), .B(
        n16413), .ZN(n13151) );
  AOI221_X1 U8175 ( .B1(\registers[1][18] ), .B2(n16386), .C1(
        \registers[19][18] ), .C2(n16383), .A(n13157), .ZN(n13152) );
  AOI221_X1 U8176 ( .B1(\registers[16][18] ), .B2(n16398), .C1(
        \registers[15][18] ), .C2(n16395), .A(n13156), .ZN(n13153) );
  NAND4_X1 U8177 ( .A1(n12857), .A2(n12858), .A3(n12859), .A4(n12860), .ZN(
        n12856) );
  AOI211_X1 U8178 ( .C1(\registers[23][25] ), .C2(n16375), .A(n12864), .B(
        n16413), .ZN(n12857) );
  AOI221_X1 U8179 ( .B1(\registers[1][25] ), .B2(n16387), .C1(
        \registers[19][25] ), .C2(n16384), .A(n12863), .ZN(n12858) );
  AOI221_X1 U8180 ( .B1(\registers[16][25] ), .B2(n16399), .C1(
        \registers[15][25] ), .C2(n16396), .A(n12862), .ZN(n12859) );
  NAND4_X1 U8181 ( .A1(n12815), .A2(n12816), .A3(n12817), .A4(n12818), .ZN(
        n12814) );
  AOI211_X1 U8182 ( .C1(\registers[23][26] ), .C2(n16375), .A(n12822), .B(
        n16413), .ZN(n12815) );
  AOI221_X1 U8183 ( .B1(\registers[1][26] ), .B2(n16387), .C1(
        \registers[19][26] ), .C2(n16384), .A(n12821), .ZN(n12816) );
  AOI221_X1 U8184 ( .B1(\registers[16][26] ), .B2(n16399), .C1(
        \registers[15][26] ), .C2(n16396), .A(n12820), .ZN(n12817) );
  NAND4_X1 U8185 ( .A1(n12773), .A2(n12774), .A3(n12775), .A4(n12776), .ZN(
        n12772) );
  AOI211_X1 U8186 ( .C1(\registers[23][27] ), .C2(n16375), .A(n12780), .B(
        n16413), .ZN(n12773) );
  AOI221_X1 U8187 ( .B1(\registers[1][27] ), .B2(n16387), .C1(
        \registers[19][27] ), .C2(n16384), .A(n12779), .ZN(n12774) );
  AOI221_X1 U8188 ( .B1(\registers[16][27] ), .B2(n16399), .C1(
        \registers[15][27] ), .C2(n16396), .A(n12778), .ZN(n12775) );
  NAND4_X1 U8189 ( .A1(n12731), .A2(n12732), .A3(n12733), .A4(n12734), .ZN(
        n12730) );
  AOI211_X1 U8190 ( .C1(\registers[23][28] ), .C2(n16375), .A(n12738), .B(
        n16412), .ZN(n12731) );
  AOI221_X1 U8191 ( .B1(\registers[1][28] ), .B2(n16387), .C1(
        \registers[19][28] ), .C2(n16384), .A(n12737), .ZN(n12732) );
  AOI221_X1 U8192 ( .B1(\registers[16][28] ), .B2(n16399), .C1(
        \registers[15][28] ), .C2(n16396), .A(n12736), .ZN(n12733) );
  NAND4_X1 U8193 ( .A1(n12689), .A2(n12690), .A3(n12691), .A4(n12692), .ZN(
        n12688) );
  AOI211_X1 U8194 ( .C1(\registers[23][29] ), .C2(n16375), .A(n12696), .B(
        n16412), .ZN(n12689) );
  AOI221_X1 U8195 ( .B1(\registers[1][29] ), .B2(n16387), .C1(
        \registers[19][29] ), .C2(n16384), .A(n12695), .ZN(n12690) );
  AOI221_X1 U8196 ( .B1(\registers[16][29] ), .B2(n16399), .C1(
        \registers[15][29] ), .C2(n16396), .A(n12694), .ZN(n12691) );
  NAND4_X1 U8197 ( .A1(n12645), .A2(n12646), .A3(n12647), .A4(n12648), .ZN(
        n12644) );
  AOI211_X1 U8198 ( .C1(\registers[23][30] ), .C2(n16375), .A(n12653), .B(
        n16412), .ZN(n12645) );
  AOI221_X1 U8199 ( .B1(\registers[1][30] ), .B2(n16387), .C1(
        \registers[19][30] ), .C2(n16384), .A(n12651), .ZN(n12646) );
  AOI221_X1 U8200 ( .B1(\registers[16][30] ), .B2(n16399), .C1(
        \registers[15][30] ), .C2(n16396), .A(n12650), .ZN(n12647) );
  NAND4_X1 U8201 ( .A1(n12533), .A2(n12534), .A3(n12535), .A4(n12536), .ZN(
        n12532) );
  AOI211_X1 U8202 ( .C1(\registers[23][31] ), .C2(n16375), .A(n12554), .B(
        n16412), .ZN(n12533) );
  AOI221_X1 U8203 ( .B1(\registers[1][31] ), .B2(n16387), .C1(
        \registers[19][31] ), .C2(n16384), .A(n12549), .ZN(n12534) );
  AOI221_X1 U8204 ( .B1(\registers[16][31] ), .B2(n16399), .C1(
        \registers[15][31] ), .C2(n16396), .A(n12544), .ZN(n12535) );
  NAND4_X1 U8205 ( .A1(n12431), .A2(n12432), .A3(n12433), .A4(n12434), .ZN(
        n12430) );
  AOI221_X1 U8206 ( .B1(\registers[16][0] ), .B2(n16649), .C1(
        \registers[19][0] ), .C2(n16646), .A(n12442), .ZN(n12433) );
  AOI211_X1 U8207 ( .C1(\registers[23][0] ), .C2(n16625), .A(n12453), .B(
        n16664), .ZN(n12431) );
  AOI221_X1 U8208 ( .B1(\registers[1][0] ), .B2(n16637), .C1(
        \registers[22][0] ), .C2(n16634), .A(n12448), .ZN(n12432) );
  NAND4_X1 U8209 ( .A1(n12269), .A2(n12270), .A3(n12271), .A4(n12272), .ZN(
        n12268) );
  AOI221_X1 U8210 ( .B1(\registers[16][1] ), .B2(n16649), .C1(
        \registers[19][1] ), .C2(n16646), .A(n12274), .ZN(n12271) );
  AOI211_X1 U8211 ( .C1(\registers[23][1] ), .C2(n16625), .A(n12276), .B(
        n16664), .ZN(n12269) );
  AOI221_X1 U8212 ( .B1(\registers[1][1] ), .B2(n16637), .C1(
        \registers[22][1] ), .C2(n16634), .A(n12275), .ZN(n12270) );
  NAND4_X1 U8213 ( .A1(n12116), .A2(n12117), .A3(n12118), .A4(n12119), .ZN(
        n12115) );
  AOI221_X1 U8214 ( .B1(\registers[16][2] ), .B2(n16649), .C1(
        \registers[19][2] ), .C2(n16646), .A(n12121), .ZN(n12118) );
  AOI211_X1 U8215 ( .C1(\registers[23][2] ), .C2(n16625), .A(n12123), .B(
        n16664), .ZN(n12116) );
  AOI221_X1 U8216 ( .B1(\registers[1][2] ), .B2(n16637), .C1(
        \registers[22][2] ), .C2(n16634), .A(n12122), .ZN(n12117) );
  NAND4_X1 U8217 ( .A1(n11963), .A2(n11964), .A3(n11965), .A4(n11966), .ZN(
        n11962) );
  AOI221_X1 U8218 ( .B1(\registers[16][3] ), .B2(n16649), .C1(
        \registers[19][3] ), .C2(n16646), .A(n11968), .ZN(n11965) );
  AOI211_X1 U8219 ( .C1(\registers[23][3] ), .C2(n16625), .A(n11970), .B(
        n16664), .ZN(n11963) );
  AOI221_X1 U8220 ( .B1(\registers[1][3] ), .B2(n16637), .C1(
        \registers[22][3] ), .C2(n16634), .A(n11969), .ZN(n11964) );
  NAND4_X1 U8221 ( .A1(n11810), .A2(n11811), .A3(n11812), .A4(n11813), .ZN(
        n11809) );
  AOI221_X1 U8222 ( .B1(\registers[16][4] ), .B2(n16649), .C1(
        \registers[19][4] ), .C2(n16646), .A(n11815), .ZN(n11812) );
  AOI211_X1 U8223 ( .C1(\registers[23][4] ), .C2(n16625), .A(n11817), .B(
        n16664), .ZN(n11810) );
  AOI221_X1 U8224 ( .B1(\registers[1][4] ), .B2(n16637), .C1(
        \registers[22][4] ), .C2(n16634), .A(n11816), .ZN(n11811) );
  NAND4_X1 U8225 ( .A1(n11767), .A2(n11768), .A3(n11769), .A4(n11770), .ZN(
        n11766) );
  AOI221_X1 U8226 ( .B1(\registers[16][5] ), .B2(n16649), .C1(
        \registers[19][5] ), .C2(n16646), .A(n11772), .ZN(n11769) );
  AOI211_X1 U8227 ( .C1(\registers[23][5] ), .C2(n16625), .A(n11774), .B(
        n16664), .ZN(n11767) );
  AOI221_X1 U8228 ( .B1(\registers[1][5] ), .B2(n16637), .C1(
        \registers[22][5] ), .C2(n16634), .A(n11773), .ZN(n11768) );
  NAND4_X1 U8229 ( .A1(n11724), .A2(n11725), .A3(n11726), .A4(n11727), .ZN(
        n11723) );
  AOI221_X1 U8230 ( .B1(\registers[16][6] ), .B2(n16649), .C1(
        \registers[19][6] ), .C2(n16646), .A(n11729), .ZN(n11726) );
  AOI211_X1 U8231 ( .C1(\registers[23][6] ), .C2(n16625), .A(n11731), .B(
        n16664), .ZN(n11724) );
  AOI221_X1 U8232 ( .B1(\registers[1][6] ), .B2(n16637), .C1(
        \registers[22][6] ), .C2(n16634), .A(n11730), .ZN(n11725) );
  NAND4_X1 U8233 ( .A1(n11681), .A2(n11682), .A3(n11683), .A4(n11684), .ZN(
        n11680) );
  AOI221_X1 U8234 ( .B1(\registers[16][7] ), .B2(n16649), .C1(
        \registers[19][7] ), .C2(n16646), .A(n11686), .ZN(n11683) );
  AOI211_X1 U8235 ( .C1(\registers[23][7] ), .C2(n16625), .A(n11688), .B(
        n16664), .ZN(n11681) );
  AOI221_X1 U8236 ( .B1(\registers[1][7] ), .B2(n16637), .C1(
        \registers[22][7] ), .C2(n16634), .A(n11687), .ZN(n11682) );
  NAND4_X1 U8237 ( .A1(n11638), .A2(n11639), .A3(n11640), .A4(n11641), .ZN(
        n11637) );
  AOI221_X1 U8238 ( .B1(\registers[16][8] ), .B2(n16649), .C1(
        \registers[19][8] ), .C2(n16646), .A(n11643), .ZN(n11640) );
  AOI211_X1 U8239 ( .C1(\registers[23][8] ), .C2(n16625), .A(n11645), .B(
        n16665), .ZN(n11638) );
  AOI221_X1 U8240 ( .B1(\registers[1][8] ), .B2(n16637), .C1(
        \registers[22][8] ), .C2(n16634), .A(n11644), .ZN(n11639) );
  NAND4_X1 U8241 ( .A1(n11595), .A2(n11596), .A3(n11597), .A4(n11598), .ZN(
        n11594) );
  AOI221_X1 U8242 ( .B1(\registers[16][9] ), .B2(n16649), .C1(
        \registers[19][9] ), .C2(n16646), .A(n11600), .ZN(n11597) );
  AOI211_X1 U8243 ( .C1(\registers[23][9] ), .C2(n16625), .A(n11602), .B(
        n16665), .ZN(n11595) );
  AOI221_X1 U8244 ( .B1(\registers[1][9] ), .B2(n16637), .C1(
        \registers[22][9] ), .C2(n16634), .A(n11601), .ZN(n11596) );
  NAND4_X1 U8245 ( .A1(n11552), .A2(n11553), .A3(n11554), .A4(n11555), .ZN(
        n11551) );
  AOI221_X1 U8246 ( .B1(\registers[16][10] ), .B2(n16649), .C1(
        \registers[19][10] ), .C2(n16646), .A(n11557), .ZN(n11554) );
  AOI211_X1 U8247 ( .C1(\registers[23][10] ), .C2(n16625), .A(n11559), .B(
        n16665), .ZN(n11552) );
  AOI221_X1 U8248 ( .B1(\registers[1][10] ), .B2(n16637), .C1(
        \registers[22][10] ), .C2(n16634), .A(n11558), .ZN(n11553) );
  NAND4_X1 U8249 ( .A1(n11509), .A2(n11510), .A3(n11511), .A4(n11512), .ZN(
        n11508) );
  AOI221_X1 U8250 ( .B1(\registers[16][11] ), .B2(n16649), .C1(
        \registers[19][11] ), .C2(n16646), .A(n11514), .ZN(n11511) );
  AOI211_X1 U8251 ( .C1(\registers[23][11] ), .C2(n16625), .A(n11516), .B(
        n16665), .ZN(n11509) );
  AOI221_X1 U8252 ( .B1(\registers[1][11] ), .B2(n16637), .C1(
        \registers[22][11] ), .C2(n16634), .A(n11515), .ZN(n11510) );
  NAND4_X1 U8253 ( .A1(n11466), .A2(n11467), .A3(n11468), .A4(n11469), .ZN(
        n11465) );
  AOI221_X1 U8254 ( .B1(\registers[16][12] ), .B2(n16650), .C1(
        \registers[19][12] ), .C2(n16647), .A(n11471), .ZN(n11468) );
  AOI211_X1 U8255 ( .C1(\registers[23][12] ), .C2(n16626), .A(n11473), .B(
        n16665), .ZN(n11466) );
  AOI221_X1 U8256 ( .B1(\registers[1][12] ), .B2(n16638), .C1(
        \registers[22][12] ), .C2(n16635), .A(n11472), .ZN(n11467) );
  NAND4_X1 U8257 ( .A1(n11422), .A2(n11423), .A3(n11424), .A4(n11425), .ZN(
        n11421) );
  AOI221_X1 U8258 ( .B1(\registers[16][13] ), .B2(n16650), .C1(
        \registers[19][13] ), .C2(n16647), .A(n11427), .ZN(n11424) );
  AOI211_X1 U8259 ( .C1(\registers[23][13] ), .C2(n16626), .A(n11429), .B(
        n16665), .ZN(n11422) );
  AOI221_X1 U8260 ( .B1(\registers[1][13] ), .B2(n16638), .C1(
        \registers[22][13] ), .C2(n16635), .A(n11428), .ZN(n11423) );
  NAND4_X1 U8261 ( .A1(n11379), .A2(n11380), .A3(n11381), .A4(n11382), .ZN(
        n11378) );
  AOI221_X1 U8262 ( .B1(\registers[16][14] ), .B2(n16650), .C1(
        \registers[19][14] ), .C2(n16647), .A(n11384), .ZN(n11381) );
  AOI211_X1 U8263 ( .C1(\registers[23][14] ), .C2(n16626), .A(n11386), .B(
        n16665), .ZN(n11379) );
  AOI221_X1 U8264 ( .B1(\registers[1][14] ), .B2(n16638), .C1(
        \registers[22][14] ), .C2(n16635), .A(n11385), .ZN(n11380) );
  NAND4_X1 U8265 ( .A1(n11336), .A2(n11337), .A3(n11338), .A4(n11339), .ZN(
        n11335) );
  AOI221_X1 U8266 ( .B1(\registers[16][15] ), .B2(n16650), .C1(
        \registers[19][15] ), .C2(n16647), .A(n11341), .ZN(n11338) );
  AOI211_X1 U8267 ( .C1(\registers[23][15] ), .C2(n16626), .A(n11343), .B(
        n16665), .ZN(n11336) );
  AOI221_X1 U8268 ( .B1(\registers[1][15] ), .B2(n16638), .C1(
        \registers[22][15] ), .C2(n16635), .A(n11342), .ZN(n11337) );
  NAND4_X1 U8269 ( .A1(n11207), .A2(n11208), .A3(n11209), .A4(n11210), .ZN(
        n11206) );
  AOI221_X1 U8270 ( .B1(\registers[16][18] ), .B2(n16650), .C1(
        \registers[19][18] ), .C2(n16647), .A(n11212), .ZN(n11209) );
  AOI211_X1 U8271 ( .C1(\registers[23][18] ), .C2(n16626), .A(n11214), .B(
        n16665), .ZN(n11207) );
  AOI221_X1 U8272 ( .B1(\registers[1][18] ), .B2(n16638), .C1(
        \registers[22][18] ), .C2(n16635), .A(n11213), .ZN(n11208) );
  NAND4_X1 U8273 ( .A1(n10906), .A2(n10907), .A3(n10908), .A4(n10909), .ZN(
        n10905) );
  AOI221_X1 U8274 ( .B1(\registers[16][25] ), .B2(n16651), .C1(
        \registers[19][25] ), .C2(n16648), .A(n10911), .ZN(n10908) );
  AOI211_X1 U8275 ( .C1(\registers[23][25] ), .C2(n16627), .A(n10913), .B(
        n16665), .ZN(n10906) );
  AOI221_X1 U8276 ( .B1(\registers[1][25] ), .B2(n16639), .C1(
        \registers[22][25] ), .C2(n16636), .A(n10912), .ZN(n10907) );
  NAND4_X1 U8277 ( .A1(n10863), .A2(n10864), .A3(n10865), .A4(n10866), .ZN(
        n10862) );
  AOI221_X1 U8278 ( .B1(\registers[16][26] ), .B2(n16651), .C1(
        \registers[19][26] ), .C2(n16648), .A(n10868), .ZN(n10865) );
  AOI211_X1 U8279 ( .C1(\registers[23][26] ), .C2(n16627), .A(n10870), .B(
        n16665), .ZN(n10863) );
  AOI221_X1 U8280 ( .B1(\registers[1][26] ), .B2(n16639), .C1(
        \registers[22][26] ), .C2(n16636), .A(n10869), .ZN(n10864) );
  NAND4_X1 U8281 ( .A1(n10820), .A2(n10821), .A3(n10822), .A4(n10823), .ZN(
        n10819) );
  AOI221_X1 U8282 ( .B1(\registers[16][27] ), .B2(n16651), .C1(
        \registers[19][27] ), .C2(n16648), .A(n10825), .ZN(n10822) );
  AOI211_X1 U8283 ( .C1(\registers[23][27] ), .C2(n16627), .A(n10827), .B(
        n16665), .ZN(n10820) );
  AOI221_X1 U8284 ( .B1(\registers[1][27] ), .B2(n16639), .C1(
        \registers[22][27] ), .C2(n16636), .A(n10826), .ZN(n10821) );
  NAND4_X1 U8285 ( .A1(n10777), .A2(n10778), .A3(n10779), .A4(n10780), .ZN(
        n10776) );
  AOI221_X1 U8286 ( .B1(\registers[16][28] ), .B2(n16651), .C1(
        \registers[19][28] ), .C2(n16648), .A(n10782), .ZN(n10779) );
  AOI211_X1 U8287 ( .C1(\registers[23][28] ), .C2(n16627), .A(n10784), .B(
        n16664), .ZN(n10777) );
  AOI221_X1 U8288 ( .B1(\registers[1][28] ), .B2(n16639), .C1(
        \registers[22][28] ), .C2(n16636), .A(n10783), .ZN(n10778) );
  NAND4_X1 U8289 ( .A1(n10734), .A2(n10735), .A3(n10736), .A4(n10737), .ZN(
        n10733) );
  AOI221_X1 U8290 ( .B1(\registers[16][29] ), .B2(n16651), .C1(
        \registers[19][29] ), .C2(n16648), .A(n10739), .ZN(n10736) );
  AOI211_X1 U8291 ( .C1(\registers[23][29] ), .C2(n16627), .A(n10741), .B(
        n16664), .ZN(n10734) );
  AOI221_X1 U8292 ( .B1(\registers[1][29] ), .B2(n16639), .C1(
        \registers[22][29] ), .C2(n16636), .A(n10740), .ZN(n10735) );
  NAND4_X1 U8293 ( .A1(n10675), .A2(n10676), .A3(n10677), .A4(n10678), .ZN(
        n10674) );
  AOI221_X1 U8294 ( .B1(\registers[16][30] ), .B2(n16651), .C1(
        \registers[19][30] ), .C2(n16648), .A(n10682), .ZN(n10677) );
  AOI211_X1 U8295 ( .C1(\registers[23][30] ), .C2(n16627), .A(n10685), .B(
        n16664), .ZN(n10675) );
  AOI221_X1 U8296 ( .B1(\registers[1][30] ), .B2(n16639), .C1(
        \registers[22][30] ), .C2(n16636), .A(n10683), .ZN(n10676) );
  NAND4_X1 U8297 ( .A1(n10531), .A2(n10532), .A3(n10533), .A4(n10534), .ZN(
        n10530) );
  AOI221_X1 U8298 ( .B1(\registers[16][31] ), .B2(n16651), .C1(
        \registers[19][31] ), .C2(n16648), .A(n10544), .ZN(n10533) );
  AOI211_X1 U8299 ( .C1(\registers[23][31] ), .C2(n16627), .A(n10557), .B(
        n16664), .ZN(n10531) );
  AOI221_X1 U8300 ( .B1(\registers[1][31] ), .B2(n16639), .C1(
        \registers[22][31] ), .C2(n16636), .A(n10551), .ZN(n10532) );
  NAND4_X1 U8301 ( .A1(n13235), .A2(n13236), .A3(n13237), .A4(n13238), .ZN(
        n13234) );
  AOI211_X1 U8302 ( .C1(\registers[23][16] ), .C2(n16374), .A(n13242), .B(
        n16414), .ZN(n13235) );
  AOI221_X1 U8303 ( .B1(\registers[1][16] ), .B2(n16386), .C1(
        \registers[19][16] ), .C2(n16383), .A(n13241), .ZN(n13236) );
  AOI221_X1 U8304 ( .B1(\registers[16][16] ), .B2(n16398), .C1(
        \registers[15][16] ), .C2(n16395), .A(n13240), .ZN(n13237) );
  NAND4_X1 U8305 ( .A1(n13193), .A2(n13194), .A3(n13195), .A4(n13196), .ZN(
        n13192) );
  AOI211_X1 U8306 ( .C1(\registers[23][17] ), .C2(n16374), .A(n13200), .B(
        n16414), .ZN(n13193) );
  AOI221_X1 U8307 ( .B1(\registers[1][17] ), .B2(n16386), .C1(
        \registers[19][17] ), .C2(n16383), .A(n13199), .ZN(n13194) );
  AOI221_X1 U8308 ( .B1(\registers[16][17] ), .B2(n16398), .C1(
        \registers[15][17] ), .C2(n16395), .A(n13198), .ZN(n13195) );
  NAND4_X1 U8309 ( .A1(n13109), .A2(n13110), .A3(n13111), .A4(n13112), .ZN(
        n13108) );
  AOI211_X1 U8310 ( .C1(\registers[23][19] ), .C2(n16374), .A(n13116), .B(
        n16414), .ZN(n13109) );
  AOI221_X1 U8311 ( .B1(\registers[1][19] ), .B2(n16386), .C1(
        \registers[19][19] ), .C2(n16383), .A(n13115), .ZN(n13110) );
  AOI221_X1 U8312 ( .B1(\registers[16][19] ), .B2(n16398), .C1(
        \registers[15][19] ), .C2(n16395), .A(n13114), .ZN(n13111) );
  NAND4_X1 U8313 ( .A1(n13067), .A2(n13068), .A3(n13069), .A4(n13070), .ZN(
        n13066) );
  AOI211_X1 U8314 ( .C1(\registers[23][20] ), .C2(n16374), .A(n13074), .B(
        n16414), .ZN(n13067) );
  AOI221_X1 U8315 ( .B1(\registers[1][20] ), .B2(n16386), .C1(
        \registers[19][20] ), .C2(n16383), .A(n13073), .ZN(n13068) );
  AOI221_X1 U8316 ( .B1(\registers[16][20] ), .B2(n16398), .C1(
        \registers[15][20] ), .C2(n16395), .A(n13072), .ZN(n13069) );
  NAND4_X1 U8317 ( .A1(n13025), .A2(n13026), .A3(n13027), .A4(n13028), .ZN(
        n13024) );
  AOI211_X1 U8318 ( .C1(\registers[23][21] ), .C2(n16374), .A(n13032), .B(
        n16414), .ZN(n13025) );
  AOI221_X1 U8319 ( .B1(\registers[1][21] ), .B2(n16386), .C1(
        \registers[19][21] ), .C2(n16383), .A(n13031), .ZN(n13026) );
  AOI221_X1 U8320 ( .B1(\registers[16][21] ), .B2(n16398), .C1(
        \registers[15][21] ), .C2(n16395), .A(n13030), .ZN(n13027) );
  NAND4_X1 U8321 ( .A1(n12983), .A2(n12984), .A3(n12985), .A4(n12986), .ZN(
        n12982) );
  AOI211_X1 U8322 ( .C1(\registers[23][22] ), .C2(n16374), .A(n12990), .B(
        n16414), .ZN(n12983) );
  AOI221_X1 U8323 ( .B1(\registers[1][22] ), .B2(n16386), .C1(
        \registers[19][22] ), .C2(n16383), .A(n12989), .ZN(n12984) );
  AOI221_X1 U8324 ( .B1(\registers[16][22] ), .B2(n16398), .C1(
        \registers[15][22] ), .C2(n16395), .A(n12988), .ZN(n12985) );
  NAND4_X1 U8325 ( .A1(n12941), .A2(n12942), .A3(n12943), .A4(n12944), .ZN(
        n12940) );
  AOI211_X1 U8326 ( .C1(\registers[23][23] ), .C2(n16374), .A(n12948), .B(
        n16414), .ZN(n12941) );
  AOI221_X1 U8327 ( .B1(\registers[1][23] ), .B2(n16386), .C1(
        \registers[19][23] ), .C2(n16383), .A(n12947), .ZN(n12942) );
  AOI221_X1 U8328 ( .B1(\registers[16][23] ), .B2(n16398), .C1(
        \registers[15][23] ), .C2(n16395), .A(n12946), .ZN(n12943) );
  NAND4_X1 U8329 ( .A1(n12899), .A2(n12900), .A3(n12901), .A4(n12902), .ZN(
        n12898) );
  AOI211_X1 U8330 ( .C1(\registers[23][24] ), .C2(n16375), .A(n12906), .B(
        n16414), .ZN(n12899) );
  AOI221_X1 U8331 ( .B1(\registers[1][24] ), .B2(n16387), .C1(
        \registers[19][24] ), .C2(n16384), .A(n12905), .ZN(n12900) );
  AOI221_X1 U8332 ( .B1(\registers[16][24] ), .B2(n16399), .C1(
        \registers[15][24] ), .C2(n16396), .A(n12904), .ZN(n12901) );
  NAND4_X1 U8333 ( .A1(n11293), .A2(n11294), .A3(n11295), .A4(n11296), .ZN(
        n11292) );
  AOI221_X1 U8334 ( .B1(\registers[16][16] ), .B2(n16650), .C1(
        \registers[19][16] ), .C2(n16647), .A(n11298), .ZN(n11295) );
  AOI211_X1 U8335 ( .C1(\registers[23][16] ), .C2(n16626), .A(n11300), .B(
        n16666), .ZN(n11293) );
  AOI221_X1 U8336 ( .B1(\registers[1][16] ), .B2(n16638), .C1(
        \registers[22][16] ), .C2(n16635), .A(n11299), .ZN(n11294) );
  NAND4_X1 U8337 ( .A1(n11250), .A2(n11251), .A3(n11252), .A4(n11253), .ZN(
        n11249) );
  AOI221_X1 U8338 ( .B1(\registers[16][17] ), .B2(n16650), .C1(
        \registers[19][17] ), .C2(n16647), .A(n11255), .ZN(n11252) );
  AOI211_X1 U8339 ( .C1(\registers[23][17] ), .C2(n16626), .A(n11257), .B(
        n16666), .ZN(n11250) );
  AOI221_X1 U8340 ( .B1(\registers[1][17] ), .B2(n16638), .C1(
        \registers[22][17] ), .C2(n16635), .A(n11256), .ZN(n11251) );
  NAND4_X1 U8341 ( .A1(n11164), .A2(n11165), .A3(n11166), .A4(n11167), .ZN(
        n11163) );
  AOI221_X1 U8342 ( .B1(\registers[16][19] ), .B2(n16650), .C1(
        \registers[19][19] ), .C2(n16647), .A(n11169), .ZN(n11166) );
  AOI211_X1 U8343 ( .C1(\registers[23][19] ), .C2(n16626), .A(n11171), .B(
        n16666), .ZN(n11164) );
  AOI221_X1 U8344 ( .B1(\registers[1][19] ), .B2(n16638), .C1(
        \registers[22][19] ), .C2(n16635), .A(n11170), .ZN(n11165) );
  NAND4_X1 U8345 ( .A1(n11121), .A2(n11122), .A3(n11123), .A4(n11124), .ZN(
        n11120) );
  AOI221_X1 U8346 ( .B1(\registers[16][20] ), .B2(n16650), .C1(
        \registers[19][20] ), .C2(n16647), .A(n11126), .ZN(n11123) );
  AOI211_X1 U8347 ( .C1(\registers[23][20] ), .C2(n16626), .A(n11128), .B(
        n16666), .ZN(n11121) );
  AOI221_X1 U8348 ( .B1(\registers[1][20] ), .B2(n16638), .C1(
        \registers[22][20] ), .C2(n16635), .A(n11127), .ZN(n11122) );
  NAND4_X1 U8349 ( .A1(n11078), .A2(n11079), .A3(n11080), .A4(n11081), .ZN(
        n11077) );
  AOI221_X1 U8350 ( .B1(\registers[16][21] ), .B2(n16650), .C1(
        \registers[19][21] ), .C2(n16647), .A(n11083), .ZN(n11080) );
  AOI211_X1 U8351 ( .C1(\registers[23][21] ), .C2(n16626), .A(n11085), .B(
        n16666), .ZN(n11078) );
  AOI221_X1 U8352 ( .B1(\registers[1][21] ), .B2(n16638), .C1(
        \registers[22][21] ), .C2(n16635), .A(n11084), .ZN(n11079) );
  NAND4_X1 U8353 ( .A1(n11035), .A2(n11036), .A3(n11037), .A4(n11038), .ZN(
        n11034) );
  AOI221_X1 U8354 ( .B1(\registers[16][22] ), .B2(n16650), .C1(
        \registers[19][22] ), .C2(n16647), .A(n11040), .ZN(n11037) );
  AOI211_X1 U8355 ( .C1(\registers[23][22] ), .C2(n16626), .A(n11042), .B(
        n16666), .ZN(n11035) );
  AOI221_X1 U8356 ( .B1(\registers[1][22] ), .B2(n16638), .C1(
        \registers[22][22] ), .C2(n16635), .A(n11041), .ZN(n11036) );
  NAND4_X1 U8357 ( .A1(n10992), .A2(n10993), .A3(n10994), .A4(n10995), .ZN(
        n10991) );
  AOI221_X1 U8358 ( .B1(\registers[16][23] ), .B2(n16650), .C1(
        \registers[19][23] ), .C2(n16647), .A(n10997), .ZN(n10994) );
  AOI211_X1 U8359 ( .C1(\registers[23][23] ), .C2(n16626), .A(n10999), .B(
        n16666), .ZN(n10992) );
  AOI221_X1 U8360 ( .B1(\registers[1][23] ), .B2(n16638), .C1(
        \registers[22][23] ), .C2(n16635), .A(n10998), .ZN(n10993) );
  NAND4_X1 U8361 ( .A1(n10949), .A2(n10950), .A3(n10951), .A4(n10952), .ZN(
        n10948) );
  AOI221_X1 U8362 ( .B1(\registers[16][24] ), .B2(n16651), .C1(
        \registers[19][24] ), .C2(n16648), .A(n10954), .ZN(n10951) );
  AOI211_X1 U8363 ( .C1(\registers[23][24] ), .C2(n16627), .A(n10956), .B(
        n16666), .ZN(n10949) );
  AOI221_X1 U8364 ( .B1(\registers[1][24] ), .B2(n16639), .C1(
        \registers[22][24] ), .C2(n16636), .A(n10955), .ZN(n10950) );
  NAND2_X1 U8365 ( .A1(n14016), .A2(call), .ZN(n14159) );
  NAND2_X1 U8366 ( .A1(n10190), .A2(N9909), .ZN(n14144) );
  INV_X1 U8367 ( .A(N46058), .ZN(n13984) );
  INV_X1 U8368 ( .A(N190), .ZN(n14229) );
  INV_X1 U8369 ( .A(N45544), .ZN(n12503) );
  AND2_X1 U8370 ( .A1(n13987), .A2(N46056), .ZN(n13901) );
  AND2_X1 U8371 ( .A1(n12506), .A2(N45542), .ZN(n12420) );
  NAND2_X1 U8372 ( .A1(n7592), .A2(n14265), .ZN(n14247) );
  OR2_X1 U8373 ( .A1(N190), .A2(N191), .ZN(n14213) );
  NOR2_X1 U8374 ( .A1(n10189), .A2(n14004), .ZN(n10179) );
  NOR2_X1 U8375 ( .A1(n10187), .A2(n14004), .ZN(n10175) );
  NOR2_X1 U8376 ( .A1(n7587), .A2(n14229), .ZN(\add_73/carry[1] ) );
  NOR2_X1 U8377 ( .A1(n10190), .A2(n14004), .ZN(n10180) );
  OAI21_X1 U8378 ( .B1(n5522), .B2(n18049), .A(n13998), .ZN(n10183) );
  NOR2_X1 U8379 ( .A1(n10188), .A2(n14004), .ZN(n10177) );
  AOI22_X1 U8380 ( .A1(net226855), .A2(n16466), .B1(\registers[68][1] ), .B2(
        n16463), .ZN(n12259) );
  AOI221_X1 U8381 ( .B1(net226854), .B2(n16687), .C1(net226853), .C2(n16682), 
        .A(n12262), .ZN(n12261) );
  AOI221_X1 U8382 ( .B1(net226856), .B2(n16675), .C1(net226865), .C2(n16670), 
        .A(n12263), .ZN(n12260) );
  AOI22_X1 U8383 ( .A1(net226876), .A2(n16466), .B1(\registers[68][2] ), .B2(
        n16463), .ZN(n12106) );
  AOI221_X1 U8384 ( .B1(net226874), .B2(n16687), .C1(net226873), .C2(n16682), 
        .A(n12109), .ZN(n12108) );
  AOI221_X1 U8385 ( .B1(net226877), .B2(n16675), .C1(net226875), .C2(n16670), 
        .A(n12110), .ZN(n12107) );
  AOI22_X1 U8386 ( .A1(net226896), .A2(n16466), .B1(\registers[68][3] ), .B2(
        n16463), .ZN(n11953) );
  AOI221_X1 U8387 ( .B1(net226894), .B2(n16687), .C1(net226893), .C2(n16682), 
        .A(n11956), .ZN(n11955) );
  AOI221_X1 U8388 ( .B1(net226897), .B2(n16675), .C1(net226895), .C2(n16670), 
        .A(n11957), .ZN(n11954) );
  AOI22_X1 U8389 ( .A1(n16214), .A2(net226843), .B1(n16213), .B2(
        \registers[68][0] ), .ZN(n13897) );
  AOI221_X1 U8390 ( .B1(n16433), .B2(net226842), .C1(n16430), .C2(net226833), 
        .A(n13900), .ZN(n13899) );
  AOI221_X1 U8391 ( .B1(n16421), .B2(net226835), .C1(n16418), .C2(net226834), 
        .A(n13906), .ZN(n13898) );
  AOI22_X1 U8392 ( .A1(n16214), .A2(net226855), .B1(n16213), .B2(
        \registers[68][1] ), .ZN(n13855) );
  AOI221_X1 U8393 ( .B1(n16433), .B2(net226854), .C1(n16430), .C2(net226853), 
        .A(n13858), .ZN(n13857) );
  AOI221_X1 U8394 ( .B1(n16421), .B2(net226856), .C1(n16418), .C2(net226865), 
        .A(n13859), .ZN(n13856) );
  AOI22_X1 U8395 ( .A1(n16214), .A2(net226876), .B1(n16213), .B2(
        \registers[68][2] ), .ZN(n13813) );
  AOI221_X1 U8396 ( .B1(n16433), .B2(net226874), .C1(n16430), .C2(net226873), 
        .A(n13816), .ZN(n13815) );
  AOI221_X1 U8397 ( .B1(n16421), .B2(net226877), .C1(n16418), .C2(net226875), 
        .A(n13817), .ZN(n13814) );
  AOI22_X1 U8398 ( .A1(n16214), .A2(net226896), .B1(n16213), .B2(
        \registers[68][3] ), .ZN(n13771) );
  AOI221_X1 U8399 ( .B1(n16433), .B2(net226894), .C1(n16430), .C2(net226893), 
        .A(n13774), .ZN(n13773) );
  AOI221_X1 U8400 ( .B1(n16421), .B2(net226897), .C1(n16418), .C2(net226895), 
        .A(n13775), .ZN(n13772) );
  AOI22_X1 U8401 ( .A1(n16214), .A2(net226970), .B1(n16213), .B2(
        \registers[68][4] ), .ZN(n13729) );
  AOI221_X1 U8402 ( .B1(n16433), .B2(net226968), .C1(n16430), .C2(net226967), 
        .A(n13732), .ZN(n13731) );
  AOI221_X1 U8403 ( .B1(n16421), .B2(net226971), .C1(n16418), .C2(net226969), 
        .A(n13733), .ZN(n13730) );
  AOI22_X1 U8404 ( .A1(n16214), .A2(net226988), .B1(n16213), .B2(
        \registers[68][5] ), .ZN(n13687) );
  AOI221_X1 U8405 ( .B1(n16433), .B2(net226986), .C1(n16430), .C2(net226985), 
        .A(n13690), .ZN(n13689) );
  AOI221_X1 U8406 ( .B1(n16421), .B2(net226989), .C1(n16418), .C2(net226987), 
        .A(n13691), .ZN(n13688) );
  AOI22_X1 U8407 ( .A1(n16214), .A2(net227006), .B1(n16213), .B2(
        \registers[68][6] ), .ZN(n13645) );
  AOI221_X1 U8408 ( .B1(n16433), .B2(net227004), .C1(n16430), .C2(net227003), 
        .A(n13648), .ZN(n13647) );
  AOI221_X1 U8409 ( .B1(n16421), .B2(net227007), .C1(n16418), .C2(net227005), 
        .A(n13649), .ZN(n13646) );
  AOI22_X1 U8410 ( .A1(n16214), .A2(net227024), .B1(n16213), .B2(
        \registers[68][7] ), .ZN(n13603) );
  AOI221_X1 U8411 ( .B1(n16433), .B2(net227022), .C1(n16430), .C2(net227021), 
        .A(n13606), .ZN(n13605) );
  AOI221_X1 U8412 ( .B1(n16421), .B2(net227025), .C1(n16418), .C2(net227023), 
        .A(n13607), .ZN(n13604) );
  AOI22_X1 U8413 ( .A1(n16214), .A2(net227042), .B1(n16212), .B2(
        \registers[68][8] ), .ZN(n13561) );
  AOI221_X1 U8414 ( .B1(n16433), .B2(net227040), .C1(n16430), .C2(net227039), 
        .A(n13564), .ZN(n13563) );
  AOI221_X1 U8415 ( .B1(n16421), .B2(net227043), .C1(n16418), .C2(net227041), 
        .A(n13565), .ZN(n13562) );
  AOI22_X1 U8416 ( .A1(n16214), .A2(net227060), .B1(n16212), .B2(
        \registers[68][9] ), .ZN(n13519) );
  AOI221_X1 U8417 ( .B1(n16433), .B2(net227058), .C1(n16430), .C2(net227057), 
        .A(n13522), .ZN(n13521) );
  AOI221_X1 U8418 ( .B1(n16421), .B2(net227061), .C1(n16418), .C2(net227059), 
        .A(n13523), .ZN(n13520) );
  AOI22_X1 U8419 ( .A1(n16214), .A2(net227078), .B1(n16212), .B2(
        \registers[68][10] ), .ZN(n13477) );
  AOI221_X1 U8420 ( .B1(n16433), .B2(net227076), .C1(n16430), .C2(net227075), 
        .A(n13480), .ZN(n13479) );
  AOI221_X1 U8421 ( .B1(n16421), .B2(net227079), .C1(n16418), .C2(net227077), 
        .A(n13481), .ZN(n13478) );
  AOI22_X1 U8422 ( .A1(n16214), .A2(net227096), .B1(n16212), .B2(
        \registers[68][11] ), .ZN(n13435) );
  AOI221_X1 U8423 ( .B1(n16433), .B2(net227094), .C1(n16430), .C2(net227093), 
        .A(n13438), .ZN(n13437) );
  AOI221_X1 U8424 ( .B1(n16421), .B2(net227097), .C1(n16418), .C2(net227095), 
        .A(n13439), .ZN(n13436) );
  AOI22_X1 U8425 ( .A1(n16215), .A2(net227114), .B1(n16212), .B2(
        \registers[68][12] ), .ZN(n13393) );
  AOI221_X1 U8426 ( .B1(n16434), .B2(net227112), .C1(n16431), .C2(net227111), 
        .A(n13396), .ZN(n13395) );
  AOI221_X1 U8427 ( .B1(n16422), .B2(net227115), .C1(n16419), .C2(net227113), 
        .A(n13397), .ZN(n13394) );
  AOI22_X1 U8428 ( .A1(n16215), .A2(net227132), .B1(n16212), .B2(
        \registers[68][13] ), .ZN(n13351) );
  AOI221_X1 U8429 ( .B1(n16434), .B2(net227130), .C1(n16431), .C2(net227129), 
        .A(n13354), .ZN(n13353) );
  AOI221_X1 U8430 ( .B1(n16422), .B2(net227133), .C1(n16419), .C2(net227131), 
        .A(n13355), .ZN(n13352) );
  AOI22_X1 U8431 ( .A1(n16215), .A2(net227150), .B1(n16212), .B2(
        \registers[68][14] ), .ZN(n13309) );
  AOI221_X1 U8432 ( .B1(n16434), .B2(net227148), .C1(n16431), .C2(net227147), 
        .A(n13312), .ZN(n13311) );
  AOI221_X1 U8433 ( .B1(n16422), .B2(net227151), .C1(n16419), .C2(net227149), 
        .A(n13313), .ZN(n13310) );
  AOI22_X1 U8434 ( .A1(n16215), .A2(net227168), .B1(n16212), .B2(
        \registers[68][15] ), .ZN(n13267) );
  AOI221_X1 U8435 ( .B1(n16434), .B2(net227166), .C1(n16431), .C2(net227165), 
        .A(n13270), .ZN(n13269) );
  AOI221_X1 U8436 ( .B1(n16422), .B2(net227169), .C1(n16419), .C2(net227167), 
        .A(n13271), .ZN(n13268) );
  AOI22_X1 U8437 ( .A1(n16215), .A2(net227186), .B1(n16212), .B2(
        \registers[68][16] ), .ZN(n13225) );
  AOI221_X1 U8438 ( .B1(n16434), .B2(net227184), .C1(n16431), .C2(net227183), 
        .A(n13228), .ZN(n13227) );
  AOI221_X1 U8439 ( .B1(n16422), .B2(net227187), .C1(n16419), .C2(net227185), 
        .A(n13229), .ZN(n13226) );
  AOI22_X1 U8440 ( .A1(n16215), .A2(net227204), .B1(n16212), .B2(
        \registers[68][17] ), .ZN(n13183) );
  AOI221_X1 U8441 ( .B1(n16434), .B2(net227202), .C1(n16431), .C2(net227201), 
        .A(n13186), .ZN(n13185) );
  AOI221_X1 U8442 ( .B1(n16422), .B2(net227205), .C1(n16419), .C2(net227203), 
        .A(n13187), .ZN(n13184) );
  AOI22_X1 U8443 ( .A1(n16215), .A2(net227222), .B1(n16212), .B2(
        \registers[68][18] ), .ZN(n13141) );
  AOI221_X1 U8444 ( .B1(n16434), .B2(net227220), .C1(n16431), .C2(net227219), 
        .A(n13144), .ZN(n13143) );
  AOI221_X1 U8445 ( .B1(n16422), .B2(net227223), .C1(n16419), .C2(net227221), 
        .A(n13145), .ZN(n13142) );
  AOI22_X1 U8446 ( .A1(n16215), .A2(net227240), .B1(n16212), .B2(
        \registers[68][19] ), .ZN(n13099) );
  AOI221_X1 U8447 ( .B1(n16434), .B2(net227238), .C1(n16431), .C2(net227237), 
        .A(n13102), .ZN(n13101) );
  AOI221_X1 U8448 ( .B1(n16422), .B2(net227241), .C1(n16419), .C2(net227239), 
        .A(n13103), .ZN(n13100) );
  AOI22_X1 U8449 ( .A1(n16215), .A2(net227258), .B1(n16211), .B2(
        \registers[68][20] ), .ZN(n13057) );
  AOI221_X1 U8450 ( .B1(n16434), .B2(net227256), .C1(n16431), .C2(net227255), 
        .A(n13060), .ZN(n13059) );
  AOI221_X1 U8451 ( .B1(n16422), .B2(net227259), .C1(n16419), .C2(net227257), 
        .A(n13061), .ZN(n13058) );
  AOI22_X1 U8452 ( .A1(n16215), .A2(net227276), .B1(n16211), .B2(
        \registers[68][21] ), .ZN(n13015) );
  AOI221_X1 U8453 ( .B1(n16434), .B2(net227274), .C1(n16431), .C2(net227273), 
        .A(n13018), .ZN(n13017) );
  AOI221_X1 U8454 ( .B1(n16422), .B2(net227277), .C1(n16419), .C2(net227275), 
        .A(n13019), .ZN(n13016) );
  AOI22_X1 U8455 ( .A1(n16215), .A2(net227294), .B1(n16211), .B2(
        \registers[68][22] ), .ZN(n12973) );
  AOI221_X1 U8456 ( .B1(n16434), .B2(net227292), .C1(n16431), .C2(net227291), 
        .A(n12976), .ZN(n12975) );
  AOI221_X1 U8457 ( .B1(n16422), .B2(net227295), .C1(n16419), .C2(net227293), 
        .A(n12977), .ZN(n12974) );
  AOI22_X1 U8458 ( .A1(n16215), .A2(net227312), .B1(n16211), .B2(
        \registers[68][23] ), .ZN(n12931) );
  AOI221_X1 U8459 ( .B1(n16434), .B2(net227310), .C1(n16431), .C2(net227309), 
        .A(n12934), .ZN(n12933) );
  AOI221_X1 U8460 ( .B1(n16422), .B2(net227313), .C1(n16419), .C2(net227311), 
        .A(n12935), .ZN(n12932) );
  AOI22_X1 U8461 ( .A1(n16466), .A2(net226970), .B1(n16463), .B2(
        \registers[68][4] ), .ZN(n11800) );
  AOI221_X1 U8462 ( .B1(n16687), .B2(net226968), .C1(n16682), .C2(net226967), 
        .A(n11803), .ZN(n11802) );
  AOI221_X1 U8463 ( .B1(n16675), .B2(net226971), .C1(n16670), .C2(net226969), 
        .A(n11804), .ZN(n11801) );
  AOI22_X1 U8464 ( .A1(n16468), .A2(net227024), .B1(n16465), .B2(
        \registers[68][7] ), .ZN(n11671) );
  AOI221_X1 U8465 ( .B1(n16686), .B2(net227022), .C1(n16684), .C2(net227021), 
        .A(n11674), .ZN(n11673) );
  AOI221_X1 U8466 ( .B1(n16674), .B2(net227025), .C1(n16672), .C2(net227023), 
        .A(n11675), .ZN(n11672) );
  AOI22_X1 U8467 ( .A1(n16468), .A2(net227042), .B1(n16465), .B2(
        \registers[68][8] ), .ZN(n11628) );
  AOI221_X1 U8468 ( .B1(n16686), .B2(net227040), .C1(n16684), .C2(net227039), 
        .A(n11631), .ZN(n11630) );
  AOI221_X1 U8469 ( .B1(n16674), .B2(net227043), .C1(n16672), .C2(net227041), 
        .A(n11632), .ZN(n11629) );
  AOI22_X1 U8470 ( .A1(n16468), .A2(net227060), .B1(n16465), .B2(
        \registers[68][9] ), .ZN(n11585) );
  AOI221_X1 U8471 ( .B1(n16686), .B2(net227058), .C1(n16684), .C2(net227057), 
        .A(n11588), .ZN(n11587) );
  AOI221_X1 U8472 ( .B1(n16674), .B2(net227061), .C1(n16672), .C2(net227059), 
        .A(n11589), .ZN(n11586) );
  AOI22_X1 U8473 ( .A1(n16468), .A2(net227078), .B1(n16465), .B2(
        \registers[68][10] ), .ZN(n11542) );
  AOI221_X1 U8474 ( .B1(n16686), .B2(net227076), .C1(n16684), .C2(net227075), 
        .A(n11545), .ZN(n11544) );
  AOI221_X1 U8475 ( .B1(n16674), .B2(net227079), .C1(n16672), .C2(net227077), 
        .A(n11546), .ZN(n11543) );
  AOI22_X1 U8476 ( .A1(n16467), .A2(net227096), .B1(n16464), .B2(
        \registers[68][11] ), .ZN(n11499) );
  AOI221_X1 U8477 ( .B1(n16686), .B2(net227094), .C1(n16683), .C2(net227093), 
        .A(n11502), .ZN(n11501) );
  AOI221_X1 U8478 ( .B1(n16674), .B2(net227097), .C1(n16671), .C2(net227095), 
        .A(n11503), .ZN(n11500) );
  AOI22_X1 U8479 ( .A1(n16467), .A2(net227114), .B1(n16464), .B2(
        \registers[68][12] ), .ZN(n11455) );
  AOI221_X1 U8480 ( .B1(n16686), .B2(net227112), .C1(n16683), .C2(net227111), 
        .A(n11458), .ZN(n11457) );
  AOI221_X1 U8481 ( .B1(n16674), .B2(net227115), .C1(n16671), .C2(net227113), 
        .A(n11459), .ZN(n11456) );
  AOI22_X1 U8482 ( .A1(n16467), .A2(net227132), .B1(n16464), .B2(
        \registers[68][13] ), .ZN(n11412) );
  AOI221_X1 U8483 ( .B1(n16686), .B2(net227130), .C1(n16683), .C2(net227129), 
        .A(n11415), .ZN(n11414) );
  AOI221_X1 U8484 ( .B1(n16674), .B2(net227133), .C1(n16671), .C2(net227131), 
        .A(n11416), .ZN(n11413) );
  AOI22_X1 U8485 ( .A1(n16467), .A2(net227150), .B1(n16464), .B2(
        \registers[68][14] ), .ZN(n11369) );
  AOI221_X1 U8486 ( .B1(n16686), .B2(net227148), .C1(n16683), .C2(net227147), 
        .A(n11372), .ZN(n11371) );
  AOI221_X1 U8487 ( .B1(n16674), .B2(net227151), .C1(n16671), .C2(net227149), 
        .A(n11373), .ZN(n11370) );
  AOI22_X1 U8488 ( .A1(n16467), .A2(net227168), .B1(n16464), .B2(
        \registers[68][15] ), .ZN(n11326) );
  AOI221_X1 U8489 ( .B1(n16686), .B2(net227166), .C1(n16683), .C2(net227165), 
        .A(n11329), .ZN(n11328) );
  AOI221_X1 U8490 ( .B1(n16674), .B2(net227169), .C1(n16671), .C2(net227167), 
        .A(n11330), .ZN(n11327) );
  AOI22_X1 U8491 ( .A1(n16467), .A2(net227186), .B1(n16464), .B2(
        \registers[68][16] ), .ZN(n11283) );
  AOI221_X1 U8492 ( .B1(n16686), .B2(net227184), .C1(n16683), .C2(net227183), 
        .A(n11286), .ZN(n11285) );
  AOI221_X1 U8493 ( .B1(n16674), .B2(net227187), .C1(n16671), .C2(net227185), 
        .A(n11287), .ZN(n11284) );
  AOI22_X1 U8494 ( .A1(n16467), .A2(net227204), .B1(n16464), .B2(
        \registers[68][17] ), .ZN(n11240) );
  AOI221_X1 U8495 ( .B1(n16686), .B2(net227202), .C1(n16683), .C2(net227201), 
        .A(n11243), .ZN(n11242) );
  AOI221_X1 U8496 ( .B1(n16674), .B2(net227205), .C1(n16671), .C2(net227203), 
        .A(n11244), .ZN(n11241) );
  AOI22_X1 U8497 ( .A1(n16467), .A2(net227222), .B1(n16464), .B2(
        \registers[68][18] ), .ZN(n11197) );
  AOI221_X1 U8498 ( .B1(n16685), .B2(net227220), .C1(n16683), .C2(net227219), 
        .A(n11200), .ZN(n11199) );
  AOI221_X1 U8499 ( .B1(n16673), .B2(net227223), .C1(n16671), .C2(net227221), 
        .A(n11201), .ZN(n11198) );
  AOI22_X1 U8500 ( .A1(n16467), .A2(net227240), .B1(n16464), .B2(
        \registers[68][19] ), .ZN(n11154) );
  AOI221_X1 U8501 ( .B1(n16685), .B2(net227238), .C1(n16683), .C2(net227237), 
        .A(n11157), .ZN(n11156) );
  AOI221_X1 U8502 ( .B1(n16673), .B2(net227241), .C1(n16671), .C2(net227239), 
        .A(n11158), .ZN(n11155) );
  AOI22_X1 U8503 ( .A1(n16467), .A2(net227258), .B1(n16464), .B2(
        \registers[68][20] ), .ZN(n11111) );
  AOI221_X1 U8504 ( .B1(n16685), .B2(net227256), .C1(n16683), .C2(net227255), 
        .A(n11114), .ZN(n11113) );
  AOI221_X1 U8505 ( .B1(n16673), .B2(net227259), .C1(n16671), .C2(net227257), 
        .A(n11115), .ZN(n11112) );
  AOI22_X1 U8506 ( .A1(n16467), .A2(net227276), .B1(n16464), .B2(
        \registers[68][21] ), .ZN(n11068) );
  AOI221_X1 U8507 ( .B1(n16685), .B2(net227274), .C1(n16683), .C2(net227273), 
        .A(n11071), .ZN(n11070) );
  AOI221_X1 U8508 ( .B1(n16673), .B2(net227277), .C1(n16671), .C2(net227275), 
        .A(n11072), .ZN(n11069) );
  AOI22_X1 U8509 ( .A1(n16467), .A2(net227294), .B1(n16464), .B2(
        \registers[68][22] ), .ZN(n11025) );
  AOI221_X1 U8510 ( .B1(n16685), .B2(net227292), .C1(n16683), .C2(net227291), 
        .A(n11028), .ZN(n11027) );
  AOI221_X1 U8511 ( .B1(n16673), .B2(net227295), .C1(n16671), .C2(net227293), 
        .A(n11029), .ZN(n11026) );
  AOI22_X1 U8512 ( .A1(n16467), .A2(net227312), .B1(n16464), .B2(
        \registers[68][23] ), .ZN(n10982) );
  AOI221_X1 U8513 ( .B1(n16686), .B2(net227310), .C1(n16683), .C2(net227309), 
        .A(n10985), .ZN(n10984) );
  AOI221_X1 U8514 ( .B1(n16674), .B2(net227313), .C1(n16671), .C2(net227311), 
        .A(n10986), .ZN(n10983) );
  AOI22_X1 U8515 ( .A1(n16466), .A2(net227330), .B1(n16463), .B2(
        \registers[68][24] ), .ZN(n10939) );
  AOI221_X1 U8516 ( .B1(n16685), .B2(net227328), .C1(n16682), .C2(net227327), 
        .A(n10942), .ZN(n10941) );
  AOI221_X1 U8517 ( .B1(n16673), .B2(net227331), .C1(n16670), .C2(net227329), 
        .A(n10943), .ZN(n10940) );
  AOI22_X1 U8518 ( .A1(n16466), .A2(net227348), .B1(n16463), .B2(
        \registers[68][25] ), .ZN(n10896) );
  AOI221_X1 U8519 ( .B1(n16685), .B2(net227346), .C1(n16682), .C2(net227345), 
        .A(n10899), .ZN(n10898) );
  AOI221_X1 U8520 ( .B1(n16673), .B2(net227349), .C1(n16670), .C2(net227347), 
        .A(n10900), .ZN(n10897) );
  AOI22_X1 U8521 ( .A1(n16466), .A2(net227366), .B1(n16463), .B2(
        \registers[68][26] ), .ZN(n10853) );
  AOI221_X1 U8522 ( .B1(n16685), .B2(net227364), .C1(n16682), .C2(net227363), 
        .A(n10856), .ZN(n10855) );
  AOI221_X1 U8523 ( .B1(n16673), .B2(net227367), .C1(n16670), .C2(net227365), 
        .A(n10857), .ZN(n10854) );
  AOI22_X1 U8524 ( .A1(n16466), .A2(net227384), .B1(n16463), .B2(
        \registers[68][27] ), .ZN(n10810) );
  AOI221_X1 U8525 ( .B1(n16685), .B2(net227382), .C1(n16682), .C2(net227381), 
        .A(n10813), .ZN(n10812) );
  AOI221_X1 U8526 ( .B1(n16673), .B2(net227385), .C1(n16670), .C2(net227383), 
        .A(n10814), .ZN(n10811) );
  AOI22_X1 U8527 ( .A1(n16466), .A2(net227402), .B1(n16463), .B2(
        \registers[68][28] ), .ZN(n10767) );
  AOI221_X1 U8528 ( .B1(n16685), .B2(net227400), .C1(n16682), .C2(net227399), 
        .A(n10770), .ZN(n10769) );
  AOI221_X1 U8529 ( .B1(n16673), .B2(net227403), .C1(n16670), .C2(net227401), 
        .A(n10771), .ZN(n10768) );
  AOI22_X1 U8530 ( .A1(n16466), .A2(net227420), .B1(n16463), .B2(
        \registers[68][29] ), .ZN(n10724) );
  AOI221_X1 U8531 ( .B1(n16685), .B2(net227418), .C1(n16682), .C2(net227417), 
        .A(n10727), .ZN(n10726) );
  AOI221_X1 U8532 ( .B1(n16673), .B2(net227421), .C1(n16670), .C2(net227419), 
        .A(n10728), .ZN(n10725) );
  AOI22_X1 U8533 ( .A1(n16466), .A2(net227438), .B1(n16463), .B2(
        \registers[68][30] ), .ZN(n10665) );
  AOI221_X1 U8534 ( .B1(n16685), .B2(net227436), .C1(n16682), .C2(net227435), 
        .A(n10668), .ZN(n10667) );
  AOI221_X1 U8535 ( .B1(n16673), .B2(net227439), .C1(n16670), .C2(net227437), 
        .A(n10669), .ZN(n10666) );
  AND4_X1 U8536 ( .A1(n14233), .A2(wr), .A3(\sub_71/carry[4] ), .A4(add_wr[4]), 
        .ZN(n14223) );
  AND2_X1 U8537 ( .A1(n14016), .A2(\r590/carry[5] ), .ZN(n14194) );
  NOR4_X1 U8538 ( .A1(n13989), .A2(N46056), .A3(add_rd2[4]), .A4(
        \sub_146/carry[4] ), .ZN(n13974) );
  INV_X1 U8539 ( .A(n13985), .ZN(n13989) );
  AND4_X1 U8540 ( .A1(n14026), .A2(n14027), .A3(n14028), .A4(n14029), .ZN(
        n14024) );
  XNOR2_X1 U8541 ( .A(swp[2]), .B(N9909), .ZN(n14027) );
  XNOR2_X1 U8542 ( .A(swp[0]), .B(N9641), .ZN(n14026) );
  XNOR2_X1 U8543 ( .A(swp[3]), .B(N9910), .ZN(n14028) );
  NOR4_X1 U8544 ( .A1(n12508), .A2(N45542), .A3(add_rd1[4]), .A4(
        \sub_132/carry[4] ), .ZN(n12493) );
  INV_X1 U8545 ( .A(n12504), .ZN(n12508) );
  INV_X1 U8546 ( .A(n11859), .ZN(n8037) );
  AOI221_X1 U8547 ( .B1(n17989), .B2(\registers[56][3] ), .C1(n17991), .C2(
        datain[3]), .A(n18049), .ZN(n11859) );
  INV_X1 U8548 ( .A(n11853), .ZN(n8043) );
  AOI221_X1 U8549 ( .B1(n16989), .B2(\registers[42][3] ), .C1(n16991), .C2(
        datain[3]), .A(n18049), .ZN(n11853) );
  INV_X1 U8550 ( .A(n11848), .ZN(n8048) );
  AOI221_X1 U8551 ( .B1(n17150), .B2(\registers[29][3] ), .C1(n17152), .C2(
        datain[3]), .A(n18048), .ZN(n11848) );
  INV_X1 U8552 ( .A(n10448), .ZN(n8134) );
  AOI221_X1 U8553 ( .B1(n17216), .B2(\registers[23][4] ), .C1(n17218), .C2(
        datain[4]), .A(n18048), .ZN(n10448) );
  INV_X1 U8554 ( .A(n10444), .ZN(n8138) );
  AOI221_X1 U8555 ( .B1(n17268), .B2(\registers[19][4] ), .C1(n17270), .C2(
        datain[4]), .A(n18048), .ZN(n10444) );
  INV_X1 U8556 ( .A(n10416), .ZN(n8165) );
  AOI221_X1 U8557 ( .B1(n17989), .B2(\registers[56][4] ), .C1(n17992), .C2(
        datain[4]), .A(n18048), .ZN(n10416) );
  INV_X1 U8558 ( .A(n10413), .ZN(n8168) );
  AOI221_X1 U8559 ( .B1(n16866), .B2(net226980), .C1(n16868), .C2(datain[4]), 
        .A(n18047), .ZN(n10413) );
  INV_X1 U8560 ( .A(n10410), .ZN(n8171) );
  AOI221_X1 U8561 ( .B1(n16900), .B2(\registers[50][4] ), .C1(n16902), .C2(
        datain[4]), .A(n18047), .ZN(n10410) );
  INV_X1 U8562 ( .A(n10405), .ZN(n8176) );
  AOI221_X1 U8563 ( .B1(n17150), .B2(\registers[29][4] ), .C1(n17152), .C2(
        datain[4]), .A(n18047), .ZN(n10405) );
  INV_X1 U8564 ( .A(n10306), .ZN(n8237) );
  AOI221_X1 U8565 ( .B1(n17989), .B2(\registers[56][5] ), .C1(n17991), .C2(
        datain[5]), .A(n18047), .ZN(n10306) );
  INV_X1 U8566 ( .A(n10303), .ZN(n8240) );
  AOI221_X1 U8567 ( .B1(n16866), .B2(net227000), .C1(n16868), .C2(datain[5]), 
        .A(n18046), .ZN(n10303) );
  INV_X1 U8568 ( .A(n10300), .ZN(n8243) );
  AOI221_X1 U8569 ( .B1(n16900), .B2(\registers[50][5] ), .C1(n16902), .C2(
        datain[5]), .A(n18046), .ZN(n10300) );
  INV_X1 U8570 ( .A(n10292), .ZN(n8251) );
  AOI221_X1 U8571 ( .B1(n16989), .B2(\registers[42][5] ), .C1(n16991), .C2(
        datain[5]), .A(n18046), .ZN(n10292) );
  INV_X1 U8572 ( .A(n10288), .ZN(n8254) );
  AOI221_X1 U8573 ( .B1(n17534), .B2(net227003), .C1(n17536), .C2(datain[6]), 
        .A(n18046), .ZN(n10288) );
  INV_X1 U8574 ( .A(n10287), .ZN(n8255) );
  AOI221_X1 U8575 ( .B1(n17548), .B2(net227004), .C1(n17550), .C2(datain[6]), 
        .A(n18045), .ZN(n10287) );
  INV_X1 U8576 ( .A(n10286), .ZN(n8256) );
  AOI221_X1 U8577 ( .B1(n17562), .B2(\registers[68][6] ), .C1(n17564), .C2(
        datain[6]), .A(n18045), .ZN(n10286) );
  INV_X1 U8578 ( .A(n10283), .ZN(n8258) );
  AOI221_X1 U8579 ( .B1(n17589), .B2(net227005), .C1(n17591), .C2(datain[6]), 
        .A(n18045), .ZN(n10283) );
  INV_X1 U8580 ( .A(n10282), .ZN(n8259) );
  AOI221_X1 U8581 ( .B1(n17603), .B2(net227006), .C1(n17605), .C2(datain[6]), 
        .A(n18045), .ZN(n10282) );
  INV_X1 U8582 ( .A(n10280), .ZN(n8260) );
  AOI221_X1 U8583 ( .B1(n17617), .B2(net227007), .C1(n17619), .C2(datain[6]), 
        .A(n18049), .ZN(n10280) );
  NOR2_X1 U8584 ( .A1(n10187), .A2(n14017), .ZN(n14021) );
  OAI22_X1 U8585 ( .A1(n14820), .A2(n14000), .B1(\r590/carry[5] ), .B2(n14001), 
        .ZN(n10182) );
  OAI22_X1 U8586 ( .A1(n3043), .A2(n14000), .B1(n14002), .B2(n14001), .ZN(
        n10181) );
  NOR2_X1 U8587 ( .A1(call), .A2(n14003), .ZN(n14002) );
  NOR2_X1 U8588 ( .A1(\r590/carry[5] ), .A2(n14021), .ZN(n14011) );
  NAND2_X1 U8589 ( .A1(N191), .A2(n14229), .ZN(n14220) );
  NAND2_X1 U8590 ( .A1(N191), .A2(N190), .ZN(n12412) );
  NOR2_X1 U8591 ( .A1(n13984), .A2(N46057), .ZN(n13905) );
  NOR2_X1 U8592 ( .A1(n12503), .A2(N45543), .ZN(n12424) );
  AND2_X1 U8593 ( .A1(N46057), .A2(n13984), .ZN(n13902) );
  AND2_X1 U8594 ( .A1(N46057), .A2(N46058), .ZN(n13903) );
  AND2_X1 U8595 ( .A1(N45543), .A2(n12503), .ZN(n12421) );
  OR2_X1 U8596 ( .A1(n14229), .A2(N191), .ZN(n14217) );
  AND2_X1 U8597 ( .A1(N45543), .A2(N45544), .ZN(n12422) );
  NAND2_X1 U8598 ( .A1(n7685), .A2(n17823), .ZN(n10148) );
  NAND2_X1 U8599 ( .A1(n7684), .A2(n17823), .ZN(n10149) );
  NAND2_X1 U8600 ( .A1(n7683), .A2(n17823), .ZN(n10150) );
  NAND2_X1 U8601 ( .A1(n7682), .A2(n17823), .ZN(n10151) );
  NAND2_X1 U8602 ( .A1(n7681), .A2(n17823), .ZN(n10152) );
  NAND2_X1 U8603 ( .A1(n7680), .A2(n17823), .ZN(n10153) );
  NAND2_X1 U8604 ( .A1(n7679), .A2(n17823), .ZN(n10154) );
  NAND2_X1 U8605 ( .A1(n7678), .A2(n17823), .ZN(n10155) );
  NAND2_X1 U8606 ( .A1(n7677), .A2(n17823), .ZN(n10156) );
  NAND2_X1 U8607 ( .A1(n7676), .A2(n17823), .ZN(n10157) );
  NAND2_X1 U8608 ( .A1(n7675), .A2(n17823), .ZN(n10158) );
  NAND2_X1 U8609 ( .A1(n7674), .A2(n17823), .ZN(n10159) );
  NAND2_X1 U8610 ( .A1(n7673), .A2(n17825), .ZN(n10160) );
  NAND2_X1 U8611 ( .A1(n7672), .A2(n17825), .ZN(n10161) );
  NAND2_X1 U8612 ( .A1(n7671), .A2(n17825), .ZN(n10162) );
  NAND2_X1 U8613 ( .A1(n7670), .A2(n17825), .ZN(n10163) );
  NAND2_X1 U8614 ( .A1(n7669), .A2(n17825), .ZN(n10164) );
  NAND2_X1 U8615 ( .A1(n7668), .A2(n17825), .ZN(n10165) );
  NAND2_X1 U8616 ( .A1(n7667), .A2(n17825), .ZN(n10166) );
  NAND2_X1 U8617 ( .A1(n7666), .A2(n17825), .ZN(n10167) );
  NAND2_X1 U8618 ( .A1(n7665), .A2(n17825), .ZN(n10168) );
  NAND2_X1 U8619 ( .A1(n7664), .A2(n17825), .ZN(n10169) );
  NAND2_X1 U8620 ( .A1(n7663), .A2(n17824), .ZN(n10170) );
  NAND2_X1 U8621 ( .A1(n7662), .A2(n17824), .ZN(n10171) );
  NAND2_X1 U8622 ( .A1(n7693), .A2(n17824), .ZN(n10140) );
  NAND2_X1 U8623 ( .A1(n7692), .A2(n17824), .ZN(n10141) );
  NAND2_X1 U8624 ( .A1(n7691), .A2(n17824), .ZN(n10142) );
  NAND2_X1 U8625 ( .A1(n7690), .A2(n17824), .ZN(n10143) );
  NAND2_X1 U8626 ( .A1(n7689), .A2(n17824), .ZN(n10144) );
  NAND2_X1 U8627 ( .A1(n7688), .A2(n17824), .ZN(n10145) );
  NAND2_X1 U8628 ( .A1(n7687), .A2(n17824), .ZN(n10146) );
  NAND2_X1 U8629 ( .A1(n7686), .A2(n17824), .ZN(n10147) );
  OR2_X1 U8630 ( .A1(n18050), .A2(swp[5]), .ZN(n10173) );
  AND2_X1 U8631 ( .A1(n18044), .A2(swp[4]), .ZN(n10172) );
  AND2_X1 U8632 ( .A1(n18044), .A2(swp[3]), .ZN(n10174) );
  AND2_X1 U8633 ( .A1(n18044), .A2(swp[2]), .ZN(n10176) );
  AND2_X1 U8634 ( .A1(n18044), .A2(swp[1]), .ZN(n10178) );
  AND2_X1 U8635 ( .A1(n18044), .A2(swp[0]), .ZN(n10184) );
  INV_X1 U8636 ( .A(call), .ZN(n14020) );
  INV_X1 U8637 ( .A(wr), .ZN(n12514) );
  NOR2_X1 U8638 ( .A1(ret), .A2(call), .ZN(n14005) );
  NAND3_X2 U8639 ( .A1(n14240), .A2(n14239), .A3(N276), .ZN(n14241) );
  CLKBUF_X1 U8640 ( .A(n12527), .Z(n16417) );
  CLKBUF_X1 U8641 ( .A(n10525), .Z(n16669) );
  INV_X1 U8642 ( .A(n16696), .ZN(n16692) );
  CLKBUF_X1 U8643 ( .A(n7652), .Z(n16730) );
  INV_X1 U8644 ( .A(n17455), .ZN(n17451) );
  INV_X1 U8645 ( .A(n17581), .ZN(n17577) );
  INV_X1 U8646 ( .A(n17834), .ZN(n17825) );
  INV_X1 U8647 ( .A(n17855), .ZN(n17838) );
  CLKBUF_X1 U8648 ( .A(n17854), .Z(n17839) );
  CLKBUF_X1 U8649 ( .A(n17856), .Z(n17840) );
  CLKBUF_X1 U8650 ( .A(n17856), .Z(n17841) );
  CLKBUF_X1 U8651 ( .A(n17856), .Z(n17842) );
  CLKBUF_X1 U8652 ( .A(n17856), .Z(n17843) );
  CLKBUF_X1 U8653 ( .A(n17856), .Z(n17844) );
  CLKBUF_X1 U8654 ( .A(n17856), .Z(n17845) );
  CLKBUF_X1 U8655 ( .A(n17856), .Z(n17846) );
  CLKBUF_X1 U8656 ( .A(n17853), .Z(n17847) );
  CLKBUF_X1 U8657 ( .A(n17840), .Z(n17848) );
  CLKBUF_X1 U8658 ( .A(n17845), .Z(n17849) );
  CLKBUF_X1 U8659 ( .A(n17856), .Z(n17850) );
  CLKBUF_X1 U8660 ( .A(n17856), .Z(n17851) );
  CLKBUF_X1 U8661 ( .A(n17856), .Z(n17852) );
  CLKBUF_X1 U8662 ( .A(n17856), .Z(n17853) );
  CLKBUF_X1 U8663 ( .A(n17856), .Z(n17854) );
  CLKBUF_X1 U8664 ( .A(n17856), .Z(n17855) );
  INV_X1 U8665 ( .A(n17835), .ZN(n17856) );
  INV_X1 U8666 ( .A(n17877), .ZN(n17860) );
  CLKBUF_X1 U8667 ( .A(n17878), .Z(n17861) );
  CLKBUF_X1 U8668 ( .A(n17878), .Z(n17862) );
  CLKBUF_X1 U8669 ( .A(n17878), .Z(n17863) );
  CLKBUF_X1 U8670 ( .A(n17878), .Z(n17864) );
  CLKBUF_X1 U8671 ( .A(n17878), .Z(n17865) );
  CLKBUF_X1 U8672 ( .A(n17878), .Z(n17866) );
  CLKBUF_X1 U8673 ( .A(n17865), .Z(n17867) );
  CLKBUF_X1 U8674 ( .A(n17861), .Z(n17868) );
  CLKBUF_X1 U8675 ( .A(n17866), .Z(n17869) );
  CLKBUF_X1 U8676 ( .A(n17864), .Z(n17870) );
  CLKBUF_X1 U8677 ( .A(n17876), .Z(n17871) );
  CLKBUF_X1 U8678 ( .A(n17878), .Z(n17872) );
  CLKBUF_X1 U8679 ( .A(n17878), .Z(n17873) );
  CLKBUF_X1 U8680 ( .A(n17878), .Z(n17874) );
  CLKBUF_X1 U8681 ( .A(n17863), .Z(n17875) );
  CLKBUF_X1 U8682 ( .A(n17878), .Z(n17876) );
  CLKBUF_X1 U8683 ( .A(n17878), .Z(n17877) );
  INV_X1 U8684 ( .A(n17857), .ZN(n17878) );
  INV_X1 U8685 ( .A(n17899), .ZN(n17882) );
  CLKBUF_X1 U8686 ( .A(n17900), .Z(n17883) );
  CLKBUF_X1 U8687 ( .A(n17887), .Z(n17884) );
  CLKBUF_X1 U8688 ( .A(n17900), .Z(n17885) );
  CLKBUF_X1 U8689 ( .A(n17900), .Z(n17886) );
  CLKBUF_X1 U8690 ( .A(n17900), .Z(n17887) );
  CLKBUF_X1 U8691 ( .A(n17900), .Z(n17888) );
  CLKBUF_X1 U8692 ( .A(n17900), .Z(n17889) );
  CLKBUF_X1 U8693 ( .A(n17900), .Z(n17890) );
  CLKBUF_X1 U8694 ( .A(n17888), .Z(n17891) );
  CLKBUF_X1 U8695 ( .A(n17890), .Z(n17892) );
  CLKBUF_X1 U8696 ( .A(n17883), .Z(n17893) );
  CLKBUF_X1 U8697 ( .A(n17900), .Z(n17894) );
  CLKBUF_X1 U8698 ( .A(n17898), .Z(n17895) );
  CLKBUF_X1 U8699 ( .A(n17900), .Z(n17896) );
  CLKBUF_X1 U8700 ( .A(n17889), .Z(n17897) );
  CLKBUF_X1 U8701 ( .A(n17900), .Z(n17898) );
  CLKBUF_X1 U8702 ( .A(n17900), .Z(n17899) );
  INV_X1 U8703 ( .A(n17879), .ZN(n17900) );
  INV_X1 U8704 ( .A(n17921), .ZN(n17904) );
  CLKBUF_X1 U8705 ( .A(n17922), .Z(n17905) );
  CLKBUF_X1 U8706 ( .A(n17922), .Z(n17906) );
  CLKBUF_X1 U8707 ( .A(n17922), .Z(n17907) );
  CLKBUF_X1 U8708 ( .A(n17922), .Z(n17908) );
  CLKBUF_X1 U8709 ( .A(n17922), .Z(n17909) );
  CLKBUF_X1 U8710 ( .A(n17922), .Z(n17910) );
  CLKBUF_X1 U8711 ( .A(n17909), .Z(n17911) );
  CLKBUF_X1 U8712 ( .A(n17905), .Z(n17912) );
  CLKBUF_X1 U8713 ( .A(n17910), .Z(n17913) );
  CLKBUF_X1 U8714 ( .A(n17908), .Z(n17914) );
  CLKBUF_X1 U8715 ( .A(n17920), .Z(n17915) );
  CLKBUF_X1 U8716 ( .A(n17922), .Z(n17916) );
  CLKBUF_X1 U8717 ( .A(n17922), .Z(n17917) );
  CLKBUF_X1 U8718 ( .A(n17922), .Z(n17918) );
  CLKBUF_X1 U8719 ( .A(n17907), .Z(n17919) );
  CLKBUF_X1 U8720 ( .A(n17922), .Z(n17920) );
  CLKBUF_X1 U8721 ( .A(n17922), .Z(n17921) );
  INV_X1 U8722 ( .A(n17901), .ZN(n17922) );
  INV_X1 U8723 ( .A(n17942), .ZN(n17925) );
  CLKBUF_X1 U8724 ( .A(n17943), .Z(n17926) );
  CLKBUF_X1 U8725 ( .A(n17930), .Z(n17927) );
  CLKBUF_X1 U8726 ( .A(n17943), .Z(n17928) );
  CLKBUF_X1 U8727 ( .A(n17943), .Z(n17929) );
  CLKBUF_X1 U8728 ( .A(n17943), .Z(n17930) );
  CLKBUF_X1 U8729 ( .A(n17943), .Z(n17931) );
  CLKBUF_X1 U8730 ( .A(n17943), .Z(n17932) );
  CLKBUF_X1 U8731 ( .A(n17943), .Z(n17933) );
  CLKBUF_X1 U8732 ( .A(n17931), .Z(n17934) );
  CLKBUF_X1 U8733 ( .A(n17933), .Z(n17935) );
  CLKBUF_X1 U8734 ( .A(n17926), .Z(n17936) );
  CLKBUF_X1 U8735 ( .A(n17943), .Z(n17937) );
  CLKBUF_X1 U8736 ( .A(n17941), .Z(n17938) );
  CLKBUF_X1 U8737 ( .A(n17943), .Z(n17939) );
  CLKBUF_X1 U8738 ( .A(n17932), .Z(n17940) );
  CLKBUF_X1 U8739 ( .A(n17943), .Z(n17941) );
  CLKBUF_X1 U8740 ( .A(n17943), .Z(n17942) );
  INV_X1 U8741 ( .A(n4076), .ZN(n17943) );
  INV_X1 U8742 ( .A(n17963), .ZN(n17946) );
  CLKBUF_X1 U8743 ( .A(n17964), .Z(n17947) );
  CLKBUF_X1 U8744 ( .A(n17964), .Z(n17948) );
  CLKBUF_X1 U8745 ( .A(n17964), .Z(n17949) );
  CLKBUF_X1 U8746 ( .A(n17964), .Z(n17950) );
  CLKBUF_X1 U8747 ( .A(n17964), .Z(n17951) );
  CLKBUF_X1 U8748 ( .A(n17964), .Z(n17952) );
  CLKBUF_X1 U8749 ( .A(n17951), .Z(n17953) );
  CLKBUF_X1 U8750 ( .A(n17947), .Z(n17954) );
  CLKBUF_X1 U8751 ( .A(n17952), .Z(n17955) );
  CLKBUF_X1 U8752 ( .A(n17950), .Z(n17956) );
  CLKBUF_X1 U8753 ( .A(n17962), .Z(n17957) );
  CLKBUF_X1 U8754 ( .A(n17964), .Z(n17958) );
  CLKBUF_X1 U8755 ( .A(n17964), .Z(n17959) );
  CLKBUF_X1 U8756 ( .A(n17964), .Z(n17960) );
  CLKBUF_X1 U8757 ( .A(n17949), .Z(n17961) );
  CLKBUF_X1 U8758 ( .A(n17964), .Z(n17962) );
  CLKBUF_X1 U8759 ( .A(n17964), .Z(n17963) );
  INV_X1 U8760 ( .A(n4073), .ZN(n17964) );
  INV_X1 U8761 ( .A(n17984), .ZN(n17967) );
  CLKBUF_X1 U8762 ( .A(n17985), .Z(n17968) );
  CLKBUF_X1 U8763 ( .A(n17972), .Z(n17969) );
  CLKBUF_X1 U8764 ( .A(n17985), .Z(n17970) );
  CLKBUF_X1 U8765 ( .A(n17985), .Z(n17971) );
  CLKBUF_X1 U8766 ( .A(n17985), .Z(n17972) );
  CLKBUF_X1 U8767 ( .A(n17985), .Z(n17973) );
  CLKBUF_X1 U8768 ( .A(n17985), .Z(n17974) );
  CLKBUF_X1 U8769 ( .A(n17985), .Z(n17975) );
  CLKBUF_X1 U8770 ( .A(n17973), .Z(n17976) );
  CLKBUF_X1 U8771 ( .A(n17975), .Z(n17977) );
  CLKBUF_X1 U8772 ( .A(n17968), .Z(n17978) );
  CLKBUF_X1 U8773 ( .A(n17983), .Z(n17979) );
  CLKBUF_X1 U8774 ( .A(n17985), .Z(n17980) );
  CLKBUF_X1 U8775 ( .A(n17985), .Z(n17981) );
  CLKBUF_X1 U8776 ( .A(n17974), .Z(n17982) );
  CLKBUF_X1 U8777 ( .A(n17985), .Z(n17983) );
  CLKBUF_X1 U8778 ( .A(n17985), .Z(n17984) );
  INV_X1 U8779 ( .A(n4070), .ZN(n17985) );
  INV_X1 U8780 ( .A(n18051), .ZN(n18033) );
endmodule


module reg_N5_1 ( clk, rst, d_in, d_out );
  input [4:0] d_in;
  output [4:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6;

  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[2]), .A2(rst), .ZN(N4) );
  AND2_X1 U4 ( .A1(d_in[3]), .A2(rst), .ZN(N5) );
  AND2_X1 U5 ( .A1(d_in[1]), .A2(rst), .ZN(N3) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U7 ( .A1(rst), .A2(d_in[4]), .ZN(N6) );
endmodule


module reg_N5_2 ( clk, rst, d_in, d_out );
  input [4:0] d_in;
  output [4:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6;

  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[2]), .A2(rst), .ZN(N4) );
  AND2_X1 U4 ( .A1(d_in[3]), .A2(rst), .ZN(N5) );
  AND2_X1 U5 ( .A1(d_in[1]), .A2(rst), .ZN(N3) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U7 ( .A1(rst), .A2(d_in[4]), .ZN(N6) );
endmodule


module reg_N5_0 ( clk, rst, d_in, d_out );
  input [4:0] d_in;
  output [4:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6;

  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[1]), .A2(rst), .ZN(N3) );
  AND2_X1 U4 ( .A1(d_in[2]), .A2(rst), .ZN(N4) );
  AND2_X1 U5 ( .A1(rst), .A2(d_in[4]), .ZN(N6) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[3]), .A2(rst), .ZN(N5) );
endmodule


module reg_N6_1 ( clk, rst, d_in, d_out );
  input [5:0] d_in;
  output [5:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7;

  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(rst), .A2(d_in[5]), .ZN(N7) );
  AND2_X1 U4 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U5 ( .A1(d_in[1]), .A2(rst), .ZN(N3) );
  AND2_X1 U6 ( .A1(d_in[2]), .A2(rst), .ZN(N4) );
  AND2_X1 U7 ( .A1(d_in[3]), .A2(rst), .ZN(N5) );
  AND2_X1 U8 ( .A1(d_in[4]), .A2(rst), .ZN(N6) );
endmodule


module reg_N6_0 ( clk, rst, d_in, d_out );
  input [5:0] d_in;
  output [5:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7;

  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  AND2_X1 U3 ( .A1(d_in[3]), .A2(rst), .ZN(N5) );
  AND2_X1 U4 ( .A1(d_in[4]), .A2(rst), .ZN(N6) );
  AND2_X1 U5 ( .A1(rst), .A2(d_in[5]), .ZN(N7) );
  AND2_X1 U6 ( .A1(d_in[2]), .A2(rst), .ZN(N4) );
  AND2_X1 U7 ( .A1(d_in[0]), .A2(rst), .ZN(N2) );
  AND2_X1 U8 ( .A1(d_in[1]), .A2(rst), .ZN(N3) );
endmodule


module reg_N32_0 ( clk, rst, d_in, d_out );
  input [31:0] d_in;
  output [31:0] d_out;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n68, n69, n70;

  DFF_X1 \d_out_reg[31]  ( .D(N33), .CK(clk), .Q(d_out[31]) );
  DFF_X1 \d_out_reg[30]  ( .D(N32), .CK(clk), .Q(d_out[30]) );
  DFF_X1 \d_out_reg[29]  ( .D(N31), .CK(clk), .Q(d_out[29]) );
  DFF_X1 \d_out_reg[28]  ( .D(N30), .CK(clk), .Q(d_out[28]) );
  DFF_X1 \d_out_reg[27]  ( .D(N29), .CK(clk), .Q(d_out[27]) );
  DFF_X1 \d_out_reg[26]  ( .D(N28), .CK(clk), .Q(d_out[26]) );
  DFF_X1 \d_out_reg[25]  ( .D(N27), .CK(clk), .Q(d_out[25]) );
  DFF_X1 \d_out_reg[24]  ( .D(N26), .CK(clk), .Q(d_out[24]) );
  DFF_X1 \d_out_reg[23]  ( .D(N25), .CK(clk), .Q(d_out[23]) );
  DFF_X1 \d_out_reg[22]  ( .D(N24), .CK(clk), .Q(d_out[22]) );
  DFF_X1 \d_out_reg[21]  ( .D(N23), .CK(clk), .Q(d_out[21]) );
  DFF_X1 \d_out_reg[20]  ( .D(N22), .CK(clk), .Q(d_out[20]) );
  DFF_X1 \d_out_reg[19]  ( .D(N21), .CK(clk), .Q(d_out[19]) );
  DFF_X1 \d_out_reg[18]  ( .D(N20), .CK(clk), .Q(d_out[18]) );
  DFF_X1 \d_out_reg[17]  ( .D(N19), .CK(clk), .Q(d_out[17]) );
  DFF_X1 \d_out_reg[16]  ( .D(N18), .CK(clk), .Q(d_out[16]) );
  DFF_X1 \d_out_reg[15]  ( .D(N17), .CK(clk), .Q(d_out[15]) );
  DFF_X1 \d_out_reg[14]  ( .D(N16), .CK(clk), .Q(d_out[14]) );
  DFF_X1 \d_out_reg[13]  ( .D(N15), .CK(clk), .Q(d_out[13]) );
  DFF_X1 \d_out_reg[12]  ( .D(N14), .CK(clk), .Q(d_out[12]) );
  DFF_X1 \d_out_reg[11]  ( .D(N13), .CK(clk), .Q(d_out[11]) );
  DFF_X1 \d_out_reg[10]  ( .D(N12), .CK(clk), .Q(d_out[10]) );
  DFF_X1 \d_out_reg[9]  ( .D(N11), .CK(clk), .Q(d_out[9]) );
  DFF_X1 \d_out_reg[8]  ( .D(N10), .CK(clk), .Q(d_out[8]) );
  DFF_X1 \d_out_reg[7]  ( .D(N9), .CK(clk), .Q(d_out[7]) );
  DFF_X1 \d_out_reg[6]  ( .D(N8), .CK(clk), .Q(d_out[6]) );
  DFF_X1 \d_out_reg[5]  ( .D(N7), .CK(clk), .Q(d_out[5]) );
  DFF_X1 \d_out_reg[4]  ( .D(N6), .CK(clk), .Q(d_out[4]) );
  DFF_X1 \d_out_reg[3]  ( .D(N5), .CK(clk), .Q(d_out[3]) );
  DFF_X1 \d_out_reg[2]  ( .D(N4), .CK(clk), .Q(d_out[2]) );
  DFF_X1 \d_out_reg[1]  ( .D(N3), .CK(clk), .Q(d_out[1]) );
  DFF_X1 \d_out_reg[0]  ( .D(N2), .CK(clk), .Q(d_out[0]) );
  BUF_X1 U3 ( .A(rst), .Z(n68) );
  BUF_X1 U4 ( .A(rst), .Z(n69) );
  BUF_X1 U5 ( .A(rst), .Z(n70) );
  AND2_X1 U6 ( .A1(d_in[0]), .A2(n68), .ZN(N2) );
  AND2_X1 U7 ( .A1(d_in[1]), .A2(n69), .ZN(N3) );
  AND2_X1 U8 ( .A1(d_in[8]), .A2(n68), .ZN(N10) );
  AND2_X1 U9 ( .A1(d_in[9]), .A2(n68), .ZN(N11) );
  AND2_X1 U10 ( .A1(d_in[10]), .A2(n68), .ZN(N12) );
  AND2_X1 U11 ( .A1(d_in[11]), .A2(n68), .ZN(N13) );
  AND2_X1 U12 ( .A1(d_in[12]), .A2(n68), .ZN(N14) );
  AND2_X1 U13 ( .A1(d_in[13]), .A2(n68), .ZN(N15) );
  AND2_X1 U14 ( .A1(d_in[14]), .A2(n68), .ZN(N16) );
  AND2_X1 U15 ( .A1(d_in[15]), .A2(n68), .ZN(N17) );
  AND2_X1 U16 ( .A1(d_in[16]), .A2(n68), .ZN(N18) );
  AND2_X1 U17 ( .A1(d_in[17]), .A2(n68), .ZN(N19) );
  AND2_X1 U18 ( .A1(d_in[18]), .A2(n68), .ZN(N20) );
  AND2_X1 U19 ( .A1(d_in[19]), .A2(n69), .ZN(N21) );
  AND2_X1 U20 ( .A1(d_in[20]), .A2(n69), .ZN(N22) );
  AND2_X1 U21 ( .A1(d_in[21]), .A2(n69), .ZN(N23) );
  AND2_X1 U22 ( .A1(d_in[22]), .A2(n69), .ZN(N24) );
  AND2_X1 U23 ( .A1(d_in[23]), .A2(n69), .ZN(N25) );
  AND2_X1 U24 ( .A1(d_in[24]), .A2(n69), .ZN(N26) );
  AND2_X1 U25 ( .A1(d_in[25]), .A2(n69), .ZN(N27) );
  AND2_X1 U26 ( .A1(d_in[26]), .A2(n69), .ZN(N28) );
  AND2_X1 U27 ( .A1(d_in[27]), .A2(n69), .ZN(N29) );
  AND2_X1 U28 ( .A1(d_in[28]), .A2(n69), .ZN(N30) );
  AND2_X1 U29 ( .A1(d_in[29]), .A2(n69), .ZN(N31) );
  AND2_X1 U30 ( .A1(n70), .A2(d_in[7]), .ZN(N9) );
  AND2_X1 U31 ( .A1(d_in[2]), .A2(n70), .ZN(N4) );
  AND2_X1 U32 ( .A1(d_in[3]), .A2(n70), .ZN(N5) );
  AND2_X1 U33 ( .A1(d_in[4]), .A2(n70), .ZN(N6) );
  AND2_X1 U34 ( .A1(d_in[5]), .A2(n70), .ZN(N7) );
  AND2_X1 U35 ( .A1(d_in[6]), .A2(n70), .ZN(N8) );
  AND2_X1 U36 ( .A1(d_in[30]), .A2(n70), .ZN(N32) );
  AND2_X1 U37 ( .A1(d_in[31]), .A2(n70), .ZN(N33) );
endmodule


module cla_adder_N32 ( A, B, Ci, Cout, Sum );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Ci;
  output Cout;

  wire   [8:0] Carry;

  carry_generator_N32_Nblocks8 CG ( .A(A), .B(B), .Ci(Ci), .Cout(Carry) );
  sum_generator_Nbits32_Nblocks8 SG ( .A(A), .B(B), .Carry(Carry), .S(Sum), 
        .Cout(Cout) );
endmodule


module alu ( A, B, .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), Y1, 
        cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y1;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  output cout;
  wire   add_sub, sign, N25, N26, N27, N28, N29, N31, N32, N33, N34, N35, N36,
         gt, get, lt, let, eq, neq, n23, n24, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98;
  wire   [31:0] A_add;
  wire   [31:0] B_add;
  wire   [15:0] A_mul;
  wire   [15:0] B_mul;
  wire   [3:0] sel_log;
  wire   [31:0] A_log;
  wire   [31:0] B_log;
  wire   [1:0] sel_shift;
  wire   [31:0] A_sht;
  wire   [31:0] B_sht;
  wire   [15:0] B_lhi;
  wire   [31:0] out_add;
  wire   [31:0] out_mul;
  wire   [31:0] out_log;
  wire   [31:0] out_shift;
  tri   [31:0] Y1;

  adder_sub_N32 adder_subtr ( .A(A_add), .B(B_add), .Ci(add_sub), .Cout(cout), 
        .Sum(out_add) );
  booth_mul_N16 mul ( .A({A_mul[15:1], n23}), .B(B_mul), .Y(out_mul) );
  logical logic ( .A(A_log), .B(B_log), .sel({1'b0, sel_log[2:0]}), .Y(out_log) );
  shifter shift ( .A(A_sht), .B(B_sht), .sel(sel_shift), .C(out_shift) );
  comparator compar ( .C(cout), .Sum(out_add), .sign(sign), .gt(gt), .get(get), 
        .lt(lt), .let(let), .eq(eq), .neq(neq) );
  mux_alu muxy1 ( .addsub(out_add), .mul(out_mul), .log(out_log), .shift(
        out_shift), .lhi({B_lhi, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .gt(gt), .get(
        get), .lt(lt), .let(let), .eq(eq), .neq(neq), .sel({\OP[4] , \OP[3] , 
        \OP[2] , \OP[1] , \OP[0] }), .out_mux(Y1) );
  DLH_X1 \B_lhi_reg[15]  ( .G(N36), .D(B[15]), .Q(B_lhi[15]) );
  DLH_X1 \B_lhi_reg[14]  ( .G(N36), .D(B[14]), .Q(B_lhi[14]) );
  DLH_X1 \B_lhi_reg[13]  ( .G(N36), .D(B[13]), .Q(B_lhi[13]) );
  DLH_X1 \B_lhi_reg[12]  ( .G(N36), .D(B[12]), .Q(B_lhi[12]) );
  DLH_X1 \B_lhi_reg[11]  ( .G(N36), .D(B[11]), .Q(B_lhi[11]) );
  DLH_X1 \B_lhi_reg[10]  ( .G(N36), .D(B[10]), .Q(B_lhi[10]) );
  DLH_X1 \B_lhi_reg[9]  ( .G(N36), .D(B[9]), .Q(B_lhi[9]) );
  DLH_X1 \B_lhi_reg[8]  ( .G(N36), .D(B[8]), .Q(B_lhi[8]) );
  DLH_X1 \B_lhi_reg[7]  ( .G(N36), .D(B[7]), .Q(B_lhi[7]) );
  DLH_X1 \B_lhi_reg[6]  ( .G(N36), .D(B[6]), .Q(B_lhi[6]) );
  DLH_X1 \B_lhi_reg[5]  ( .G(N36), .D(B[5]), .Q(B_lhi[5]) );
  DLH_X1 \B_lhi_reg[4]  ( .G(N36), .D(B[4]), .Q(B_lhi[4]) );
  DLH_X1 \B_lhi_reg[3]  ( .G(N36), .D(B[3]), .Q(B_lhi[3]) );
  DLH_X1 \B_lhi_reg[2]  ( .G(N36), .D(B[2]), .Q(B_lhi[2]) );
  DLH_X1 \B_lhi_reg[1]  ( .G(N36), .D(B[1]), .Q(B_lhi[1]) );
  DLH_X1 \B_lhi_reg[0]  ( .G(N36), .D(B[0]), .Q(B_lhi[0]) );
  DLH_X1 \A_add_reg[31]  ( .G(n98), .D(A[31]), .Q(A_add[31]) );
  DLH_X1 \A_add_reg[30]  ( .G(n98), .D(A[30]), .Q(A_add[30]) );
  DLH_X1 \A_add_reg[29]  ( .G(n98), .D(A[29]), .Q(A_add[29]) );
  DLH_X1 \A_add_reg[28]  ( .G(n98), .D(A[28]), .Q(A_add[28]) );
  DLH_X1 \A_add_reg[27]  ( .G(n98), .D(A[27]), .Q(A_add[27]) );
  DLH_X1 \A_add_reg[26]  ( .G(n98), .D(A[26]), .Q(A_add[26]) );
  DLH_X1 \A_add_reg[25]  ( .G(n98), .D(A[25]), .Q(A_add[25]) );
  DLH_X1 \A_add_reg[24]  ( .G(n98), .D(A[24]), .Q(A_add[24]) );
  DLH_X1 \A_add_reg[23]  ( .G(n98), .D(A[23]), .Q(A_add[23]) );
  DLH_X1 \A_add_reg[22]  ( .G(n98), .D(A[22]), .Q(A_add[22]) );
  DLH_X1 \A_add_reg[21]  ( .G(n97), .D(A[21]), .Q(A_add[21]) );
  DLH_X1 \A_add_reg[20]  ( .G(n97), .D(A[20]), .Q(A_add[20]) );
  DLH_X1 \A_add_reg[19]  ( .G(n97), .D(A[19]), .Q(A_add[19]) );
  DLH_X1 \A_add_reg[18]  ( .G(n97), .D(A[18]), .Q(A_add[18]) );
  DLH_X1 \A_add_reg[17]  ( .G(n97), .D(A[17]), .Q(A_add[17]) );
  DLH_X1 \A_add_reg[16]  ( .G(n97), .D(A[16]), .Q(A_add[16]) );
  DLH_X1 \A_add_reg[15]  ( .G(n97), .D(A[15]), .Q(A_add[15]) );
  DLH_X1 \A_add_reg[14]  ( .G(n97), .D(A[14]), .Q(A_add[14]) );
  DLH_X1 \A_add_reg[13]  ( .G(n97), .D(A[13]), .Q(A_add[13]) );
  DLH_X1 \A_add_reg[12]  ( .G(n97), .D(A[12]), .Q(A_add[12]) );
  DLH_X1 \A_add_reg[11]  ( .G(n97), .D(A[11]), .Q(A_add[11]) );
  DLH_X1 \A_add_reg[10]  ( .G(n96), .D(A[10]), .Q(A_add[10]) );
  DLH_X1 \A_add_reg[9]  ( .G(n96), .D(A[9]), .Q(A_add[9]) );
  DLH_X1 \A_add_reg[8]  ( .G(n96), .D(A[8]), .Q(A_add[8]) );
  DLH_X1 \A_add_reg[7]  ( .G(n96), .D(A[7]), .Q(A_add[7]) );
  DLH_X1 \A_add_reg[6]  ( .G(n96), .D(A[6]), .Q(A_add[6]) );
  DLH_X1 \A_add_reg[5]  ( .G(n96), .D(A[5]), .Q(A_add[5]) );
  DLH_X1 \A_add_reg[4]  ( .G(n96), .D(A[4]), .Q(A_add[4]) );
  DLH_X1 \A_add_reg[3]  ( .G(n96), .D(A[3]), .Q(A_add[3]) );
  DLH_X1 \A_add_reg[2]  ( .G(n96), .D(A[2]), .Q(A_add[2]) );
  DLH_X1 \A_add_reg[1]  ( .G(n96), .D(A[1]), .Q(A_add[1]) );
  DLH_X1 \A_add_reg[0]  ( .G(n96), .D(A[0]), .Q(A_add[0]) );
  DLH_X1 \B_add_reg[31]  ( .G(n95), .D(B[31]), .Q(B_add[31]) );
  DLH_X1 \B_add_reg[30]  ( .G(n95), .D(B[30]), .Q(B_add[30]) );
  DLH_X1 \B_add_reg[29]  ( .G(n95), .D(B[29]), .Q(B_add[29]) );
  DLH_X1 \B_add_reg[28]  ( .G(n95), .D(B[28]), .Q(B_add[28]) );
  DLH_X1 \B_add_reg[27]  ( .G(n95), .D(B[27]), .Q(B_add[27]) );
  DLH_X1 \B_add_reg[26]  ( .G(n95), .D(B[26]), .Q(B_add[26]) );
  DLH_X1 \B_add_reg[25]  ( .G(n95), .D(B[25]), .Q(B_add[25]) );
  DLH_X1 \B_add_reg[24]  ( .G(n95), .D(B[24]), .Q(B_add[24]) );
  DLH_X1 \B_add_reg[23]  ( .G(n95), .D(B[23]), .Q(B_add[23]) );
  DLH_X1 \B_add_reg[22]  ( .G(n95), .D(B[22]), .Q(B_add[22]) );
  DLH_X1 \B_add_reg[21]  ( .G(n95), .D(B[21]), .Q(B_add[21]) );
  DLH_X1 \B_add_reg[20]  ( .G(n94), .D(B[20]), .Q(B_add[20]) );
  DLH_X1 \B_add_reg[19]  ( .G(n94), .D(B[19]), .Q(B_add[19]) );
  DLH_X1 \B_add_reg[18]  ( .G(n94), .D(B[18]), .Q(B_add[18]) );
  DLH_X1 \B_add_reg[17]  ( .G(n94), .D(B[17]), .Q(B_add[17]) );
  DLH_X1 \B_add_reg[16]  ( .G(n94), .D(B[16]), .Q(B_add[16]) );
  DLH_X1 \B_add_reg[15]  ( .G(n94), .D(B[15]), .Q(B_add[15]) );
  DLH_X1 \B_add_reg[14]  ( .G(n94), .D(B[14]), .Q(B_add[14]) );
  DLH_X1 \B_add_reg[13]  ( .G(n94), .D(B[13]), .Q(B_add[13]) );
  DLH_X1 \B_add_reg[12]  ( .G(n94), .D(B[12]), .Q(B_add[12]) );
  DLH_X1 \B_add_reg[11]  ( .G(n94), .D(B[11]), .Q(B_add[11]) );
  DLH_X1 \B_add_reg[10]  ( .G(n94), .D(B[10]), .Q(B_add[10]) );
  DLH_X1 \B_add_reg[9]  ( .G(n93), .D(B[9]), .Q(B_add[9]) );
  DLH_X1 \B_add_reg[8]  ( .G(n93), .D(B[8]), .Q(B_add[8]) );
  DLH_X1 \B_add_reg[7]  ( .G(n93), .D(B[7]), .Q(B_add[7]) );
  DLH_X1 \B_add_reg[6]  ( .G(n93), .D(B[6]), .Q(B_add[6]) );
  DLH_X1 \B_add_reg[5]  ( .G(n93), .D(B[5]), .Q(B_add[5]) );
  DLH_X1 \B_add_reg[4]  ( .G(n93), .D(B[4]), .Q(B_add[4]) );
  DLH_X1 \B_add_reg[3]  ( .G(n93), .D(B[3]), .Q(B_add[3]) );
  DLH_X1 \B_add_reg[2]  ( .G(n93), .D(B[2]), .Q(B_add[2]) );
  DLH_X1 \B_add_reg[1]  ( .G(n93), .D(B[1]), .Q(B_add[1]) );
  DLH_X1 \B_add_reg[0]  ( .G(n93), .D(B[0]), .Q(B_add[0]) );
  DLH_X1 \A_mul_reg[15]  ( .G(n92), .D(A[15]), .Q(A_mul[15]) );
  DLH_X1 \A_mul_reg[0]  ( .G(n92), .D(A[0]), .Q(n23) );
  DLH_X1 \B_mul_reg[15]  ( .G(n92), .D(B[15]), .Q(B_mul[15]) );
  DLH_X1 \B_mul_reg[14]  ( .G(n92), .D(B[14]), .Q(B_mul[14]) );
  DLH_X1 \B_mul_reg[13]  ( .G(n92), .D(B[13]), .Q(B_mul[13]) );
  DLH_X1 \B_mul_reg[12]  ( .G(n92), .D(B[12]), .Q(B_mul[12]) );
  DLH_X1 \B_mul_reg[11]  ( .G(n92), .D(B[11]), .Q(B_mul[11]) );
  DLH_X1 \B_mul_reg[10]  ( .G(n92), .D(B[10]), .Q(B_mul[10]) );
  DLH_X1 \B_mul_reg[9]  ( .G(n92), .D(B[9]), .Q(B_mul[9]) );
  DLH_X1 \B_mul_reg[8]  ( .G(n92), .D(B[8]), .Q(B_mul[8]) );
  DLH_X1 \B_mul_reg[7]  ( .G(n91), .D(B[7]), .Q(B_mul[7]) );
  DLH_X1 \B_mul_reg[6]  ( .G(n91), .D(B[6]), .Q(B_mul[6]) );
  DLH_X1 \B_mul_reg[5]  ( .G(n91), .D(B[5]), .Q(B_mul[5]) );
  DLH_X1 \B_mul_reg[4]  ( .G(n91), .D(B[4]), .Q(B_mul[4]) );
  DLH_X1 \B_mul_reg[3]  ( .G(n91), .D(B[3]), .Q(B_mul[3]) );
  DLH_X1 \B_mul_reg[2]  ( .G(n91), .D(B[2]), .Q(B_mul[2]) );
  DLH_X1 \B_mul_reg[1]  ( .G(n91), .D(B[1]), .Q(B_mul[1]) );
  DLH_X1 \B_mul_reg[0]  ( .G(n91), .D(B[0]), .Q(B_mul[0]) );
  DLH_X1 \sel_log_reg[2]  ( .G(n78), .D(N29), .Q(sel_log[2]) );
  DLH_X1 \sel_log_reg[1]  ( .G(n78), .D(N29), .Q(sel_log[1]) );
  DLH_X1 \sel_log_reg[0]  ( .G(n78), .D(N28), .Q(sel_log[0]) );
  DLH_X1 \A_log_reg[31]  ( .G(n78), .D(A[31]), .Q(A_log[31]) );
  DLH_X1 \A_log_reg[30]  ( .G(n78), .D(A[30]), .Q(A_log[30]) );
  DLH_X1 \A_log_reg[29]  ( .G(n78), .D(A[29]), .Q(A_log[29]) );
  DLH_X1 \A_log_reg[28]  ( .G(n78), .D(A[28]), .Q(A_log[28]) );
  DLH_X1 \A_log_reg[27]  ( .G(n78), .D(A[27]), .Q(A_log[27]) );
  DLH_X1 \A_log_reg[26]  ( .G(n78), .D(A[26]), .Q(A_log[26]) );
  DLH_X1 \A_log_reg[25]  ( .G(n78), .D(A[25]), .Q(A_log[25]) );
  DLH_X1 \A_log_reg[24]  ( .G(n78), .D(A[24]), .Q(A_log[24]) );
  DLH_X1 \A_log_reg[23]  ( .G(n79), .D(A[23]), .Q(A_log[23]) );
  DLH_X1 \A_log_reg[22]  ( .G(n79), .D(A[22]), .Q(A_log[22]) );
  DLH_X1 \A_log_reg[21]  ( .G(n79), .D(A[21]), .Q(A_log[21]) );
  DLH_X1 \A_log_reg[20]  ( .G(n79), .D(A[20]), .Q(A_log[20]) );
  DLH_X1 \A_log_reg[19]  ( .G(n79), .D(A[19]), .Q(A_log[19]) );
  DLH_X1 \A_log_reg[18]  ( .G(n79), .D(A[18]), .Q(A_log[18]) );
  DLH_X1 \A_log_reg[17]  ( .G(n79), .D(A[17]), .Q(A_log[17]) );
  DLH_X1 \A_log_reg[16]  ( .G(n79), .D(A[16]), .Q(A_log[16]) );
  DLH_X1 \A_log_reg[15]  ( .G(n79), .D(A[15]), .Q(A_log[15]) );
  DLH_X1 \A_log_reg[14]  ( .G(n79), .D(A[14]), .Q(A_log[14]) );
  DLH_X1 \A_log_reg[13]  ( .G(n79), .D(A[13]), .Q(A_log[13]) );
  DLH_X1 \A_log_reg[12]  ( .G(n80), .D(A[12]), .Q(A_log[12]) );
  DLH_X1 \A_log_reg[11]  ( .G(n80), .D(A[11]), .Q(A_log[11]) );
  DLH_X1 \A_log_reg[10]  ( .G(n80), .D(A[10]), .Q(A_log[10]) );
  DLH_X1 \A_log_reg[9]  ( .G(n80), .D(A[9]), .Q(A_log[9]) );
  DLH_X1 \A_log_reg[8]  ( .G(n80), .D(A[8]), .Q(A_log[8]) );
  DLH_X1 \A_log_reg[7]  ( .G(n80), .D(A[7]), .Q(A_log[7]) );
  DLH_X1 \A_log_reg[6]  ( .G(n80), .D(A[6]), .Q(A_log[6]) );
  DLH_X1 \A_log_reg[5]  ( .G(n80), .D(A[5]), .Q(A_log[5]) );
  DLH_X1 \A_log_reg[4]  ( .G(n80), .D(A[4]), .Q(A_log[4]) );
  DLH_X1 \A_log_reg[3]  ( .G(n80), .D(A[3]), .Q(A_log[3]) );
  DLH_X1 \A_log_reg[2]  ( .G(n80), .D(A[2]), .Q(A_log[2]) );
  DLH_X1 \A_log_reg[1]  ( .G(n81), .D(A[1]), .Q(A_log[1]) );
  DLH_X1 \A_log_reg[0]  ( .G(n81), .D(A[0]), .Q(A_log[0]) );
  DLH_X1 \B_log_reg[31]  ( .G(n81), .D(B[31]), .Q(B_log[31]) );
  DLH_X1 \B_log_reg[30]  ( .G(n81), .D(B[30]), .Q(B_log[30]) );
  DLH_X1 \B_log_reg[29]  ( .G(n81), .D(B[29]), .Q(B_log[29]) );
  DLH_X1 \B_log_reg[28]  ( .G(n81), .D(B[28]), .Q(B_log[28]) );
  DLH_X1 \B_log_reg[27]  ( .G(n81), .D(B[27]), .Q(B_log[27]) );
  DLH_X1 \B_log_reg[26]  ( .G(n81), .D(B[26]), .Q(B_log[26]) );
  DLH_X1 \B_log_reg[25]  ( .G(n81), .D(B[25]), .Q(B_log[25]) );
  DLH_X1 \B_log_reg[24]  ( .G(n81), .D(B[24]), .Q(B_log[24]) );
  DLH_X1 \B_log_reg[23]  ( .G(n81), .D(B[23]), .Q(B_log[23]) );
  DLH_X1 \B_log_reg[22]  ( .G(n82), .D(B[22]), .Q(B_log[22]) );
  DLH_X1 \B_log_reg[21]  ( .G(n82), .D(B[21]), .Q(B_log[21]) );
  DLH_X1 \B_log_reg[20]  ( .G(n82), .D(B[20]), .Q(B_log[20]) );
  DLH_X1 \B_log_reg[19]  ( .G(n82), .D(B[19]), .Q(B_log[19]) );
  DLH_X1 \B_log_reg[18]  ( .G(n82), .D(B[18]), .Q(B_log[18]) );
  DLH_X1 \B_log_reg[17]  ( .G(n82), .D(B[17]), .Q(B_log[17]) );
  DLH_X1 \B_log_reg[16]  ( .G(n82), .D(B[16]), .Q(B_log[16]) );
  DLH_X1 \B_log_reg[15]  ( .G(n82), .D(B[15]), .Q(B_log[15]) );
  DLH_X1 \B_log_reg[14]  ( .G(n82), .D(B[14]), .Q(B_log[14]) );
  DLH_X1 \B_log_reg[13]  ( .G(n82), .D(B[13]), .Q(B_log[13]) );
  DLH_X1 \B_log_reg[12]  ( .G(n82), .D(B[12]), .Q(B_log[12]) );
  DLH_X1 \B_log_reg[11]  ( .G(n83), .D(B[11]), .Q(B_log[11]) );
  DLH_X1 \B_log_reg[10]  ( .G(n83), .D(B[10]), .Q(B_log[10]) );
  DLH_X1 \B_log_reg[9]  ( .G(n83), .D(B[9]), .Q(B_log[9]) );
  DLH_X1 \B_log_reg[8]  ( .G(n83), .D(B[8]), .Q(B_log[8]) );
  DLH_X1 \B_log_reg[7]  ( .G(n83), .D(B[7]), .Q(B_log[7]) );
  DLH_X1 \B_log_reg[6]  ( .G(n83), .D(B[6]), .Q(B_log[6]) );
  DLH_X1 \B_log_reg[5]  ( .G(n83), .D(B[5]), .Q(B_log[5]) );
  DLH_X1 \B_log_reg[4]  ( .G(n83), .D(B[4]), .Q(B_log[4]) );
  DLH_X1 \B_log_reg[3]  ( .G(n83), .D(B[3]), .Q(B_log[3]) );
  DLH_X1 \B_log_reg[2]  ( .G(n83), .D(B[2]), .Q(B_log[2]) );
  DLH_X1 \B_log_reg[1]  ( .G(n83), .D(B[1]), .Q(B_log[1]) );
  DLH_X1 \B_log_reg[0]  ( .G(n24), .D(B[0]), .Q(B_log[0]) );
  DLH_X1 \sel_shift_reg[1]  ( .G(n89), .D(N32), .Q(sel_shift[1]) );
  DLH_X1 \sel_shift_reg[0]  ( .G(n89), .D(N31), .Q(sel_shift[0]) );
  DLH_X1 \A_sht_reg[31]  ( .G(n89), .D(A[31]), .Q(A_sht[31]) );
  DLH_X1 \A_sht_reg[30]  ( .G(n89), .D(A[30]), .Q(A_sht[30]) );
  DLH_X1 \A_sht_reg[29]  ( .G(n89), .D(A[29]), .Q(A_sht[29]) );
  DLH_X1 \A_sht_reg[28]  ( .G(n89), .D(A[28]), .Q(A_sht[28]) );
  DLH_X1 \A_sht_reg[27]  ( .G(n89), .D(A[27]), .Q(A_sht[27]) );
  DLH_X1 \A_sht_reg[26]  ( .G(n89), .D(A[26]), .Q(A_sht[26]) );
  DLH_X1 \A_sht_reg[25]  ( .G(n89), .D(A[25]), .Q(A_sht[25]) );
  DLH_X1 \A_sht_reg[24]  ( .G(n89), .D(A[24]), .Q(A_sht[24]) );
  DLH_X1 \A_sht_reg[23]  ( .G(n89), .D(A[23]), .Q(A_sht[23]) );
  DLH_X1 \A_sht_reg[22]  ( .G(n88), .D(A[22]), .Q(A_sht[22]) );
  DLH_X1 \A_sht_reg[21]  ( .G(n88), .D(A[21]), .Q(A_sht[21]) );
  DLH_X1 \A_sht_reg[20]  ( .G(n88), .D(A[20]), .Q(A_sht[20]) );
  DLH_X1 \A_sht_reg[19]  ( .G(n88), .D(A[19]), .Q(A_sht[19]) );
  DLH_X1 \A_sht_reg[18]  ( .G(n88), .D(A[18]), .Q(A_sht[18]) );
  DLH_X1 \A_sht_reg[17]  ( .G(n88), .D(A[17]), .Q(A_sht[17]) );
  DLH_X1 \A_sht_reg[16]  ( .G(n88), .D(A[16]), .Q(A_sht[16]) );
  DLH_X1 \A_sht_reg[15]  ( .G(n88), .D(A[15]), .Q(A_sht[15]) );
  DLH_X1 \A_sht_reg[14]  ( .G(n88), .D(A[14]), .Q(A_sht[14]) );
  DLH_X1 \A_sht_reg[13]  ( .G(n88), .D(A[13]), .Q(A_sht[13]) );
  DLH_X1 \A_sht_reg[12]  ( .G(n88), .D(A[12]), .Q(A_sht[12]) );
  DLH_X1 \A_sht_reg[11]  ( .G(n87), .D(A[11]), .Q(A_sht[11]) );
  DLH_X1 \A_sht_reg[10]  ( .G(n87), .D(A[10]), .Q(A_sht[10]) );
  DLH_X1 \A_sht_reg[9]  ( .G(n87), .D(A[9]), .Q(A_sht[9]) );
  DLH_X1 \A_sht_reg[8]  ( .G(n87), .D(A[8]), .Q(A_sht[8]) );
  DLH_X1 \A_sht_reg[7]  ( .G(n87), .D(A[7]), .Q(A_sht[7]) );
  DLH_X1 \A_sht_reg[6]  ( .G(n87), .D(A[6]), .Q(A_sht[6]) );
  DLH_X1 \A_sht_reg[5]  ( .G(n87), .D(A[5]), .Q(A_sht[5]) );
  DLH_X1 \A_sht_reg[4]  ( .G(n87), .D(A[4]), .Q(A_sht[4]) );
  DLH_X1 \A_sht_reg[3]  ( .G(n87), .D(A[3]), .Q(A_sht[3]) );
  DLH_X1 \A_sht_reg[2]  ( .G(n87), .D(A[2]), .Q(A_sht[2]) );
  DLH_X1 \A_sht_reg[1]  ( .G(n87), .D(A[1]), .Q(A_sht[1]) );
  DLH_X1 \A_sht_reg[0]  ( .G(n86), .D(A[0]), .Q(A_sht[0]) );
  DLH_X1 \B_sht_reg[31]  ( .G(n86), .D(B[31]), .Q(B_sht[31]) );
  DLH_X1 \B_sht_reg[30]  ( .G(n86), .D(B[30]), .Q(B_sht[30]) );
  DLH_X1 \B_sht_reg[29]  ( .G(n86), .D(B[29]), .Q(B_sht[29]) );
  DLH_X1 \B_sht_reg[28]  ( .G(n86), .D(B[28]), .Q(B_sht[28]) );
  DLH_X1 \B_sht_reg[27]  ( .G(n86), .D(B[27]), .Q(B_sht[27]) );
  DLH_X1 \B_sht_reg[26]  ( .G(n86), .D(B[26]), .Q(B_sht[26]) );
  DLH_X1 \B_sht_reg[25]  ( .G(n86), .D(B[25]), .Q(B_sht[25]) );
  DLH_X1 \B_sht_reg[24]  ( .G(n86), .D(B[24]), .Q(B_sht[24]) );
  DLH_X1 \B_sht_reg[23]  ( .G(n86), .D(B[23]), .Q(B_sht[23]) );
  DLH_X1 \B_sht_reg[22]  ( .G(n86), .D(B[22]), .Q(B_sht[22]) );
  DLH_X1 \B_sht_reg[21]  ( .G(n85), .D(B[21]), .Q(B_sht[21]) );
  DLH_X1 \B_sht_reg[20]  ( .G(n85), .D(B[20]), .Q(B_sht[20]) );
  DLH_X1 \B_sht_reg[19]  ( .G(n85), .D(B[19]), .Q(B_sht[19]) );
  DLH_X1 \B_sht_reg[18]  ( .G(n85), .D(B[18]), .Q(B_sht[18]) );
  DLH_X1 \B_sht_reg[17]  ( .G(n85), .D(B[17]), .Q(B_sht[17]) );
  DLH_X1 \B_sht_reg[16]  ( .G(n85), .D(B[16]), .Q(B_sht[16]) );
  DLH_X1 \B_sht_reg[15]  ( .G(n85), .D(B[15]), .Q(B_sht[15]) );
  DLH_X1 \B_sht_reg[14]  ( .G(n85), .D(B[14]), .Q(B_sht[14]) );
  DLH_X1 \B_sht_reg[13]  ( .G(n85), .D(B[13]), .Q(B_sht[13]) );
  DLH_X1 \B_sht_reg[12]  ( .G(n85), .D(B[12]), .Q(B_sht[12]) );
  DLH_X1 \B_sht_reg[11]  ( .G(n85), .D(B[11]), .Q(B_sht[11]) );
  DLH_X1 \B_sht_reg[10]  ( .G(n84), .D(B[10]), .Q(B_sht[10]) );
  DLH_X1 \B_sht_reg[9]  ( .G(n84), .D(B[9]), .Q(B_sht[9]) );
  DLH_X1 \B_sht_reg[8]  ( .G(n84), .D(B[8]), .Q(B_sht[8]) );
  DLH_X1 \B_sht_reg[7]  ( .G(n84), .D(B[7]), .Q(B_sht[7]) );
  DLH_X1 \B_sht_reg[6]  ( .G(n84), .D(B[6]), .Q(B_sht[6]) );
  DLH_X1 \B_sht_reg[5]  ( .G(n84), .D(B[5]), .Q(B_sht[5]) );
  DLH_X1 \B_sht_reg[4]  ( .G(n84), .D(B[4]), .Q(B_sht[4]) );
  DLH_X1 \B_sht_reg[3]  ( .G(n84), .D(B[3]), .Q(B_sht[3]) );
  DLH_X1 \B_sht_reg[2]  ( .G(n84), .D(B[2]), .Q(B_sht[2]) );
  DLH_X1 \B_sht_reg[1]  ( .G(n84), .D(B[1]), .Q(B_sht[1]) );
  DLH_X1 \B_sht_reg[0]  ( .G(n84), .D(B[0]), .Q(B_sht[0]) );
  DLH_X1 sign_reg ( .G(N34), .D(N35), .Q(sign) );
  NAND3_X1 U63 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n58) );
  XOR2_X1 U64 ( .A(n66), .B(OP[2]), .Z(n63) );
  NAND3_X1 U65 ( .A1(n70), .A2(OP[2]), .A3(OP[0]), .ZN(n69) );
  NAND3_X1 U66 ( .A1(OP[2]), .A2(n59), .A3(n70), .ZN(n72) );
  NAND3_X1 U67 ( .A1(n66), .A2(n60), .A3(n61), .ZN(n57) );
  NAND3_X1 U68 ( .A1(n65), .A2(n60), .A3(OP[1]), .ZN(n73) );
  DLH_X1 \A_mul_reg[13]  ( .G(n91), .D(A[13]), .Q(A_mul[13]) );
  DLH_X1 \A_mul_reg[3]  ( .G(n91), .D(A[3]), .Q(A_mul[3]) );
  DLH_X1 \A_mul_reg[5]  ( .G(n91), .D(A[5]), .Q(A_mul[5]) );
  DLH_X1 \A_mul_reg[9]  ( .G(n90), .D(A[9]), .Q(A_mul[9]) );
  DLH_X1 \A_mul_reg[7]  ( .G(n90), .D(A[7]), .Q(A_mul[7]) );
  DLH_X1 \A_mul_reg[14]  ( .G(n90), .D(A[14]), .Q(A_mul[14]) );
  DLH_X1 \A_mul_reg[11]  ( .G(n90), .D(A[11]), .Q(A_mul[11]) );
  DLH_X1 \A_mul_reg[1]  ( .G(n90), .D(A[1]), .Q(A_mul[1]) );
  DLH_X1 \A_mul_reg[12]  ( .G(n90), .D(A[12]), .Q(A_mul[12]) );
  DLH_X1 \A_mul_reg[8]  ( .G(n90), .D(A[8]), .Q(A_mul[8]) );
  DLH_X1 \A_mul_reg[10]  ( .G(n90), .D(A[10]), .Q(A_mul[10]) );
  DLH_X1 \A_mul_reg[6]  ( .G(n90), .D(A[6]), .Q(A_mul[6]) );
  DLH_X1 \A_mul_reg[4]  ( .G(n90), .D(A[4]), .Q(A_mul[4]) );
  DLH_X1 add_sub_reg ( .G(n93), .D(N25), .Q(add_sub) );
  DLH_X1 \A_mul_reg[2]  ( .G(n90), .D(A[2]), .Q(A_mul[2]) );
  NOR4_X4 U69 ( .A1(OP[1]), .A2(OP[0]), .A3(n62), .A4(n60), .ZN(N36) );
  INV_X1 U70 ( .A(n57), .ZN(N28) );
  OAI21_X1 U71 ( .B1(n73), .B2(n76), .A(n67), .ZN(N25) );
  NAND2_X1 U72 ( .A1(n59), .A2(n71), .ZN(n76) );
  NAND2_X1 U73 ( .A1(n57), .A2(n58), .ZN(n24) );
  BUF_X1 U74 ( .A(N27), .Z(n90) );
  BUF_X1 U75 ( .A(N27), .Z(n91) );
  BUF_X1 U76 ( .A(N27), .Z(n92) );
  INV_X1 U77 ( .A(n73), .ZN(n70) );
  NOR2_X1 U78 ( .A1(n59), .A2(n68), .ZN(N32) );
  INV_X1 U79 ( .A(n67), .ZN(N34) );
  INV_X1 U80 ( .A(n62), .ZN(n61) );
  OAI221_X1 U81 ( .B1(n77), .B2(n65), .C1(OP[4]), .C2(OP[3]), .A(n62), .ZN(n67) );
  AOI21_X1 U82 ( .B1(n66), .B2(n71), .A(OP[4]), .ZN(n77) );
  NOR3_X1 U83 ( .A1(n59), .A2(OP[2]), .A3(n73), .ZN(N27) );
  NOR4_X1 U84 ( .A1(OP[4]), .A2(n63), .A3(n64), .A4(n65), .ZN(N35) );
  XNOR2_X1 U85 ( .A(B[31]), .B(A[31]), .ZN(n64) );
  NAND4_X1 U86 ( .A1(OP[3]), .A2(n66), .A3(n71), .A4(n60), .ZN(n68) );
  INV_X1 U87 ( .A(OP[0]), .ZN(n59) );
  INV_X1 U88 ( .A(OP[3]), .ZN(n65) );
  INV_X1 U89 ( .A(OP[1]), .ZN(n66) );
  INV_X1 U90 ( .A(OP[2]), .ZN(n71) );
  INV_X1 U91 ( .A(OP[4]), .ZN(n60) );
  NAND2_X1 U92 ( .A1(OP[2]), .A2(n65), .ZN(n62) );
  OAI21_X1 U93 ( .B1(n59), .B2(n57), .A(n72), .ZN(N29) );
  NAND2_X1 U94 ( .A1(n68), .A2(n69), .ZN(N33) );
  NAND2_X1 U95 ( .A1(n74), .A2(n75), .ZN(N26) );
  INV_X1 U96 ( .A(N25), .ZN(n75) );
  NAND4_X1 U97 ( .A1(OP[0]), .A2(n66), .A3(n71), .A4(n65), .ZN(n74) );
  NOR2_X1 U98 ( .A1(OP[0]), .A2(n68), .ZN(N31) );
  CLKBUF_X1 U99 ( .A(n24), .Z(n78) );
  CLKBUF_X1 U100 ( .A(n24), .Z(n79) );
  CLKBUF_X1 U101 ( .A(n24), .Z(n80) );
  CLKBUF_X1 U102 ( .A(n24), .Z(n81) );
  CLKBUF_X1 U103 ( .A(n24), .Z(n82) );
  CLKBUF_X1 U104 ( .A(n24), .Z(n83) );
  CLKBUF_X1 U105 ( .A(N33), .Z(n84) );
  CLKBUF_X1 U106 ( .A(N33), .Z(n85) );
  CLKBUF_X1 U107 ( .A(N33), .Z(n86) );
  CLKBUF_X1 U108 ( .A(N33), .Z(n87) );
  CLKBUF_X1 U109 ( .A(N33), .Z(n88) );
  CLKBUF_X1 U110 ( .A(N33), .Z(n89) );
  CLKBUF_X1 U111 ( .A(N26), .Z(n93) );
  CLKBUF_X1 U112 ( .A(N26), .Z(n94) );
  CLKBUF_X1 U113 ( .A(N26), .Z(n95) );
  CLKBUF_X1 U114 ( .A(N26), .Z(n96) );
  CLKBUF_X1 U115 ( .A(N26), .Z(n97) );
  CLKBUF_X1 U116 ( .A(N26), .Z(n98) );
endmodule


module CU_HW ( Clk, Rst, IR_IN, flush, JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, 
        CALL, RET, IMM_SEL, MUXA_SEL, MUXB_SEL, EQ_COND, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), SEL_STORE1, SEL_STORE0, SEL_LOAD2, SEL_LOAD1, 
        SEL_LOAD0, DRAM_WR, WB_MUX_SEL, RF_WR );
  input [31:0] IR_IN;
  input [1:0] flush;
  input Clk, Rst;
  output JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL, MUXA_SEL,
         MUXB_SEL, EQ_COND, \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] ,
         \ALU_OPCODE[1] , \ALU_OPCODE[0] , SEL_STORE1, SEL_STORE0, SEL_LOAD2,
         SEL_LOAD1, SEL_LOAD0, DRAM_WR, WB_MUX_SEL, RF_WR;

  assign JUMP_EN = 1'b0;
  assign RF_RD1_EN = 1'b0;
  assign RF_RD2_EN = 1'b0;
  assign RF_EN = 1'b0;
  assign CALL = 1'b0;
  assign RET = 1'b0;
  assign IMM_SEL = 1'b0;
  assign MUXA_SEL = 1'b0;
  assign MUXB_SEL = 1'b0;
  assign EQ_COND = 1'b0;
  assign \ALU_OPCODE[4]  = 1'b0;
  assign \ALU_OPCODE[3]  = 1'b0;
  assign \ALU_OPCODE[2]  = 1'b0;
  assign \ALU_OPCODE[1]  = 1'b0;
  assign \ALU_OPCODE[0]  = 1'b0;
  assign SEL_STORE1 = 1'b0;
  assign SEL_STORE0 = 1'b0;
  assign SEL_LOAD2 = 1'b0;
  assign SEL_LOAD1 = 1'b0;
  assign SEL_LOAD0 = 1'b0;
  assign DRAM_WR = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign RF_WR = 1'b0;

endmodule


module datapath ( Clk, Rst, Instr, JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, 
        RET, IMM_SEL, MUXA_SEL, MUXB_SEL, EQ_COND, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), SEL_STORE1, SEL_STORE0, SEL_LOAD2, SEL_LOAD1, 
        SEL_LOAD0, DRAM_WR, WB_MUX_SEL, RF_WR, flush, PC_out );
  input [31:0] Instr;
  output [1:0] flush;
  output [31:0] PC_out;
  input Clk, Rst, JUMP_EN, RF_RD1_EN, RF_RD2_EN, RF_EN, CALL, RET, IMM_SEL,
         MUXA_SEL, MUXB_SEL, EQ_COND, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , SEL_STORE1,
         SEL_STORE0, SEL_LOAD2, SEL_LOAD1, SEL_LOAD0, DRAM_WR, WB_MUX_SEL,
         RF_WR;
  wire   PC_out_31, PC_enable1, SPILL, FILL, JAL_op2, JAL_op4, PC_enable_fixed,
         JUMP_EN1, JUMP_EN2, BRANCH_op2, forward_branch, forward_branch1,
         forward_branch2, JR_op, BRANCH_op, JR_op1, PC_enable, LOAD_op1,
         STORE_op, bootstrap, JAL_op, JAL_op1, JAL_op3, BRANCH_op1, LOAD_op,
         LOAD_op2, STORE_op1, STORE_op2, FWD_A_mem_dec, FWD_A_exe_dec,
         FWD_A_wb_dec, FWD_B_mem_exe, FWD_B_exe_dec, FWD_B_wb_dec,
         FWD_B_exe_mem, FWD_B_exe_mem1, FWD_B_exe_mem2, FWD_B_wb_mem,
         FWD_B_wb_mem1, FWD_B_wb_mem2, FWD_B_mem_mem, FWD_B_mem_mem1,
         FWD_B_mem_mem2, FWD_B_lmd1_mem, FWD_B_lmd1_mem1, FWD_B_lmd1_mem2,
         FWD_exe_branch, FWD_exe_branch1, FWD_wb_branch, FWD_wb_branch1, n39,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n97, n98, n99, n100, n101, n102, n113,
         n210, n312, n313, n314, n330, n331, n332, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453;
  wire   [31:0] Instr_reg_out;
  wire   [5:0] OPCODE1;
  wire   [5:0] OPCODE2;
  wire   [4:0] RD;
  wire   [4:0] RD1;
  wire   [4:0] RD2;
  wire   [4:0] RD3;
  wire   [31:0] RF_write_data;
  wire   [31:0] RF_out_A;
  wire   [31:0] RF_out_B;
  wire   [31:0] fill_from_stack;
  wire   [31:0] A_reg_out;
  wire   [31:0] B_reg_out;
  wire   [31:0] Immediate_16_extended;
  wire   [31:0] Immediate_26_extended;
  wire   [31:0] Immediate_selected;
  wire   [31:0] Immediate_clocked;
  wire   [31:0] NPC2;
  wire   [31:0] ALU_operand_1;
  wire   [31:0] ALU_operand_2;
  wire   [4:0] ALU_OPCODE_in;
  wire   [31:0] ALU_operand_1_FWD;
  wire   [31:0] ALU_operand_2_FWD;
  wire   [31:0] ALU_output_FWD;
  wire   [31:0] ALU_reg_out;
  wire   [31:0] DRAM_write_data;
  wire   [31:0] DRAM_write_data_FWD;
  wire   [31:0] DRAM_read_data;
  wire   [31:0] LMD_reg_out;
  wire   [31:0] LMD_reg_out1;
  wire   [31:0] ALU_WB_out;
  wire   [31:0] ALU_WB_out1;
  wire   [31:0] WB_mux_out;
  wire   [31:0] NPC4;
  wire   [1:0] PC_reg_out;
  wire   [31:0] NPC;
  wire   [31:0] NPC1;
  wire   [31:0] NPC3;
  wire   [2:0] PC_mux_sel;
  wire   [31:0] PC_displaced;
  wire   [31:0] RF_out_A_FWD;
  wire   [31:16] PC_Immediate_displacement;
  wire   [1:0] flush0;
  wire   [1:0] flush2;
  wire   [2:0] FWD_A_sel;
  wire   [2:0] FWD_B_sel;
  tri   [31:0] spill_to_stack;
  tri   [31:0] ALU_output;
  tri   [31:0] PC_reg_in;
  assign PC_out[31] = PC_out_31;
  assign PC_out[30] = PC_out_31;
  assign PC_out[29] = PC_out_31;
  assign n39 = Rst;

  alu ALU_block ( .A(ALU_operand_1_FWD), .B(ALU_operand_2_FWD), .OP(
        ALU_OPCODE_in), .Y1(ALU_output) );
  cla_adder_N32 jump_adder ( .A(NPC), .B({PC_Immediate_displacement[31], 
        PC_Immediate_displacement[31], PC_Immediate_displacement[31], 
        PC_Immediate_displacement[31], PC_Immediate_displacement[31], 
        PC_Immediate_displacement[31], PC_Immediate_displacement[31], 
        PC_Immediate_displacement[24:16], Instr[15:0]}), .Ci(1'b0), .Sum(
        PC_displaced) );
  NAND3_X1 U456 ( .A1(Instr_reg_out[31]), .A2(Instr_reg_out[29]), .A3(n228), 
        .ZN(n109) );
  OAI33_X1 U457 ( .A1(n232), .A2(FWD_exe_branch1), .A3(n233), .B1(n234), .B2(
        n235), .B3(n236), .ZN(n231) );
  NAND3_X1 U458 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n296) );
  NAND3_X1 U459 ( .A1(Instr_reg_out[27]), .A2(n278), .A3(Instr_reg_out[26]), 
        .ZN(n311) );
  NAND3_X1 U460 ( .A1(n306), .A2(n307), .A3(n305), .ZN(n327) );
  XOR2_X1 U461 ( .A(RD2[0]), .B(Instr_reg_out[21]), .Z(n341) );
  XOR2_X1 U462 ( .A(RD2[1]), .B(Instr_reg_out[22]), .Z(n340) );
  XOR2_X1 U463 ( .A(RD1[0]), .B(Instr_reg_out[21]), .Z(n349) );
  XOR2_X1 U464 ( .A(RD1[1]), .B(Instr_reg_out[22]), .Z(n348) );
  reg_N32_0 IR ( .clk(Clk), .rst(n451), .d_in(Instr), .d_out(Instr_reg_out) );
  reg_N6_0 OPC1 ( .clk(Clk), .rst(n451), .d_in(Instr_reg_out[31:26]), .d_out(
        OPCODE1) );
  reg_N6_1 OPC2 ( .clk(Clk), .rst(n451), .d_in(OPCODE1), .d_out(OPCODE2) );
  reg_N5_0 RDreg1 ( .clk(Clk), .rst(n451), .d_in(RD), .d_out(RD1) );
  reg_N5_2 RDreg2 ( .clk(Clk), .rst(n451), .d_in(RD1), .d_out(RD2) );
  reg_N5_1 RDreg3 ( .clk(Clk), .rst(n451), .d_in(RD2), .d_out(RD3) );
  w_reg_file_M8_N8_F4_Nbit32 RF ( .clk(Clk), .reset(n451), .enable(RF_EN), 
        .rd1(RF_RD1_EN), .rd2(RF_RD2_EN), .wr(RF_WR), .add_wr(RD3), .add_rd1(
        Instr_reg_out[25:21]), .add_rd2(Instr_reg_out[20:16]), .datain(
        RF_write_data), .out1(RF_out_A), .out2(RF_out_B), .call(CALL), .ret(
        RET), .spill(SPILL), .fill(FILL), .to_mem(spill_to_stack), .from_mem(
        fill_from_stack) );
  stack WRF_stack ( .clk(Clk), .reset(n453), .enable(1'b1), .RD(FILL), .wr(
        SPILL), .datain(spill_to_stack), .dataout(fill_from_stack) );
  reg_N32_13 A ( .clk(Clk), .rst(n451), .d_in(RF_out_A), .d_out(A_reg_out) );
  reg_N32_12 B ( .clk(Clk), .rst(n452), .d_in(RF_out_B), .d_out(B_reg_out) );
  sign_ext_Nstart16_Nend32 Imm16ext ( .Ain(Instr_reg_out[15:0]), .Aout(
        Immediate_16_extended) );
  sign_ext_Nstart26_Nend32 Imm26ext ( .Ain(Instr_reg_out[25:0]), .Aout(
        Immediate_26_extended) );
  MUX21_GENERIC_N32_0 mux_imm ( .A(Immediate_16_extended), .B(
        Immediate_26_extended), .SEL(IMM_SEL), .Y(Immediate_selected) );
  reg_N32_11 Immreg ( .clk(Clk), .rst(n452), .d_in(Immediate_selected), 
        .d_out(Immediate_clocked) );
  MUX21_GENERIC_N32_4 MUX_A ( .A(NPC2), .B(A_reg_out), .SEL(MUXA_SEL), .Y(
        ALU_operand_1) );
  MUX21_GENERIC_N32_3 MUX_B ( .A(B_reg_out), .B(Immediate_clocked), .SEL(
        MUXB_SEL), .Y(ALU_operand_2) );
  reg_N32_10 ALU_REG ( .clk(Clk), .rst(n451), .d_in(ALU_output_FWD), .d_out(
        ALU_reg_out) );
  reg_N32_9 BREG ( .clk(Clk), .rst(n452), .d_in(B_reg_out), .d_out(
        DRAM_write_data) );
  DRAM dataram ( .clk(Clk), .rst(n453), .WR(DRAM_WR), .sel_store({SEL_STORE1, 
        SEL_STORE0}), .sel_load({SEL_LOAD2, SEL_LOAD1, SEL_LOAD0}), .addr(
        ALU_reg_out[11:0]), .d_in(DRAM_write_data_FWD), .d_out(DRAM_read_data)
         );
  reg_N32_8 LMD ( .clk(Clk), .rst(n452), .d_in(DRAM_read_data), .d_out(
        LMD_reg_out) );
  reg_N32_7 LMD1 ( .clk(Clk), .rst(n452), .d_in(LMD_reg_out), .d_out(
        LMD_reg_out1) );
  reg_N32_6 ALUWB ( .clk(Clk), .rst(n451), .d_in(ALU_reg_out), .d_out(
        ALU_WB_out) );
  reg_N32_5 ALUWB1 ( .clk(Clk), .rst(n451), .d_in(ALU_WB_out), .d_out(
        ALU_WB_out1) );
  MUX21_GENERIC_N32_2 mux_WB ( .A(LMD_reg_out), .B(ALU_WB_out), .SEL(
        WB_MUX_SEL), .Y(WB_mux_out) );
  MUX21_GENERIC_N32_1 RFin_mux ( .A(NPC4), .B(WB_mux_out), .SEL(JAL_op4), .Y(
        RF_write_data) );
  reg_en_N32 PC ( .clk(Clk), .rst(n451), .en(PC_enable_fixed), .d_in(PC_reg_in), .d_out({PC_out_31, PC_out[28:0], PC_reg_out}) );
  PC_incr PCi ( .PC({PC_out_31, PC_out[28:0], PC_reg_out}), .NPC(NPC) );
  reg_N32_4 NPCreg1 ( .clk(Clk), .rst(n451), .d_in(NPC), .d_out(NPC1) );
  reg_N32_3 NPCreg2 ( .clk(Clk), .rst(n452), .d_in(NPC1), .d_out(NPC2) );
  reg_N32_2 NPCreg3 ( .clk(Clk), .rst(n452), .d_in(NPC2), .d_out(NPC3) );
  reg_N32_1 NPCreg4 ( .clk(Clk), .rst(n452), .d_in(NPC3), .d_out(NPC4) );
  ff_0 JUMPENREG1 ( .clk(Clk), .rst(n452), .d_in(JUMP_EN), .d_out(JUMP_EN1) );
  ff_31 JUMPENREG2 ( .clk(Clk), .rst(n452), .d_in(JUMP_EN1), .d_out(JUMP_EN2)
         );
  ff_30 forward_branchREG1 ( .clk(Clk), .rst(n453), .d_in(forward_branch), 
        .d_out(forward_branch1) );
  ff_29 forward_branchREG2 ( .clk(Clk), .rst(n453), .d_in(forward_branch1), 
        .d_out(forward_branch2) );
  mux_pc pc_mux ( .A(NPC), .B(PC_displaced), .C(RF_out_A_FWD), .D(NPC2), .E(
        ALU_output_FWD), .F(NPC2), .sel({PC_mux_sel[2], flush0[0], 
        PC_mux_sel[0]}), .Y(PC_reg_in) );
  reg_N2_0 flushreg1 ( .clk(Clk), .rst(n452), .d_in(flush0), .d_out(flush) );
  reg_N2_1 flushreg2 ( .clk(Clk), .rst(n452), .d_in(flush), .d_out(flush2) );
  ff_28 pcen1 ( .clk(Clk), .rst(n453), .d_in(PC_enable), .d_out(PC_enable1) );
  counter cnt ( .clk(Clk), .rst(n452), .tc(bootstrap) );
  ff_27 JALreg1 ( .clk(Clk), .rst(n453), .d_in(JAL_op), .d_out(JAL_op1) );
  ff_26 JALreg2 ( .clk(Clk), .rst(n453), .d_in(JAL_op1), .d_out(JAL_op2) );
  ff_25 JALreg3 ( .clk(Clk), .rst(n453), .d_in(JAL_op2), .d_out(JAL_op3) );
  ff_24 JALreg4 ( .clk(Clk), .rst(n453), .d_in(JAL_op3), .d_out(JAL_op4) );
  ff_23 JRreg1 ( .clk(Clk), .rst(n453), .d_in(JR_op), .d_out(JR_op1) );
  ff_22 BRANCH_opREG1 ( .clk(Clk), .rst(n453), .d_in(BRANCH_op), .d_out(
        BRANCH_op1) );
  ff_21 BRANCH_opREG2 ( .clk(Clk), .rst(n453), .d_in(BRANCH_op1), .d_out(
        BRANCH_op2) );
  ff_20 LOADREG1 ( .clk(Clk), .rst(n452), .d_in(LOAD_op), .d_out(LOAD_op1) );
  ff_19 LOADREG2 ( .clk(Clk), .rst(n452), .d_in(LOAD_op1), .d_out(LOAD_op2) );
  ff_18 STOREREG1 ( .clk(Clk), .rst(n452), .d_in(STORE_op), .d_out(STORE_op1)
         );
  ff_17 STOREREG2 ( .clk(Clk), .rst(n452), .d_in(STORE_op1), .d_out(STORE_op2)
         );
  ff_16 FWDAREG3 ( .clk(Clk), .rst(n452), .d_in(FWD_A_mem_dec), .d_out(
        FWD_A_sel[0]) );
  ff_15 FWDAREG ( .clk(Clk), .rst(n452), .d_in(FWD_A_exe_dec), .d_out(
        FWD_A_sel[2]) );
  ff_14 FWDAREG2 ( .clk(Clk), .rst(n452), .d_in(FWD_A_wb_dec), .d_out(
        FWD_A_sel[1]) );
  mux_fwd_0 FWDAMUX ( .OP(ALU_operand_1), .alu_out(ALU_reg_out), .alu_wb_in(
        ALU_WB_out), .lmd_out(LMD_reg_out), .OPF(ALU_operand_1_FWD), .sel(
        FWD_A_sel) );
  ff_13 FWDBREG3a ( .clk(Clk), .rst(n452), .d_in(FWD_B_mem_exe), .d_out(
        FWD_B_sel[0]) );
  ff_12 FWDBREG ( .clk(Clk), .rst(n452), .d_in(FWD_B_exe_dec), .d_out(
        FWD_B_sel[2]) );
  ff_11 FWDBREG2 ( .clk(Clk), .rst(n452), .d_in(FWD_B_wb_dec), .d_out(
        FWD_B_sel[1]) );
  mux_fwd_1 FWDBMUX ( .OP(ALU_operand_2), .alu_out(ALU_reg_out), .alu_wb_in(
        ALU_WB_out), .lmd_out(LMD_reg_out), .OPF(ALU_operand_2_FWD), .sel(
        FWD_B_sel) );
  ff_10 FWDBREG3 ( .clk(Clk), .rst(n452), .d_in(FWD_B_exe_mem), .d_out(
        FWD_B_exe_mem1) );
  ff_9 FWDBREG4 ( .clk(Clk), .rst(n452), .d_in(FWD_B_exe_mem1), .d_out(
        FWD_B_exe_mem2) );
  ff_8 FWDBREG5 ( .clk(Clk), .rst(n452), .d_in(FWD_B_wb_mem), .d_out(
        FWD_B_wb_mem1) );
  ff_7 FWDBREG6 ( .clk(Clk), .rst(n452), .d_in(FWD_B_wb_mem1), .d_out(
        FWD_B_wb_mem2) );
  ff_6 FWDBREG7 ( .clk(Clk), .rst(n452), .d_in(FWD_B_mem_mem), .d_out(
        FWD_B_mem_mem1) );
  ff_5 FWDBREG8 ( .clk(Clk), .rst(n452), .d_in(FWD_B_mem_mem1), .d_out(
        FWD_B_mem_mem2) );
  ff_4 FWDBREG9 ( .clk(Clk), .rst(n452), .d_in(FWD_B_lmd1_mem), .d_out(
        FWD_B_lmd1_mem1) );
  ff_3 FWDBREG10 ( .clk(Clk), .rst(n452), .d_in(FWD_B_lmd1_mem1), .d_out(
        FWD_B_lmd1_mem2) );
  ff_2 FWDBRANCH1 ( .clk(Clk), .rst(n452), .d_in(FWD_exe_branch), .d_out(
        FWD_exe_branch1) );
  ff_1 FWDBRANCH2 ( .clk(Clk), .rst(n452), .d_in(FWD_wb_branch), .d_out(
        FWD_wb_branch1) );
  NOR4_X1 U3 ( .A1(RD2[3]), .A2(RD2[4]), .A3(RD2[2]), .A4(n342), .ZN(n290) );
  BUF_X1 U4 ( .A(n110), .Z(n434) );
  BUF_X1 U5 ( .A(n110), .Z(n435) );
  INV_X1 U6 ( .A(n449), .ZN(n440) );
  BUF_X1 U7 ( .A(n110), .Z(n436) );
  BUF_X1 U8 ( .A(n115), .Z(n429) );
  BUF_X1 U9 ( .A(n115), .Z(n430) );
  BUF_X1 U10 ( .A(n115), .Z(n431) );
  BUF_X1 U11 ( .A(n450), .Z(n449) );
  NAND2_X1 U12 ( .A1(n209), .A2(n432), .ZN(n110) );
  BUF_X1 U13 ( .A(n446), .Z(n447) );
  BUF_X1 U14 ( .A(n445), .Z(n448) );
  BUF_X1 U15 ( .A(n450), .Z(n445) );
  BUF_X1 U16 ( .A(n450), .Z(n446) );
  BUF_X1 U17 ( .A(n450), .Z(n444) );
  BUF_X1 U18 ( .A(n450), .Z(n441) );
  BUF_X1 U19 ( .A(n450), .Z(n443) );
  BUF_X1 U20 ( .A(n450), .Z(n442) );
  BUF_X1 U21 ( .A(n355), .Z(n210) );
  BUF_X1 U22 ( .A(n355), .Z(n312) );
  BUF_X1 U23 ( .A(n355), .Z(n313) );
  AOI21_X1 U24 ( .B1(n106), .B2(n107), .A(n108), .ZN(flush0[0]) );
  INV_X1 U25 ( .A(n97), .ZN(n432) );
  INV_X1 U26 ( .A(n97), .ZN(n433) );
  NOR2_X1 U27 ( .A1(n209), .A2(n97), .ZN(n115) );
  OAI21_X1 U28 ( .B1(n218), .B2(PC_enable), .A(n107), .ZN(n103) );
  NOR2_X1 U29 ( .A1(n212), .A2(n106), .ZN(n209) );
  INV_X1 U30 ( .A(n221), .ZN(PC_mux_sel[0]) );
  AOI21_X1 U31 ( .B1(n106), .B2(n103), .A(n108), .ZN(n221) );
  INV_X1 U32 ( .A(n104), .ZN(PC_mux_sel[2]) );
  INV_X1 U33 ( .A(n230), .ZN(n211) );
  INV_X1 U34 ( .A(n120), .ZN(ALU_output_FWD[7]) );
  INV_X1 U35 ( .A(n162), .ZN(ALU_output_FWD[23]) );
  INV_X1 U36 ( .A(n168), .ZN(ALU_output_FWD[21]) );
  INV_X1 U37 ( .A(n180), .ZN(ALU_output_FWD[18]) );
  INV_X1 U38 ( .A(n186), .ZN(ALU_output_FWD[16]) );
  INV_X1 U39 ( .A(n189), .ZN(ALU_output_FWD[15]) );
  INV_X1 U40 ( .A(n192), .ZN(ALU_output_FWD[14]) );
  INV_X1 U41 ( .A(n195), .ZN(ALU_output_FWD[13]) );
  INV_X1 U42 ( .A(n198), .ZN(ALU_output_FWD[12]) );
  INV_X1 U43 ( .A(n201), .ZN(ALU_output_FWD[11]) );
  INV_X1 U44 ( .A(n204), .ZN(ALU_output_FWD[10]) );
  INV_X1 U45 ( .A(n174), .ZN(ALU_output_FWD[1]) );
  INV_X1 U46 ( .A(n207), .ZN(ALU_output_FWD[0]) );
  INV_X1 U47 ( .A(n147), .ZN(ALU_output_FWD[28]) );
  INV_X1 U48 ( .A(n153), .ZN(ALU_output_FWD[26]) );
  INV_X1 U49 ( .A(n159), .ZN(ALU_output_FWD[24]) );
  INV_X1 U50 ( .A(n165), .ZN(ALU_output_FWD[22]) );
  INV_X1 U51 ( .A(n171), .ZN(ALU_output_FWD[20]) );
  INV_X1 U52 ( .A(n177), .ZN(ALU_output_FWD[19]) );
  INV_X1 U53 ( .A(n183), .ZN(ALU_output_FWD[17]) );
  INV_X1 U54 ( .A(n117), .ZN(ALU_output_FWD[8]) );
  INV_X1 U55 ( .A(n123), .ZN(ALU_output_FWD[6]) );
  INV_X1 U56 ( .A(n129), .ZN(ALU_output_FWD[4]) );
  INV_X1 U57 ( .A(n141), .ZN(ALU_output_FWD[2]) );
  INV_X1 U58 ( .A(n150), .ZN(ALU_output_FWD[27]) );
  INV_X1 U59 ( .A(n156), .ZN(ALU_output_FWD[25]) );
  INV_X1 U60 ( .A(n112), .ZN(ALU_output_FWD[9]) );
  INV_X1 U61 ( .A(n126), .ZN(ALU_output_FWD[5]) );
  INV_X1 U62 ( .A(n132), .ZN(ALU_output_FWD[3]) );
  INV_X1 U63 ( .A(n138), .ZN(ALU_output_FWD[30]) );
  INV_X1 U64 ( .A(n144), .ZN(ALU_output_FWD[29]) );
  INV_X1 U65 ( .A(n135), .ZN(ALU_output_FWD[31]) );
  OAI21_X1 U66 ( .B1(n103), .B2(n104), .A(n105), .ZN(flush0[1]) );
  INV_X1 U67 ( .A(flush0[0]), .ZN(n105) );
  INV_X1 U68 ( .A(n304), .ZN(n303) );
  INV_X1 U69 ( .A(n216), .ZN(RD[1]) );
  INV_X1 U70 ( .A(n215), .ZN(RD[2]) );
  INV_X1 U71 ( .A(n109), .ZN(STORE_op) );
  NOR3_X1 U72 ( .A1(n335), .A2(n290), .A3(n212), .ZN(FWD_A_mem_dec) );
  NOR3_X1 U73 ( .A1(n327), .A2(n304), .A3(n328), .ZN(FWD_B_exe_dec) );
  INV_X1 U74 ( .A(n308), .ZN(FWD_B_lmd1_mem) );
  NOR2_X1 U75 ( .A1(n230), .A2(n284), .ZN(FWD_exe_branch) );
  NOR2_X1 U76 ( .A1(n212), .A2(n284), .ZN(FWD_wb_branch) );
  INV_X1 U77 ( .A(n213), .ZN(RD[4]) );
  INV_X1 U78 ( .A(n217), .ZN(RD[0]) );
  INV_X1 U79 ( .A(n214), .ZN(RD[3]) );
  INV_X1 U80 ( .A(JAL_op2), .ZN(n450) );
  BUF_X1 U81 ( .A(n353), .Z(n332) );
  BUF_X1 U82 ( .A(n353), .Z(n424) );
  NOR2_X1 U83 ( .A1(n420), .A2(n418), .ZN(n355) );
  BUF_X1 U84 ( .A(n354), .Z(n314) );
  BUF_X1 U85 ( .A(n354), .Z(n330) );
  BUF_X1 U86 ( .A(n352), .Z(n426) );
  BUF_X1 U87 ( .A(n352), .Z(n427) );
  BUF_X1 U88 ( .A(n353), .Z(n425) );
  BUF_X1 U89 ( .A(n354), .Z(n331) );
  BUF_X1 U90 ( .A(n352), .Z(n428) );
  INV_X1 U91 ( .A(n419), .ZN(n418) );
  OAI22_X1 U92 ( .A1(Instr_reg_out[20]), .A2(n322), .B1(Instr_reg_out[15]), 
        .B2(n304), .ZN(n213) );
  OAI22_X1 U93 ( .A1(Instr_reg_out[19]), .A2(n322), .B1(Instr_reg_out[14]), 
        .B2(n304), .ZN(n214) );
  OAI22_X1 U94 ( .A1(Instr_reg_out[18]), .A2(n322), .B1(Instr_reg_out[13]), 
        .B2(n304), .ZN(n215) );
  OAI22_X1 U95 ( .A1(Instr_reg_out[16]), .A2(n322), .B1(Instr_reg_out[11]), 
        .B2(n304), .ZN(n217) );
  OAI22_X1 U96 ( .A1(Instr_reg_out[17]), .A2(n322), .B1(Instr_reg_out[12]), 
        .B2(n304), .ZN(n216) );
  NOR3_X1 U97 ( .A1(n222), .A2(JR_op), .A3(n223), .ZN(n108) );
  AOI21_X1 U98 ( .B1(Instr[15]), .B2(BRANCH_op), .A(JUMP_EN), .ZN(n222) );
  INV_X1 U99 ( .A(n224), .ZN(n223) );
  OAI221_X1 U100 ( .B1(n435), .B2(n137), .C1(n138), .C2(n433), .A(n139), .ZN(
        RF_out_A_FWD[30]) );
  OAI221_X1 U101 ( .B1(n435), .B2(n143), .C1(n144), .C2(n433), .A(n145), .ZN(
        RF_out_A_FWD[29]) );
  OAI221_X1 U102 ( .B1(n435), .B2(n161), .C1(n162), .C2(n433), .A(n163), .ZN(
        RF_out_A_FWD[23]) );
  OAI221_X1 U103 ( .B1(n435), .B2(n146), .C1(n147), .C2(n433), .A(n148), .ZN(
        RF_out_A_FWD[28]) );
  OAI221_X1 U104 ( .B1(n435), .B2(n152), .C1(n153), .C2(n433), .A(n154), .ZN(
        RF_out_A_FWD[26]) );
  OAI221_X1 U105 ( .B1(n435), .B2(n158), .C1(n159), .C2(n433), .A(n160), .ZN(
        RF_out_A_FWD[24]) );
  OAI221_X1 U106 ( .B1(n435), .B2(n149), .C1(n150), .C2(n433), .A(n151), .ZN(
        RF_out_A_FWD[27]) );
  OAI221_X1 U107 ( .B1(n435), .B2(n155), .C1(n156), .C2(n433), .A(n157), .ZN(
        RF_out_A_FWD[25]) );
  NOR4_X1 U108 ( .A1(ALU_reg_out[22]), .A2(ALU_reg_out[21]), .A3(
        ALU_reg_out[20]), .A4(ALU_reg_out[1]), .ZN(n244) );
  NOR4_X1 U109 ( .A1(A_reg_out[9]), .A2(A_reg_out[8]), .A3(A_reg_out[7]), .A4(
        A_reg_out[6]), .ZN(n261) );
  NOR4_X1 U110 ( .A1(A_reg_out[23]), .A2(A_reg_out[22]), .A3(A_reg_out[21]), 
        .A4(A_reg_out[20]), .ZN(n265) );
  NOR4_X1 U111 ( .A1(A_reg_out[5]), .A2(A_reg_out[4]), .A3(A_reg_out[3]), .A4(
        A_reg_out[31]), .ZN(n260) );
  NOR4_X1 U112 ( .A1(A_reg_out[1]), .A2(A_reg_out[19]), .A3(A_reg_out[18]), 
        .A4(A_reg_out[17]), .ZN(n264) );
  AOI21_X1 U113 ( .B1(n245), .B2(n246), .A(n247), .ZN(n233) );
  INV_X1 U114 ( .A(FWD_wb_branch1), .ZN(n247) );
  NOR4_X1 U115 ( .A1(n252), .A2(n253), .A3(n254), .A4(n255), .ZN(n245) );
  NOR4_X1 U116 ( .A1(n248), .A2(n249), .A3(n250), .A4(n251), .ZN(n246) );
  NOR4_X1 U117 ( .A1(ALU_reg_out[19]), .A2(ALU_reg_out[18]), .A3(
        ALU_reg_out[17]), .A4(ALU_reg_out[16]), .ZN(n243) );
  NOR4_X1 U118 ( .A1(ALU_reg_out[2]), .A2(ALU_reg_out[29]), .A3(
        ALU_reg_out[28]), .A4(ALU_reg_out[27]), .ZN(n238) );
  NOR4_X1 U119 ( .A1(ALU_reg_out[15]), .A2(ALU_reg_out[14]), .A3(
        ALU_reg_out[13]), .A4(ALU_reg_out[12]), .ZN(n242) );
  NOR4_X1 U120 ( .A1(A_reg_out[30]), .A2(A_reg_out[2]), .A3(A_reg_out[29]), 
        .A4(A_reg_out[28]), .ZN(n259) );
  NOR4_X1 U121 ( .A1(A_reg_out[16]), .A2(A_reg_out[15]), .A3(A_reg_out[14]), 
        .A4(A_reg_out[13]), .ZN(n263) );
  NOR4_X1 U122 ( .A1(ALU_reg_out[26]), .A2(ALU_reg_out[25]), .A3(
        ALU_reg_out[24]), .A4(ALU_reg_out[23]), .ZN(n237) );
  NOR4_X1 U123 ( .A1(A_reg_out[27]), .A2(A_reg_out[26]), .A3(A_reg_out[25]), 
        .A4(A_reg_out[24]), .ZN(n258) );
  BUF_X2 U124 ( .A(n39), .Z(n451) );
  NAND4_X1 U125 ( .A1(n336), .A2(n337), .A3(n338), .A4(n339), .ZN(n212) );
  XNOR2_X1 U126 ( .A(Instr_reg_out[23]), .B(RD2[2]), .ZN(n336) );
  XNOR2_X1 U127 ( .A(Instr_reg_out[24]), .B(RD2[3]), .ZN(n338) );
  NOR2_X1 U128 ( .A1(n340), .A2(n341), .ZN(n339) );
  NOR3_X1 U129 ( .A1(Instr[31]), .A2(Instr[29]), .A3(n423), .ZN(n282) );
  INV_X1 U130 ( .A(PC_enable1), .ZN(n423) );
  NAND2_X1 U131 ( .A1(n304), .A2(n326), .ZN(n322) );
  OR3_X1 U132 ( .A1(Instr_reg_out[28]), .A2(Instr_reg_out[29]), .A3(n311), 
        .ZN(n326) );
  AND2_X1 U133 ( .A1(ALU_OPCODE[2]), .A2(PC_enable1), .ZN(ALU_OPCODE_in[2]) );
  AOI22_X1 U134 ( .A1(ALU_output[16]), .A2(n447), .B1(NPC2[16]), .B2(JAL_op2), 
        .ZN(n186) );
  AOI22_X1 U135 ( .A1(ALU_output[15]), .A2(n447), .B1(NPC2[15]), .B2(JAL_op2), 
        .ZN(n189) );
  AOI22_X1 U136 ( .A1(ALU_output[14]), .A2(n447), .B1(NPC2[14]), .B2(JAL_op2), 
        .ZN(n192) );
  AOI22_X1 U137 ( .A1(ALU_output[13]), .A2(n447), .B1(NPC2[13]), .B2(n440), 
        .ZN(n195) );
  AOI22_X1 U138 ( .A1(ALU_output[12]), .A2(n448), .B1(NPC2[12]), .B2(JAL_op2), 
        .ZN(n198) );
  AOI22_X1 U139 ( .A1(ALU_output[11]), .A2(n448), .B1(NPC2[11]), .B2(n440), 
        .ZN(n201) );
  AOI22_X1 U140 ( .A1(ALU_output[10]), .A2(n448), .B1(NPC2[10]), .B2(JAL_op2), 
        .ZN(n204) );
  AOI22_X1 U141 ( .A1(ALU_output[0]), .A2(n448), .B1(NPC2[0]), .B2(n440), .ZN(
        n207) );
  AOI22_X1 U142 ( .A1(ALU_output[23]), .A2(n445), .B1(NPC2[23]), .B2(n440), 
        .ZN(n162) );
  AOI22_X1 U143 ( .A1(ALU_output[21]), .A2(n445), .B1(NPC2[21]), .B2(n440), 
        .ZN(n168) );
  AOI22_X1 U144 ( .A1(ALU_output[18]), .A2(n446), .B1(NPC2[18]), .B2(n440), 
        .ZN(n180) );
  AOI22_X1 U145 ( .A1(ALU_output[1]), .A2(n446), .B1(NPC2[1]), .B2(n440), .ZN(
        n174) );
  AOI22_X1 U146 ( .A1(ALU_output[28]), .A2(n443), .B1(NPC2[28]), .B2(JAL_op2), 
        .ZN(n147) );
  AOI22_X1 U147 ( .A1(ALU_output[26]), .A2(n444), .B1(NPC2[26]), .B2(n440), 
        .ZN(n153) );
  AOI22_X1 U148 ( .A1(ALU_output[24]), .A2(n444), .B1(NPC2[24]), .B2(n440), 
        .ZN(n159) );
  AOI22_X1 U149 ( .A1(ALU_output[22]), .A2(n445), .B1(NPC2[22]), .B2(n440), 
        .ZN(n165) );
  AOI22_X1 U150 ( .A1(ALU_output[20]), .A2(n445), .B1(NPC2[20]), .B2(n440), 
        .ZN(n171) );
  AOI22_X1 U151 ( .A1(ALU_output[19]), .A2(n446), .B1(NPC2[19]), .B2(n440), 
        .ZN(n177) );
  AOI22_X1 U152 ( .A1(ALU_output[17]), .A2(n446), .B1(NPC2[17]), .B2(n440), 
        .ZN(n183) );
  AOI22_X1 U153 ( .A1(ALU_output[8]), .A2(n441), .B1(NPC2[8]), .B2(n440), .ZN(
        n117) );
  AOI22_X1 U154 ( .A1(ALU_output[6]), .A2(n441), .B1(NPC2[6]), .B2(JAL_op2), 
        .ZN(n123) );
  AOI22_X1 U155 ( .A1(ALU_output[4]), .A2(n442), .B1(NPC2[4]), .B2(JAL_op2), 
        .ZN(n129) );
  AOI22_X1 U156 ( .A1(ALU_output[2]), .A2(n443), .B1(NPC2[2]), .B2(JAL_op2), 
        .ZN(n141) );
  AOI22_X1 U157 ( .A1(ALU_output[27]), .A2(n444), .B1(NPC2[27]), .B2(n440), 
        .ZN(n150) );
  AOI22_X1 U158 ( .A1(ALU_output[25]), .A2(n444), .B1(NPC2[25]), .B2(n440), 
        .ZN(n156) );
  AOI22_X1 U159 ( .A1(ALU_output[9]), .A2(n441), .B1(NPC2[9]), .B2(n440), .ZN(
        n112) );
  AOI22_X1 U160 ( .A1(ALU_output[7]), .A2(n441), .B1(NPC2[7]), .B2(JAL_op2), 
        .ZN(n120) );
  AOI22_X1 U161 ( .A1(ALU_output[5]), .A2(n442), .B1(NPC2[5]), .B2(JAL_op2), 
        .ZN(n126) );
  AOI22_X1 U162 ( .A1(ALU_output[3]), .A2(n442), .B1(NPC2[3]), .B2(JAL_op2), 
        .ZN(n132) );
  AOI22_X1 U163 ( .A1(ALU_output[30]), .A2(n443), .B1(NPC2[30]), .B2(JAL_op2), 
        .ZN(n138) );
  AOI22_X1 U164 ( .A1(ALU_output[29]), .A2(n443), .B1(NPC2[29]), .B2(JAL_op2), 
        .ZN(n144) );
  AOI22_X1 U165 ( .A1(ALU_output[31]), .A2(n442), .B1(NPC2[31]), .B2(n440), 
        .ZN(n135) );
  AND2_X1 U166 ( .A1(ALU_OPCODE[0]), .A2(PC_enable1), .ZN(ALU_OPCODE_in[0]) );
  NAND4_X1 U167 ( .A1(n280), .A2(n279), .A3(n229), .A4(n329), .ZN(n304) );
  NOR3_X1 U168 ( .A1(Instr_reg_out[29]), .A2(Instr_reg_out[31]), .A3(
        Instr_reg_out[30]), .ZN(n329) );
  OAI211_X1 U169 ( .C1(n218), .C2(n219), .A(n107), .B(n220), .ZN(n104) );
  INV_X1 U170 ( .A(PC_enable), .ZN(n219) );
  NOR2_X1 U171 ( .A1(JR_op1), .A2(n108), .ZN(n220) );
  AOI22_X1 U172 ( .A1(LOAD_op1), .A2(n211), .B1(n109), .B2(FWD_B_mem_mem), 
        .ZN(n224) );
  NAND4_X1 U173 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .ZN(n230) );
  XNOR2_X1 U174 ( .A(Instr_reg_out[23]), .B(RD1[2]), .ZN(n344) );
  XNOR2_X1 U175 ( .A(Instr_reg_out[24]), .B(RD1[3]), .ZN(n346) );
  XNOR2_X1 U176 ( .A(Instr_reg_out[25]), .B(RD1[4]), .ZN(n345) );
  NOR2_X1 U177 ( .A1(SPILL), .A2(FILL), .ZN(PC_enable) );
  XNOR2_X1 U178 ( .A(Instr_reg_out[25]), .B(RD2[4]), .ZN(n337) );
  NOR3_X1 U179 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n286) );
  XNOR2_X1 U180 ( .A(RD2[2]), .B(n215), .ZN(n289) );
  XNOR2_X1 U181 ( .A(RD2[3]), .B(n214), .ZN(n291) );
  NOR3_X1 U182 ( .A1(n319), .A2(n320), .A3(n321), .ZN(n316) );
  XNOR2_X1 U183 ( .A(RD1[4]), .B(n213), .ZN(n319) );
  XNOR2_X1 U184 ( .A(RD1[3]), .B(n214), .ZN(n321) );
  NOR3_X1 U185 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n285) );
  XNOR2_X1 U186 ( .A(RD2[1]), .B(n216), .ZN(n292) );
  XNOR2_X1 U187 ( .A(RD2[0]), .B(n217), .ZN(n293) );
  XNOR2_X1 U188 ( .A(RD2[4]), .B(n213), .ZN(n294) );
  XNOR2_X1 U189 ( .A(Instr_reg_out[20]), .B(RD1[4]), .ZN(n307) );
  XNOR2_X1 U190 ( .A(Instr_reg_out[19]), .B(RD1[3]), .ZN(n306) );
  AOI211_X1 U191 ( .C1(Instr_reg_out[27]), .C2(n229), .A(Instr_reg_out[30]), 
        .B(Instr_reg_out[28]), .ZN(n228) );
  AND2_X1 U192 ( .A1(JR_op1), .A2(n211), .ZN(n97) );
  XNOR2_X1 U193 ( .A(n231), .B(EQ_COND), .ZN(n226) );
  NAND2_X1 U194 ( .A1(n237), .A2(n238), .ZN(n236) );
  NAND4_X1 U195 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n234) );
  AND2_X1 U196 ( .A1(ALU_OPCODE[1]), .A2(PC_enable1), .ZN(ALU_OPCODE_in[1]) );
  NOR3_X1 U197 ( .A1(n323), .A2(n324), .A3(n325), .ZN(n315) );
  XNOR2_X1 U198 ( .A(RD1[1]), .B(n216), .ZN(n323) );
  XNOR2_X1 U199 ( .A(RD1[0]), .B(n217), .ZN(n324) );
  XNOR2_X1 U200 ( .A(RD1[2]), .B(n215), .ZN(n325) );
  AND2_X1 U201 ( .A1(ALU_OPCODE[4]), .A2(PC_enable1), .ZN(ALU_OPCODE_in[4]) );
  AND2_X1 U202 ( .A1(ALU_OPCODE[3]), .A2(PC_enable1), .ZN(ALU_OPCODE_in[3]) );
  AOI21_X1 U203 ( .B1(n256), .B2(n257), .A(FWD_wb_branch1), .ZN(n232) );
  AND4_X1 U204 ( .A1(n262), .A2(n263), .A3(n264), .A4(n265), .ZN(n256) );
  AND4_X1 U205 ( .A1(n258), .A2(n259), .A3(n260), .A4(n261), .ZN(n257) );
  NOR4_X1 U206 ( .A1(A_reg_out[12]), .A2(A_reg_out[11]), .A3(A_reg_out[10]), 
        .A4(A_reg_out[0]), .ZN(n262) );
  NOR2_X1 U207 ( .A1(n348), .A2(n349), .ZN(n347) );
  AND2_X1 U208 ( .A1(n224), .A2(n225), .ZN(n107) );
  OR3_X1 U209 ( .A1(n226), .A2(forward_branch2), .A3(n227), .ZN(n225) );
  INV_X1 U210 ( .A(BRANCH_op2), .ZN(n227) );
  OR4_X1 U211 ( .A1(ALU_WB_out[24]), .A2(ALU_WB_out[25]), .A3(ALU_WB_out[26]), 
        .A4(ALU_WB_out[27]), .ZN(n251) );
  OR4_X1 U212 ( .A1(ALU_WB_out[0]), .A2(ALU_WB_out[10]), .A3(ALU_WB_out[11]), 
        .A4(ALU_WB_out[12]), .ZN(n255) );
  OR4_X1 U213 ( .A1(ALU_WB_out[28]), .A2(ALU_WB_out[29]), .A3(ALU_WB_out[2]), 
        .A4(ALU_WB_out[30]), .ZN(n250) );
  OR4_X1 U214 ( .A1(ALU_WB_out[13]), .A2(ALU_WB_out[14]), .A3(ALU_WB_out[15]), 
        .A4(ALU_WB_out[16]), .ZN(n254) );
  OR4_X1 U215 ( .A1(ALU_WB_out[31]), .A2(ALU_WB_out[3]), .A3(ALU_WB_out[4]), 
        .A4(ALU_WB_out[5]), .ZN(n249) );
  OR4_X1 U216 ( .A1(ALU_WB_out[17]), .A2(ALU_WB_out[18]), .A3(ALU_WB_out[19]), 
        .A4(ALU_WB_out[1]), .ZN(n253) );
  OR4_X1 U217 ( .A1(ALU_WB_out[6]), .A2(ALU_WB_out[7]), .A3(ALU_WB_out[8]), 
        .A4(ALU_WB_out[9]), .ZN(n248) );
  OR4_X1 U218 ( .A1(ALU_WB_out[20]), .A2(ALU_WB_out[21]), .A3(ALU_WB_out[22]), 
        .A4(ALU_WB_out[23]), .ZN(n252) );
  INV_X1 U219 ( .A(Instr_reg_out[28]), .ZN(n279) );
  NAND4_X1 U220 ( .A1(n125), .A2(n122), .A3(n239), .A4(n240), .ZN(n235) );
  NOR3_X1 U221 ( .A1(ALU_reg_out[7]), .A2(ALU_reg_out[9]), .A3(ALU_reg_out[8]), 
        .ZN(n239) );
  NOR4_X1 U222 ( .A1(ALU_reg_out[4]), .A2(ALU_reg_out[3]), .A3(ALU_reg_out[31]), .A4(ALU_reg_out[30]), .ZN(n240) );
  INV_X1 U223 ( .A(JR_op1), .ZN(n106) );
  OAI221_X1 U224 ( .B1(n434), .B2(n173), .C1(n174), .C2(n432), .A(n175), .ZN(
        RF_out_A_FWD[1]) );
  OAI221_X1 U225 ( .B1(n434), .B2(n206), .C1(n207), .C2(n432), .A(n208), .ZN(
        RF_out_A_FWD[0]) );
  OAI221_X1 U226 ( .B1(n436), .B2(n122), .C1(n123), .C2(n433), .A(n124), .ZN(
        RF_out_A_FWD[6]) );
  OAI221_X1 U227 ( .B1(n436), .B2(n128), .C1(n129), .C2(n433), .A(n130), .ZN(
        RF_out_A_FWD[4]) );
  OAI221_X1 U228 ( .B1(n435), .B2(n140), .C1(n141), .C2(n433), .A(n142), .ZN(
        RF_out_A_FWD[2]) );
  OAI221_X1 U229 ( .B1(n436), .B2(n119), .C1(n120), .C2(n433), .A(n121), .ZN(
        RF_out_A_FWD[7]) );
  OAI221_X1 U230 ( .B1(n436), .B2(n125), .C1(n126), .C2(n433), .A(n127), .ZN(
        RF_out_A_FWD[5]) );
  OAI221_X1 U231 ( .B1(n436), .B2(n131), .C1(n132), .C2(n433), .A(n133), .ZN(
        RF_out_A_FWD[3]) );
  OAI221_X1 U232 ( .B1(n436), .B2(n134), .C1(n135), .C2(n433), .A(n136), .ZN(
        RF_out_A_FWD[31]) );
  OAI221_X1 U233 ( .B1(n435), .B2(n167), .C1(n168), .C2(n433), .A(n169), .ZN(
        RF_out_A_FWD[21]) );
  OAI221_X1 U234 ( .B1(n434), .B2(n179), .C1(n180), .C2(n432), .A(n181), .ZN(
        RF_out_A_FWD[18]) );
  OAI221_X1 U235 ( .B1(n434), .B2(n185), .C1(n186), .C2(n432), .A(n187), .ZN(
        RF_out_A_FWD[16]) );
  OAI221_X1 U236 ( .B1(n434), .B2(n188), .C1(n189), .C2(n432), .A(n190), .ZN(
        RF_out_A_FWD[15]) );
  OAI221_X1 U237 ( .B1(n434), .B2(n191), .C1(n192), .C2(n432), .A(n193), .ZN(
        RF_out_A_FWD[14]) );
  OAI221_X1 U238 ( .B1(n434), .B2(n194), .C1(n195), .C2(n432), .A(n196), .ZN(
        RF_out_A_FWD[13]) );
  OAI221_X1 U239 ( .B1(n434), .B2(n197), .C1(n198), .C2(n432), .A(n199), .ZN(
        RF_out_A_FWD[12]) );
  OAI221_X1 U240 ( .B1(n434), .B2(n200), .C1(n201), .C2(n432), .A(n202), .ZN(
        RF_out_A_FWD[11]) );
  OAI221_X1 U241 ( .B1(n434), .B2(n203), .C1(n204), .C2(n432), .A(n205), .ZN(
        RF_out_A_FWD[10]) );
  OAI221_X1 U242 ( .B1(n435), .B2(n164), .C1(n165), .C2(n433), .A(n166), .ZN(
        RF_out_A_FWD[22]) );
  OAI221_X1 U243 ( .B1(n435), .B2(n170), .C1(n171), .C2(n433), .A(n172), .ZN(
        RF_out_A_FWD[20]) );
  OAI221_X1 U244 ( .B1(n434), .B2(n176), .C1(n177), .C2(n432), .A(n178), .ZN(
        RF_out_A_FWD[19]) );
  OAI221_X1 U245 ( .B1(n434), .B2(n182), .C1(n183), .C2(n432), .A(n184), .ZN(
        RF_out_A_FWD[17]) );
  OAI221_X1 U246 ( .B1(n436), .B2(n116), .C1(n117), .C2(n433), .A(n118), .ZN(
        RF_out_A_FWD[8]) );
  OAI221_X1 U247 ( .B1(n436), .B2(n111), .C1(n112), .C2(n433), .A(n114), .ZN(
        RF_out_A_FWD[9]) );
  AND3_X1 U248 ( .A1(BRANCH_op2), .A2(n226), .A3(forward_branch2), .ZN(n218)
         );
  NAND2_X1 U249 ( .A1(RF_out_A[8]), .A2(n431), .ZN(n118) );
  NAND2_X1 U250 ( .A1(RF_out_A[6]), .A2(n431), .ZN(n124) );
  NAND2_X1 U251 ( .A1(RF_out_A[4]), .A2(n431), .ZN(n130) );
  NAND2_X1 U252 ( .A1(RF_out_A[9]), .A2(n431), .ZN(n114) );
  NAND2_X1 U253 ( .A1(RF_out_A[7]), .A2(n431), .ZN(n121) );
  NAND2_X1 U254 ( .A1(RF_out_A[5]), .A2(n431), .ZN(n127) );
  NAND2_X1 U255 ( .A1(RF_out_A[3]), .A2(n431), .ZN(n133) );
  NAND2_X1 U256 ( .A1(RF_out_A[31]), .A2(n431), .ZN(n136) );
  NOR3_X1 U257 ( .A1(n98), .A2(n99), .A3(n100), .ZN(n305) );
  XOR2_X1 U258 ( .A(Instr_reg_out[18]), .B(RD1[2]), .Z(n98) );
  XOR2_X1 U259 ( .A(Instr_reg_out[16]), .B(RD1[0]), .Z(n99) );
  XOR2_X1 U260 ( .A(Instr_reg_out[17]), .B(RD1[1]), .Z(n100) );
  INV_X1 U261 ( .A(Instr_reg_out[26]), .ZN(n229) );
  INV_X1 U262 ( .A(ALU_reg_out[0]), .ZN(n206) );
  INV_X1 U263 ( .A(ALU_reg_out[6]), .ZN(n122) );
  INV_X1 U264 ( .A(ALU_reg_out[10]), .ZN(n203) );
  INV_X1 U265 ( .A(ALU_reg_out[11]), .ZN(n200) );
  INV_X1 U266 ( .A(ALU_reg_out[5]), .ZN(n125) );
  AND3_X1 U267 ( .A1(n282), .A2(n283), .A3(Instr[27]), .ZN(n281) );
  INV_X1 U268 ( .A(Instr_reg_out[27]), .ZN(n280) );
  AND4_X1 U269 ( .A1(LOAD_op1), .A2(n305), .A3(n306), .A4(n307), .ZN(
        FWD_B_mem_mem) );
  AND2_X1 U270 ( .A1(n281), .A2(Instr[30]), .ZN(JR_op) );
  INV_X1 U271 ( .A(Instr_reg_out[31]), .ZN(n278) );
  NAND2_X1 U272 ( .A1(RF_out_A[23]), .A2(n430), .ZN(n163) );
  NAND2_X1 U273 ( .A1(RF_out_A[21]), .A2(n430), .ZN(n169) );
  NAND2_X1 U274 ( .A1(RF_out_A[18]), .A2(n429), .ZN(n181) );
  NAND2_X1 U275 ( .A1(RF_out_A[16]), .A2(n429), .ZN(n187) );
  NAND2_X1 U276 ( .A1(RF_out_A[15]), .A2(n429), .ZN(n190) );
  NAND2_X1 U277 ( .A1(RF_out_A[14]), .A2(n429), .ZN(n193) );
  NAND2_X1 U278 ( .A1(RF_out_A[13]), .A2(n429), .ZN(n196) );
  NAND2_X1 U279 ( .A1(RF_out_A[12]), .A2(n429), .ZN(n199) );
  NAND2_X1 U280 ( .A1(RF_out_A[11]), .A2(n429), .ZN(n202) );
  NAND2_X1 U281 ( .A1(RF_out_A[10]), .A2(n429), .ZN(n205) );
  NAND2_X1 U282 ( .A1(RF_out_A[1]), .A2(n429), .ZN(n175) );
  NAND2_X1 U283 ( .A1(RF_out_A[0]), .A2(n429), .ZN(n208) );
  NAND2_X1 U284 ( .A1(RF_out_A[28]), .A2(n430), .ZN(n148) );
  NAND2_X1 U285 ( .A1(RF_out_A[26]), .A2(n430), .ZN(n154) );
  NAND2_X1 U286 ( .A1(RF_out_A[24]), .A2(n430), .ZN(n160) );
  NAND2_X1 U287 ( .A1(RF_out_A[22]), .A2(n430), .ZN(n166) );
  NAND2_X1 U288 ( .A1(RF_out_A[20]), .A2(n430), .ZN(n172) );
  NAND2_X1 U289 ( .A1(RF_out_A[19]), .A2(n429), .ZN(n178) );
  NAND2_X1 U290 ( .A1(RF_out_A[17]), .A2(n429), .ZN(n184) );
  NAND2_X1 U291 ( .A1(RF_out_A[2]), .A2(n430), .ZN(n142) );
  NAND2_X1 U292 ( .A1(RF_out_A[27]), .A2(n430), .ZN(n151) );
  NAND2_X1 U293 ( .A1(RF_out_A[25]), .A2(n430), .ZN(n157) );
  NAND2_X1 U294 ( .A1(RF_out_A[30]), .A2(n430), .ZN(n139) );
  NAND2_X1 U295 ( .A1(RF_out_A[29]), .A2(n430), .ZN(n145) );
  NOR4_X1 U296 ( .A1(n283), .A2(n422), .A3(Instr[27]), .A4(Instr[30]), .ZN(
        BRANCH_op) );
  INV_X1 U297 ( .A(n282), .ZN(n422) );
  AND4_X1 U298 ( .A1(n200), .A2(n203), .A3(n206), .A4(FWD_exe_branch1), .ZN(
        n241) );
  INV_X1 U299 ( .A(Instr[28]), .ZN(n283) );
  AND4_X1 U300 ( .A1(n315), .A2(n316), .A3(n317), .A4(n318), .ZN(FWD_B_exe_mem) );
  NOR3_X1 U301 ( .A1(OPCODE1[0]), .A2(OPCODE1[2]), .A3(OPCODE1[1]), .ZN(n317)
         );
  NOR3_X1 U302 ( .A1(OPCODE1[3]), .A2(OPCODE1[5]), .A3(OPCODE1[4]), .ZN(n318)
         );
  AND4_X1 U303 ( .A1(n285), .A2(n286), .A3(n287), .A4(n288), .ZN(FWD_B_wb_mem)
         );
  NOR3_X1 U304 ( .A1(OPCODE2[0]), .A2(OPCODE2[2]), .A3(OPCODE2[1]), .ZN(n287)
         );
  NOR3_X1 U305 ( .A1(OPCODE2[3]), .A2(OPCODE2[5]), .A3(OPCODE2[4]), .ZN(n288)
         );
  NOR4_X1 U306 ( .A1(RD1[3]), .A2(RD1[4]), .A3(RD1[2]), .A4(n343), .ZN(n320)
         );
  OR2_X1 U307 ( .A1(RD1[1]), .A2(RD1[0]), .ZN(n343) );
  NAND2_X1 U308 ( .A1(n266), .A2(n267), .ZN(PC_Immediate_displacement[31]) );
  NAND2_X1 U309 ( .A1(JUMP_EN), .A2(Instr[25]), .ZN(n267) );
  BUF_X2 U310 ( .A(n39), .Z(n452) );
  XNOR2_X1 U311 ( .A(Instr_reg_out[20]), .B(RD2[4]), .ZN(n302) );
  XNOR2_X1 U312 ( .A(Instr_reg_out[19]), .B(RD2[3]), .ZN(n300) );
  NAND4_X1 U313 ( .A1(LOAD_op2), .A2(n301), .A3(n300), .A4(n302), .ZN(n308) );
  OR2_X1 U314 ( .A1(forward_branch), .A2(JUMP_EN), .ZN(n266) );
  OR2_X1 U315 ( .A1(PC_enable1), .A2(bootstrap), .ZN(PC_enable_fixed) );
  BUF_X1 U316 ( .A(n39), .Z(n453) );
  NOR3_X1 U317 ( .A1(n101), .A2(n102), .A3(n113), .ZN(n301) );
  XOR2_X1 U318 ( .A(Instr_reg_out[18]), .B(RD2[2]), .Z(n101) );
  XOR2_X1 U319 ( .A(Instr_reg_out[16]), .B(RD2[0]), .Z(n102) );
  XOR2_X1 U320 ( .A(Instr_reg_out[17]), .B(RD2[1]), .Z(n113) );
  OR3_X1 U321 ( .A1(STORE_op1), .A2(LOAD_op1), .A3(n320), .ZN(n328) );
  INV_X1 U322 ( .A(BRANCH_op1), .ZN(n284) );
  INV_X1 U323 ( .A(LOAD_op2), .ZN(n335) );
  INV_X1 U324 ( .A(ALU_reg_out[9]), .ZN(n111) );
  INV_X1 U325 ( .A(ALU_reg_out[1]), .ZN(n173) );
  INV_X1 U326 ( .A(ALU_reg_out[8]), .ZN(n116) );
  INV_X1 U327 ( .A(ALU_reg_out[7]), .ZN(n119) );
  INV_X1 U328 ( .A(ALU_reg_out[3]), .ZN(n131) );
  INV_X1 U329 ( .A(ALU_reg_out[4]), .ZN(n128) );
  INV_X1 U330 ( .A(ALU_reg_out[2]), .ZN(n140) );
  INV_X1 U331 ( .A(ALU_reg_out[23]), .ZN(n161) );
  INV_X1 U332 ( .A(ALU_reg_out[16]), .ZN(n185) );
  INV_X1 U333 ( .A(ALU_reg_out[12]), .ZN(n197) );
  INV_X1 U334 ( .A(ALU_reg_out[27]), .ZN(n149) );
  INV_X1 U335 ( .A(ALU_reg_out[30]), .ZN(n137) );
  INV_X1 U336 ( .A(ALU_reg_out[13]), .ZN(n194) );
  INV_X1 U337 ( .A(ALU_reg_out[28]), .ZN(n146) );
  INV_X1 U338 ( .A(ALU_reg_out[24]), .ZN(n158) );
  INV_X1 U339 ( .A(ALU_reg_out[20]), .ZN(n170) );
  INV_X1 U340 ( .A(ALU_reg_out[17]), .ZN(n182) );
  INV_X1 U341 ( .A(ALU_reg_out[31]), .ZN(n134) );
  INV_X1 U342 ( .A(ALU_reg_out[21]), .ZN(n167) );
  INV_X1 U343 ( .A(ALU_reg_out[18]), .ZN(n179) );
  INV_X1 U344 ( .A(ALU_reg_out[14]), .ZN(n191) );
  INV_X1 U345 ( .A(ALU_reg_out[25]), .ZN(n155) );
  INV_X1 U346 ( .A(ALU_reg_out[29]), .ZN(n143) );
  INV_X1 U347 ( .A(ALU_reg_out[15]), .ZN(n188) );
  INV_X1 U348 ( .A(ALU_reg_out[26]), .ZN(n152) );
  INV_X1 U349 ( .A(ALU_reg_out[22]), .ZN(n164) );
  INV_X1 U350 ( .A(ALU_reg_out[19]), .ZN(n176) );
  NAND2_X1 U351 ( .A1(n266), .A2(n268), .ZN(PC_Immediate_displacement[24]) );
  NAND2_X1 U352 ( .A1(Instr[24]), .A2(JUMP_EN), .ZN(n268) );
  NAND2_X1 U353 ( .A1(n266), .A2(n269), .ZN(PC_Immediate_displacement[23]) );
  NAND2_X1 U354 ( .A1(Instr[23]), .A2(JUMP_EN), .ZN(n269) );
  NAND2_X1 U355 ( .A1(n266), .A2(n270), .ZN(PC_Immediate_displacement[22]) );
  NAND2_X1 U356 ( .A1(Instr[22]), .A2(JUMP_EN), .ZN(n270) );
  NAND2_X1 U357 ( .A1(n266), .A2(n271), .ZN(PC_Immediate_displacement[21]) );
  NAND2_X1 U358 ( .A1(Instr[21]), .A2(JUMP_EN), .ZN(n271) );
  NAND2_X1 U359 ( .A1(n266), .A2(n272), .ZN(PC_Immediate_displacement[20]) );
  NAND2_X1 U360 ( .A1(Instr[20]), .A2(JUMP_EN), .ZN(n272) );
  NAND2_X1 U361 ( .A1(n266), .A2(n273), .ZN(PC_Immediate_displacement[19]) );
  NAND2_X1 U362 ( .A1(Instr[19]), .A2(JUMP_EN), .ZN(n273) );
  NAND2_X1 U363 ( .A1(n266), .A2(n274), .ZN(PC_Immediate_displacement[18]) );
  NAND2_X1 U364 ( .A1(Instr[18]), .A2(JUMP_EN), .ZN(n274) );
  NAND2_X1 U365 ( .A1(n266), .A2(n275), .ZN(PC_Immediate_displacement[17]) );
  NAND2_X1 U366 ( .A1(Instr[17]), .A2(JUMP_EN), .ZN(n275) );
  NAND2_X1 U367 ( .A1(n266), .A2(n276), .ZN(PC_Immediate_displacement[16]) );
  NAND2_X1 U368 ( .A1(Instr[16]), .A2(JUMP_EN), .ZN(n276) );
  INV_X1 U369 ( .A(flush2[1]), .ZN(n298) );
  INV_X1 U370 ( .A(flush2[0]), .ZN(n297) );
  INV_X1 U371 ( .A(STORE_op2), .ZN(n299) );
  INV_X1 U372 ( .A(Instr[15]), .ZN(forward_branch) );
  OR2_X1 U373 ( .A1(RD2[1]), .A2(RD2[0]), .ZN(n342) );
  NOR4_X1 U374 ( .A1(Instr_reg_out[30]), .A2(Instr_reg_out[29]), .A3(n277), 
        .A4(n278), .ZN(LOAD_op) );
  AOI21_X1 U375 ( .B1(Instr_reg_out[26]), .B2(n279), .A(n280), .ZN(n277) );
  NOR4_X1 U376 ( .A1(JUMP_EN2), .A2(BRANCH_op1), .A3(n230), .A4(n328), .ZN(
        FWD_A_exe_dec) );
  NOR4_X1 U377 ( .A1(n333), .A2(n334), .A3(n290), .A4(n212), .ZN(FWD_A_wb_dec)
         );
  OR2_X1 U378 ( .A1(BRANCH_op1), .A2(JUMP_EN2), .ZN(n334) );
  NAND4_X1 U379 ( .A1(n335), .A2(n299), .A3(n297), .A4(n298), .ZN(n333) );
  NOR3_X1 U380 ( .A1(n308), .A2(n290), .A3(n309), .ZN(FWD_B_mem_exe) );
  NOR4_X1 U381 ( .A1(Instr_reg_out[30]), .A2(n310), .A3(n311), .A4(n279), .ZN(
        n309) );
  INV_X1 U382 ( .A(Instr_reg_out[29]), .ZN(n310) );
  NOR4_X1 U383 ( .A1(n295), .A2(n296), .A3(LOAD_op2), .A4(n290), .ZN(
        FWD_B_wb_dec) );
  NAND4_X1 U384 ( .A1(n300), .A2(n301), .A3(n302), .A4(n303), .ZN(n295) );
  AND2_X1 U385 ( .A1(Instr[26]), .A2(n281), .ZN(JAL_op) );
  NOR3_X1 U386 ( .A1(FWD_B_lmd1_mem2), .A2(FWD_B_mem_mem2), .A3(n418), .ZN(
        n354) );
  BUF_X1 U387 ( .A(FWD_B_exe_mem2), .Z(n439) );
  NOR2_X1 U388 ( .A1(n421), .A2(n439), .ZN(n352) );
  INV_X1 U389 ( .A(FWD_B_wb_mem2), .ZN(n421) );
  BUF_X1 U390 ( .A(FWD_B_exe_mem2), .Z(n438) );
  BUF_X1 U391 ( .A(FWD_B_exe_mem2), .Z(n437) );
  NOR2_X1 U392 ( .A1(n439), .A2(FWD_B_wb_mem2), .ZN(n419) );
  AND3_X1 U393 ( .A1(n419), .A2(n420), .A3(FWD_B_lmd1_mem2), .ZN(n353) );
  INV_X1 U394 ( .A(FWD_B_mem_mem2), .ZN(n420) );
  NAND2_X1 U395 ( .A1(n366), .A2(n367), .ZN(DRAM_write_data_FWD[3]) );
  AOI22_X1 U396 ( .A1(LMD_reg_out[3]), .A2(n313), .B1(ALU_WB_out[3]), .B2(n437), .ZN(n366) );
  AOI222_X1 U397 ( .A1(ALU_WB_out1[3]), .A2(n428), .B1(LMD_reg_out1[3]), .B2(
        n425), .C1(DRAM_write_data[3]), .C2(n331), .ZN(n367) );
  NAND2_X1 U398 ( .A1(n364), .A2(n365), .ZN(DRAM_write_data_FWD[4]) );
  AOI22_X1 U399 ( .A1(LMD_reg_out[4]), .A2(n313), .B1(ALU_WB_out[4]), .B2(n437), .ZN(n364) );
  AOI222_X1 U400 ( .A1(ALU_WB_out1[4]), .A2(n428), .B1(LMD_reg_out1[4]), .B2(
        n425), .C1(DRAM_write_data[4]), .C2(n331), .ZN(n365) );
  NAND2_X1 U401 ( .A1(n362), .A2(n363), .ZN(DRAM_write_data_FWD[5]) );
  AOI22_X1 U402 ( .A1(LMD_reg_out[5]), .A2(n313), .B1(ALU_WB_out[5]), .B2(n437), .ZN(n362) );
  AOI222_X1 U403 ( .A1(ALU_WB_out1[5]), .A2(n428), .B1(LMD_reg_out1[5]), .B2(
        n425), .C1(DRAM_write_data[5]), .C2(n331), .ZN(n363) );
  NAND2_X1 U404 ( .A1(n360), .A2(n361), .ZN(DRAM_write_data_FWD[6]) );
  AOI22_X1 U405 ( .A1(LMD_reg_out[6]), .A2(n313), .B1(ALU_WB_out[6]), .B2(n437), .ZN(n360) );
  AOI222_X1 U406 ( .A1(ALU_WB_out1[6]), .A2(n428), .B1(LMD_reg_out1[6]), .B2(
        n425), .C1(DRAM_write_data[6]), .C2(n331), .ZN(n361) );
  NAND2_X1 U407 ( .A1(n358), .A2(n359), .ZN(DRAM_write_data_FWD[7]) );
  AOI22_X1 U408 ( .A1(LMD_reg_out[7]), .A2(n313), .B1(ALU_WB_out[7]), .B2(n437), .ZN(n358) );
  AOI222_X1 U409 ( .A1(ALU_WB_out1[7]), .A2(n428), .B1(LMD_reg_out1[7]), .B2(
        n425), .C1(DRAM_write_data[7]), .C2(n331), .ZN(n359) );
  NAND2_X1 U410 ( .A1(n356), .A2(n357), .ZN(DRAM_write_data_FWD[8]) );
  AOI22_X1 U411 ( .A1(LMD_reg_out[8]), .A2(n313), .B1(ALU_WB_out[8]), .B2(n437), .ZN(n356) );
  AOI222_X1 U412 ( .A1(ALU_WB_out1[8]), .A2(n428), .B1(LMD_reg_out1[8]), .B2(
        n425), .C1(DRAM_write_data[8]), .C2(n331), .ZN(n357) );
  NAND2_X1 U413 ( .A1(n350), .A2(n351), .ZN(DRAM_write_data_FWD[9]) );
  AOI22_X1 U414 ( .A1(LMD_reg_out[9]), .A2(n313), .B1(n439), .B2(ALU_WB_out[9]), .ZN(n350) );
  AOI222_X1 U415 ( .A1(ALU_WB_out1[9]), .A2(n428), .B1(LMD_reg_out1[9]), .B2(
        n425), .C1(DRAM_write_data[9]), .C2(n331), .ZN(n351) );
  NAND2_X1 U416 ( .A1(n368), .A2(n369), .ZN(DRAM_write_data_FWD[31]) );
  AOI22_X1 U417 ( .A1(LMD_reg_out[31]), .A2(n313), .B1(ALU_WB_out[31]), .B2(
        n437), .ZN(n368) );
  AOI222_X1 U418 ( .A1(ALU_WB_out1[31]), .A2(n428), .B1(LMD_reg_out1[31]), 
        .B2(n425), .C1(DRAM_write_data[31]), .C2(n331), .ZN(n369) );
  NAND2_X1 U419 ( .A1(n416), .A2(n417), .ZN(DRAM_write_data_FWD[0]) );
  AOI22_X1 U420 ( .A1(LMD_reg_out[0]), .A2(n210), .B1(ALU_WB_out[0]), .B2(n439), .ZN(n416) );
  AOI222_X1 U421 ( .A1(ALU_WB_out1[0]), .A2(n426), .B1(LMD_reg_out1[0]), .B2(
        n332), .C1(DRAM_write_data[0]), .C2(n314), .ZN(n417) );
  NAND2_X1 U422 ( .A1(n394), .A2(n395), .ZN(DRAM_write_data_FWD[1]) );
  AOI22_X1 U423 ( .A1(LMD_reg_out[1]), .A2(n210), .B1(ALU_WB_out[1]), .B2(n438), .ZN(n394) );
  AOI222_X1 U424 ( .A1(ALU_WB_out1[1]), .A2(n426), .B1(LMD_reg_out1[1]), .B2(
        n332), .C1(DRAM_write_data[1]), .C2(n314), .ZN(n395) );
  NAND2_X1 U425 ( .A1(n372), .A2(n373), .ZN(DRAM_write_data_FWD[2]) );
  AOI22_X1 U426 ( .A1(LMD_reg_out[2]), .A2(n312), .B1(ALU_WB_out[2]), .B2(n437), .ZN(n372) );
  AOI222_X1 U427 ( .A1(ALU_WB_out1[2]), .A2(n427), .B1(LMD_reg_out1[2]), .B2(
        n424), .C1(DRAM_write_data[2]), .C2(n330), .ZN(n373) );
  NAND2_X1 U428 ( .A1(n414), .A2(n415), .ZN(DRAM_write_data_FWD[10]) );
  AOI22_X1 U429 ( .A1(LMD_reg_out[10]), .A2(n210), .B1(ALU_WB_out[10]), .B2(
        n439), .ZN(n414) );
  AOI222_X1 U430 ( .A1(ALU_WB_out1[10]), .A2(n426), .B1(LMD_reg_out1[10]), 
        .B2(n332), .C1(DRAM_write_data[10]), .C2(n314), .ZN(n415) );
  NAND2_X1 U431 ( .A1(n412), .A2(n413), .ZN(DRAM_write_data_FWD[11]) );
  AOI22_X1 U432 ( .A1(LMD_reg_out[11]), .A2(n210), .B1(ALU_WB_out[11]), .B2(
        n439), .ZN(n412) );
  AOI222_X1 U433 ( .A1(ALU_WB_out1[11]), .A2(n426), .B1(LMD_reg_out1[11]), 
        .B2(n332), .C1(DRAM_write_data[11]), .C2(n314), .ZN(n413) );
  NAND2_X1 U434 ( .A1(n410), .A2(n411), .ZN(DRAM_write_data_FWD[12]) );
  AOI22_X1 U435 ( .A1(LMD_reg_out[12]), .A2(n210), .B1(ALU_WB_out[12]), .B2(
        n439), .ZN(n410) );
  AOI222_X1 U436 ( .A1(ALU_WB_out1[12]), .A2(n426), .B1(LMD_reg_out1[12]), 
        .B2(n332), .C1(DRAM_write_data[12]), .C2(n314), .ZN(n411) );
  NAND2_X1 U437 ( .A1(n408), .A2(n409), .ZN(DRAM_write_data_FWD[13]) );
  AOI22_X1 U438 ( .A1(LMD_reg_out[13]), .A2(n210), .B1(ALU_WB_out[13]), .B2(
        n439), .ZN(n408) );
  AOI222_X1 U439 ( .A1(ALU_WB_out1[13]), .A2(n426), .B1(LMD_reg_out1[13]), 
        .B2(n332), .C1(DRAM_write_data[13]), .C2(n314), .ZN(n409) );
  NAND2_X1 U440 ( .A1(n406), .A2(n407), .ZN(DRAM_write_data_FWD[14]) );
  AOI22_X1 U441 ( .A1(LMD_reg_out[14]), .A2(n210), .B1(ALU_WB_out[14]), .B2(
        n439), .ZN(n406) );
  AOI222_X1 U442 ( .A1(ALU_WB_out1[14]), .A2(n426), .B1(LMD_reg_out1[14]), 
        .B2(n332), .C1(DRAM_write_data[14]), .C2(n314), .ZN(n407) );
  NAND2_X1 U443 ( .A1(n404), .A2(n405), .ZN(DRAM_write_data_FWD[15]) );
  AOI22_X1 U444 ( .A1(LMD_reg_out[15]), .A2(n210), .B1(ALU_WB_out[15]), .B2(
        n439), .ZN(n404) );
  AOI222_X1 U445 ( .A1(ALU_WB_out1[15]), .A2(n426), .B1(LMD_reg_out1[15]), 
        .B2(n332), .C1(DRAM_write_data[15]), .C2(n314), .ZN(n405) );
  NAND2_X1 U446 ( .A1(n402), .A2(n403), .ZN(DRAM_write_data_FWD[16]) );
  AOI22_X1 U447 ( .A1(LMD_reg_out[16]), .A2(n210), .B1(ALU_WB_out[16]), .B2(
        n438), .ZN(n402) );
  AOI222_X1 U448 ( .A1(ALU_WB_out1[16]), .A2(n426), .B1(LMD_reg_out1[16]), 
        .B2(n332), .C1(DRAM_write_data[16]), .C2(n314), .ZN(n403) );
  NAND2_X1 U449 ( .A1(n400), .A2(n401), .ZN(DRAM_write_data_FWD[17]) );
  AOI22_X1 U450 ( .A1(LMD_reg_out[17]), .A2(n210), .B1(ALU_WB_out[17]), .B2(
        n438), .ZN(n400) );
  AOI222_X1 U451 ( .A1(ALU_WB_out1[17]), .A2(n426), .B1(LMD_reg_out1[17]), 
        .B2(n332), .C1(DRAM_write_data[17]), .C2(n314), .ZN(n401) );
  NAND2_X1 U452 ( .A1(n398), .A2(n399), .ZN(DRAM_write_data_FWD[18]) );
  AOI22_X1 U453 ( .A1(LMD_reg_out[18]), .A2(n210), .B1(ALU_WB_out[18]), .B2(
        n438), .ZN(n398) );
  AOI222_X1 U454 ( .A1(ALU_WB_out1[18]), .A2(n426), .B1(LMD_reg_out1[18]), 
        .B2(n332), .C1(DRAM_write_data[18]), .C2(n314), .ZN(n399) );
  NAND2_X1 U455 ( .A1(n396), .A2(n397), .ZN(DRAM_write_data_FWD[19]) );
  AOI22_X1 U465 ( .A1(LMD_reg_out[19]), .A2(n210), .B1(ALU_WB_out[19]), .B2(
        n438), .ZN(n396) );
  AOI222_X1 U466 ( .A1(ALU_WB_out1[19]), .A2(n426), .B1(LMD_reg_out1[19]), 
        .B2(n332), .C1(DRAM_write_data[19]), .C2(n314), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n392), .A2(n393), .ZN(DRAM_write_data_FWD[20]) );
  AOI22_X1 U468 ( .A1(LMD_reg_out[20]), .A2(n312), .B1(ALU_WB_out[20]), .B2(
        n438), .ZN(n392) );
  AOI222_X1 U469 ( .A1(ALU_WB_out1[20]), .A2(n427), .B1(LMD_reg_out1[20]), 
        .B2(n424), .C1(DRAM_write_data[20]), .C2(n330), .ZN(n393) );
  NAND2_X1 U470 ( .A1(n390), .A2(n391), .ZN(DRAM_write_data_FWD[21]) );
  AOI22_X1 U471 ( .A1(LMD_reg_out[21]), .A2(n312), .B1(ALU_WB_out[21]), .B2(
        n438), .ZN(n390) );
  AOI222_X1 U472 ( .A1(ALU_WB_out1[21]), .A2(n427), .B1(LMD_reg_out1[21]), 
        .B2(n424), .C1(DRAM_write_data[21]), .C2(n330), .ZN(n391) );
  NAND2_X1 U473 ( .A1(n388), .A2(n389), .ZN(DRAM_write_data_FWD[22]) );
  AOI22_X1 U474 ( .A1(LMD_reg_out[22]), .A2(n312), .B1(ALU_WB_out[22]), .B2(
        n438), .ZN(n388) );
  AOI222_X1 U475 ( .A1(ALU_WB_out1[22]), .A2(n427), .B1(LMD_reg_out1[22]), 
        .B2(n424), .C1(DRAM_write_data[22]), .C2(n330), .ZN(n389) );
  NAND2_X1 U476 ( .A1(n386), .A2(n387), .ZN(DRAM_write_data_FWD[23]) );
  AOI22_X1 U477 ( .A1(LMD_reg_out[23]), .A2(n312), .B1(ALU_WB_out[23]), .B2(
        n438), .ZN(n386) );
  AOI222_X1 U478 ( .A1(ALU_WB_out1[23]), .A2(n427), .B1(LMD_reg_out1[23]), 
        .B2(n424), .C1(DRAM_write_data[23]), .C2(n330), .ZN(n387) );
  NAND2_X1 U479 ( .A1(n384), .A2(n385), .ZN(DRAM_write_data_FWD[24]) );
  AOI22_X1 U480 ( .A1(LMD_reg_out[24]), .A2(n312), .B1(ALU_WB_out[24]), .B2(
        n438), .ZN(n384) );
  AOI222_X1 U481 ( .A1(ALU_WB_out1[24]), .A2(n427), .B1(LMD_reg_out1[24]), 
        .B2(n424), .C1(DRAM_write_data[24]), .C2(n330), .ZN(n385) );
  NAND2_X1 U482 ( .A1(n382), .A2(n383), .ZN(DRAM_write_data_FWD[25]) );
  AOI22_X1 U483 ( .A1(LMD_reg_out[25]), .A2(n312), .B1(ALU_WB_out[25]), .B2(
        n438), .ZN(n382) );
  AOI222_X1 U484 ( .A1(ALU_WB_out1[25]), .A2(n427), .B1(LMD_reg_out1[25]), 
        .B2(n424), .C1(DRAM_write_data[25]), .C2(n330), .ZN(n383) );
  NAND2_X1 U485 ( .A1(n380), .A2(n381), .ZN(DRAM_write_data_FWD[26]) );
  AOI22_X1 U486 ( .A1(LMD_reg_out[26]), .A2(n312), .B1(ALU_WB_out[26]), .B2(
        n437), .ZN(n380) );
  AOI222_X1 U487 ( .A1(ALU_WB_out1[26]), .A2(n427), .B1(LMD_reg_out1[26]), 
        .B2(n424), .C1(DRAM_write_data[26]), .C2(n330), .ZN(n381) );
  NAND2_X1 U488 ( .A1(n378), .A2(n379), .ZN(DRAM_write_data_FWD[27]) );
  AOI22_X1 U489 ( .A1(LMD_reg_out[27]), .A2(n312), .B1(ALU_WB_out[27]), .B2(
        n437), .ZN(n378) );
  AOI222_X1 U490 ( .A1(ALU_WB_out1[27]), .A2(n427), .B1(LMD_reg_out1[27]), 
        .B2(n424), .C1(DRAM_write_data[27]), .C2(n330), .ZN(n379) );
  NAND2_X1 U491 ( .A1(n376), .A2(n377), .ZN(DRAM_write_data_FWD[28]) );
  AOI22_X1 U492 ( .A1(LMD_reg_out[28]), .A2(n312), .B1(ALU_WB_out[28]), .B2(
        n437), .ZN(n376) );
  AOI222_X1 U493 ( .A1(ALU_WB_out1[28]), .A2(n427), .B1(LMD_reg_out1[28]), 
        .B2(n424), .C1(DRAM_write_data[28]), .C2(n330), .ZN(n377) );
  NAND2_X1 U494 ( .A1(n374), .A2(n375), .ZN(DRAM_write_data_FWD[29]) );
  AOI22_X1 U495 ( .A1(LMD_reg_out[29]), .A2(n312), .B1(ALU_WB_out[29]), .B2(
        n437), .ZN(n374) );
  AOI222_X1 U496 ( .A1(ALU_WB_out1[29]), .A2(n427), .B1(LMD_reg_out1[29]), 
        .B2(n424), .C1(DRAM_write_data[29]), .C2(n330), .ZN(n375) );
  NAND2_X1 U497 ( .A1(n370), .A2(n371), .ZN(DRAM_write_data_FWD[30]) );
  AOI22_X1 U498 ( .A1(LMD_reg_out[30]), .A2(n312), .B1(ALU_WB_out[30]), .B2(
        n438), .ZN(n370) );
  AOI222_X1 U499 ( .A1(ALU_WB_out1[30]), .A2(n427), .B1(LMD_reg_out1[30]), 
        .B2(n424), .C1(DRAM_write_data[30]), .C2(n330), .ZN(n371) );
endmodule


module dlx ( Clk, Rst, IR, PC );
  input [31:0] IR;
  output [31:0] PC;
  input Clk, Rst;

  wire   [4:0] ALU_OPCODE;
  wire   [1:0] flush;

  datapath DTP ( .Clk(Clk), .Rst(Rst), .Instr(IR), .JUMP_EN(1'b0), .RF_RD1_EN(
        1'b0), .RF_RD2_EN(1'b0), .RF_EN(1'b0), .CALL(1'b0), .RET(1'b0), 
        .IMM_SEL(1'b0), .MUXA_SEL(1'b0), .MUXB_SEL(1'b0), .EQ_COND(1'b0), 
        .ALU_OPCODE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_STORE1(1'b0), 
        .SEL_STORE0(1'b0), .SEL_LOAD2(1'b0), .SEL_LOAD1(1'b0), .SEL_LOAD0(1'b0), .DRAM_WR(1'b0), .WB_MUX_SEL(1'b0), .RF_WR(1'b0), .flush(flush), .PC_out(PC)
         );
  CU_HW CTRLU ( .Clk(Clk), .Rst(Rst), .IR_IN(IR), .flush(flush) );
endmodule

