
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_alu is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
subtype bus32 is std_logic_vector (31 downto 0);
type aluOp is (NOP, ADDOP, SUBOP, MULOP, ANDOP, OROP, XOROP, SLLOP, SRLOP, 
   SRAOP, GTOP, GETOP, LTOP, LETOP, EQOP, NEQOP, GTUOP, GETUOP, LTUOP, LETUOP, 
   LHIOP);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_alu;

package body CONV_PACK_alu is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when ADDOP => return "00001";
         when SUBOP => return "00010";
         when MULOP => return "00011";
         when ANDOP => return "00100";
         when OROP => return "00101";
         when XOROP => return "00110";
         when SLLOP => return "00111";
         when SRLOP => return "01000";
         when SRAOP => return "01001";
         when GTOP => return "01010";
         when GETOP => return "01011";
         when LTOP => return "01100";
         when LETOP => return "01101";
         when EQOP => return "01110";
         when NEQOP => return "01111";
         when GTUOP => return "10000";
         when GETUOP => return "10001";
         when LTUOP => return "10010";
         when LETUOP => return "10011";
         when LHIOP => return "10100";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_alu;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n17, n18 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n18, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n18);
   U1 : INV_X1 port map( A => n17, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n18, B2 => Ci, ZN => n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_23;

architecture SYN_STRUCTURAL of rca_generic_N4_23 is

   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_287 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_286 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_285 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_284 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_22;

architecture SYN_STRUCTURAL of rca_generic_N4_22 is

   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_283 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_282 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_281 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_280 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_9;

architecture SYN_STRUCTURAL of rca_generic_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_8;

architecture SYN_STRUCTURAL of rca_generic_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_7;

architecture SYN_STRUCTURAL of rca_generic_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_27;

architecture SYN_STRUCTURAL of rca_generic_N4_27 is

   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_303 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_302 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_301 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_300 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_26;

architecture SYN_STRUCTURAL of rca_generic_N4_26 is

   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_299 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_298 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_297 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_296 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_25;

architecture SYN_STRUCTURAL of rca_generic_N4_25 is

   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_295 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_294 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_293 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_292 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_21;

architecture SYN_STRUCTURAL of rca_generic_N4_21 is

   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_279 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_278 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_277 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_276 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_20;

architecture SYN_STRUCTURAL of rca_generic_N4_20 is

   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_275 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_274 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_273 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_272 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_13;

architecture SYN_STRUCTURAL of rca_generic_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_12;

architecture SYN_STRUCTURAL of rca_generic_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_11;

architecture SYN_STRUCTURAL of rca_generic_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_10;

architecture SYN_STRUCTURAL of rca_generic_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_6;

architecture SYN_STRUCTURAL of rca_generic_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_5;

architecture SYN_STRUCTURAL of rca_generic_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_4;

architecture SYN_STRUCTURAL of rca_generic_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_3;

architecture SYN_STRUCTURAL of rca_generic_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_2;

architecture SYN_STRUCTURAL of rca_generic_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_1;

architecture SYN_STRUCTURAL of rca_generic_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_35 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_35;

architecture SYN_STRUCTURAL of PG_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_17 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_17;

architecture SYN_STRUCTURAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_16 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_16;

architecture SYN_STRUCTURAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n10);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_32 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_32;

architecture SYN_STRUCTURAL of PG_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_20 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_20;

architecture SYN_STRUCTURAL of PG_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n9, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_6 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_6;

architecture SYN_STRUCTURAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_43 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_43;

architecture SYN_STRUCTURAL of PG_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_41 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_41;

architecture SYN_STRUCTURAL of PG_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_40 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_40;

architecture SYN_STRUCTURAL of PG_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_39 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_39;

architecture SYN_STRUCTURAL of PG_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_38 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_38;

architecture SYN_STRUCTURAL of PG_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_31 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_31;

architecture SYN_STRUCTURAL of PG_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_29 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_29;

architecture SYN_STRUCTURAL of PG_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_27 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_27;

architecture SYN_STRUCTURAL of PG_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_12 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_12;

architecture SYN_STRUCTURAL of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_11 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_11;

architecture SYN_STRUCTURAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_10 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_10;

architecture SYN_STRUCTURAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_9 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_9;

architecture SYN_STRUCTURAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_8 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_8;

architecture SYN_STRUCTURAL of PG_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_7 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_7;

architecture SYN_STRUCTURAL of PG_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_5 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_5;

architecture SYN_STRUCTURAL of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_3 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_3;

architecture SYN_STRUCTURAL of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_2 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_2;

architecture SYN_STRUCTURAL of PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_11 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_11;

architecture SYN_STRUCTURAL of G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_2 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_2;

architecture SYN_STRUCTURAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_4 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_4;

architecture SYN_STRUCTURAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_12 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_12;

architecture SYN_STRUCTURAL of G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_10 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_10;

architecture SYN_STRUCTURAL of G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_9 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_9;

architecture SYN_STRUCTURAL of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_7 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_7;

architecture SYN_STRUCTURAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_3 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_3;

architecture SYN_STRUCTURAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_59 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_59;

architecture SYN_STRUCTURAL of PGnet_block_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_58 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_58;

architecture SYN_STRUCTURAL of PGnet_block_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_57 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_57;

architecture SYN_STRUCTURAL of PGnet_block_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_56 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_56;

architecture SYN_STRUCTURAL of PGnet_block_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_55 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_55;

architecture SYN_STRUCTURAL of PGnet_block_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_54 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_54;

architecture SYN_STRUCTURAL of PGnet_block_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_53 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_53;

architecture SYN_STRUCTURAL of PGnet_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_52 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_52;

architecture SYN_STRUCTURAL of PGnet_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_51 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_51;

architecture SYN_STRUCTURAL of PGnet_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_50 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_50;

architecture SYN_STRUCTURAL of PGnet_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_49 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_49;

architecture SYN_STRUCTURAL of PGnet_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_48 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_48;

architecture SYN_STRUCTURAL of PGnet_block_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_47 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_47;

architecture SYN_STRUCTURAL of PGnet_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_46 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_46;

architecture SYN_STRUCTURAL of PGnet_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_45 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_45;

architecture SYN_STRUCTURAL of PGnet_block_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_44 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_44;

architecture SYN_STRUCTURAL of PGnet_block_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_43 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_43;

architecture SYN_STRUCTURAL of PGnet_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_42 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_42;

architecture SYN_STRUCTURAL of PGnet_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_41 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_41;

architecture SYN_STRUCTURAL of PGnet_block_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_40 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_40;

architecture SYN_STRUCTURAL of PGnet_block_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_39 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_39;

architecture SYN_STRUCTURAL of PGnet_block_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_38 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_38;

architecture SYN_STRUCTURAL of PGnet_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_37 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_37;

architecture SYN_STRUCTURAL of PGnet_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_36 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_36;

architecture SYN_STRUCTURAL of PGnet_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_35 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_35;

architecture SYN_STRUCTURAL of PGnet_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_34 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_34;

architecture SYN_STRUCTURAL of PGnet_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_33 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_33;

architecture SYN_STRUCTURAL of PGnet_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_32 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_32;

architecture SYN_STRUCTURAL of PGnet_block_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_29 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_29;

architecture SYN_STRUCTURAL of PGnet_block_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_28 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_28;

architecture SYN_STRUCTURAL of PGnet_block_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_27 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_27;

architecture SYN_STRUCTURAL of PGnet_block_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_26 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_26;

architecture SYN_STRUCTURAL of PGnet_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_25 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_25;

architecture SYN_STRUCTURAL of PGnet_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_24 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_24;

architecture SYN_STRUCTURAL of PGnet_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_23 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_23;

architecture SYN_STRUCTURAL of PGnet_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_22 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_22;

architecture SYN_STRUCTURAL of PGnet_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_21 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_21;

architecture SYN_STRUCTURAL of PGnet_block_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_20 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_20;

architecture SYN_STRUCTURAL of PGnet_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_19 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_19;

architecture SYN_STRUCTURAL of PGnet_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_18 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_18;

architecture SYN_STRUCTURAL of PGnet_block_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_17 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_17;

architecture SYN_STRUCTURAL of PGnet_block_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_16 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_16;

architecture SYN_STRUCTURAL of PGnet_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_15 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_15;

architecture SYN_STRUCTURAL of PGnet_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_14 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_14;

architecture SYN_STRUCTURAL of PGnet_block_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_13 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_13;

architecture SYN_STRUCTURAL of PGnet_block_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_12 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_12;

architecture SYN_STRUCTURAL of PGnet_block_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_11 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_11;

architecture SYN_STRUCTURAL of PGnet_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_10 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_10;

architecture SYN_STRUCTURAL of PGnet_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_9 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_9;

architecture SYN_STRUCTURAL of PGnet_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_8 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_8;

architecture SYN_STRUCTURAL of PGnet_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_7 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_7;

architecture SYN_STRUCTURAL of PGnet_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_6 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_6;

architecture SYN_STRUCTURAL of PGnet_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_5 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_5;

architecture SYN_STRUCTURAL of PGnet_block_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_4 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_4;

architecture SYN_STRUCTURAL of PGnet_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_3 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_3;

architecture SYN_STRUCTURAL of PGnet_block_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_2 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_2;

architecture SYN_STRUCTURAL of PGnet_block_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_1;

architecture SYN_STRUCTURAL of PGnet_block_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH1 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH1 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH1 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH1 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH1 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH1 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH1 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH1 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH1 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH1 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH1 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH1 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH1 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH1 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH1 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH1 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH1 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH1 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH1 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH1 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH1 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH1 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH1 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH1 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH1 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH1 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH1 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH1 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH1 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH1 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH1 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH1 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH1 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH1 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH1 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH1 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH1 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH1 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH1 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH1 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH1 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH1 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH1 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH1 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH1 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH1 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH1 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH1 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH1 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH1 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH1 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH1 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH1 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH1 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH1 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH1 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH1 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH1 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH1 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH1 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH1 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH1 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH1 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH1 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH1 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH1 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH1 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH1 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH1 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH1 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH1 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH1 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH1 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH1 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH1 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH1 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH1 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH1 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH1 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH1 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH1 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH1 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH1 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH1 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH1 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH1 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH1 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH1 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH1 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH1 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH1 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH1 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH1 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH1 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH1 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH1 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH1 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH1 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH1 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH1 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH1 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH1 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH1 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH1 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH1 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH1 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH1 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH1 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH1 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH1 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH1 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH1 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH1 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH1 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH1 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH1 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH1 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH1 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH1 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH1 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH1 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH1 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH1 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH1 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH1 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH1 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH1 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH1 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH1 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH1 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH1 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH1 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH1 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH1 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH1 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH1 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH1 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH1 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH1 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH1 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH1 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH1 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH1 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH1 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH1 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH1 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH1 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH1 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH1 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH1 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH1 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH1 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH1 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH1 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH1 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH1 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH1 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH1 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH1 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH1 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH1 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH1 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH1 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH1 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH1 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH1 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH1 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH1 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH1 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH1 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH1 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH1 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH1 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH1 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH1 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH1 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH1 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH1 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH1 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH1 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH1 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH1 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH1 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH1 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH1 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_179 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_178 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_177 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_176 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_175 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_174 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_173 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_172 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_171 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_170 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_169 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_168 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_167 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_166 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_165 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_164 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_163 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_162 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_161 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_160 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_159 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_158 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_157 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_156 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_155 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_154 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_153 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_152 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_151 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_150 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_149 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_148 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_147 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_146 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_145 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_144 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_143 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_142 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_141 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_140 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_139 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_138 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_137 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_136 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_135 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_134 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_133 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_132 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_131 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_130 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_129 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_128 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_127 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_126 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_125 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_124 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_123 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_122 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_121 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_120 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_119 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_118 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_117 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_116 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_115 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_114 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_113 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_112 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_111 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_110 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_109 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_108 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_107 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_106 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_105 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_104 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_103 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_102 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_101 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_100 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_99 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_98 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_97 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_96 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_11;

architecture SYN_struct of MUX21_GENERIC_N4_11 is

   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_47 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_46 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_45 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_44 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_10;

architecture SYN_struct of MUX21_GENERIC_N4_10 is

   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_43 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_42 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_41 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_40 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_9;

architecture SYN_struct of MUX21_GENERIC_N4_9 is

   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_39 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_38 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_37 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_36 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_8;

architecture SYN_struct of MUX21_GENERIC_N4_8 is

   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_35 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_34 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_33 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_32 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_5;

architecture SYN_struct of MUX21_GENERIC_N4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_4;

architecture SYN_struct of MUX21_GENERIC_N4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_3;

architecture SYN_struct of MUX21_GENERIC_N4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_2;

architecture SYN_struct of MUX21_GENERIC_N4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_1;

architecture SYN_struct of MUX21_GENERIC_N4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_5;

architecture SYN_STRUCTURAL of carry_select_N4_5 is

   component MUX21_GENERIC_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_5 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_4;

architecture SYN_STRUCTURAL of carry_select_N4_4 is

   component MUX21_GENERIC_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_4 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_3;

architecture SYN_STRUCTURAL of carry_select_N4_3 is

   component MUX21_GENERIC_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_3 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_2;

architecture SYN_STRUCTURAL of carry_select_N4_2 is

   component MUX21_GENERIC_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_2 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_1;

architecture SYN_STRUCTURAL of carry_select_N4_1 is

   component MUX21_GENERIC_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_62_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62_1;

architecture SYN_BEHAVIORAL of FA_62_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_14_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_14_1;

architecture SYN_STRUCTURAL of rca_generic_N4_14_1 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_21_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_21_1;

architecture SYN_STRUCTURAL of PG_21_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_24_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_24_1;

architecture SYN_STRUCTURAL of PG_24_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n6);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_5_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_5_1;

architecture SYN_STRUCTURAL of G_5_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_30_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_30_1;

architecture SYN_STRUCTURAL of PGnet_block_30_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_94_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94_1;

architecture SYN_ARCH1 of ND2_94_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_30_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30_1;

architecture SYN_BEHAVIORAL of IV_30_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_30_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30_1;

architecture SYN_STRUCTURAL of MUX21_30_1 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30_1 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_6_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6_1;

architecture SYN_struct of MUX21_GENERIC_N4_6_1 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_6_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_6_1;

architecture SYN_STRUCTURAL of carry_select_N4_6_1 is

   component MUX21_GENERIC_N4_6_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_6_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_63_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63_1;

architecture SYN_BEHAVIORAL of FA_63_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_15_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_15_1;

architecture SYN_STRUCTURAL of rca_generic_N4_15_1 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_25_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_25_1;

architecture SYN_STRUCTURAL of PG_25_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n9);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_22_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_22_1;

architecture SYN_STRUCTURAL of PG_22_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_26_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_26_1;

architecture SYN_STRUCTURAL of PG_26_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n7);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_18_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_18_1;

architecture SYN_STRUCTURAL of PG_18_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n8, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_37 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_37;

architecture SYN_STRUCTURAL of PG_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_34 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_34;

architecture SYN_STRUCTURAL of PG_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_33 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_33;

architecture SYN_STRUCTURAL of PG_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_30 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_30;

architecture SYN_STRUCTURAL of PG_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_28 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_28;

architecture SYN_STRUCTURAL of PG_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_23 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_23;

architecture SYN_STRUCTURAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_19 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_19;

architecture SYN_STRUCTURAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U2 : INV_X1 port map( A => n8, ZN => gout);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_15 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_15;

architecture SYN_STRUCTURAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_14 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_14;

architecture SYN_STRUCTURAL of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_13 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_13;

architecture SYN_STRUCTURAL of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_1;

architecture SYN_STRUCTURAL of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_4_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_4_1;

architecture SYN_STRUCTURAL of PG_4_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n6);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_1;

architecture SYN_STRUCTURAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n11 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n11, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n11);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_8_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_8_1;

architecture SYN_STRUCTURAL of G_8_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n6);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_6_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_6_1;

architecture SYN_STRUCTURAL of G_6_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n6);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_31_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_31_1;

architecture SYN_STRUCTURAL of PGnet_block_31_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_95_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95_1;

architecture SYN_ARCH1 of ND2_95_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_31_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31_1;

architecture SYN_BEHAVIORAL of IV_31_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_31_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31_1;

architecture SYN_STRUCTURAL of MUX21_31_1 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31_1 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_7_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7_1;

architecture SYN_struct of MUX21_GENERIC_N4_7_1 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_7_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_7_1;

architecture SYN_STRUCTURAL of carry_select_N4_7_1 is

   component MUX21_GENERIC_N4_7_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_14_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_14_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_7_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_0_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_1;

architecture SYN_BEHAVIORAL of FA_0_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n7, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_0_1;

architecture SYN_STRUCTURAL of rca_generic_N4_0_1 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0_1 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63_1 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_62_1 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_0_1 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_0_1;

architecture SYN_STRUCTURAL of PG_0_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n8);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_0_1 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_0_1;

architecture SYN_STRUCTURAL of G_0_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_0_1 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_0_1;

architecture SYN_STRUCTURAL of PGnet_block_0_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_0_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0_1;

architecture SYN_ARCH1 of ND2_0_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_0_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0_1;

architecture SYN_BEHAVIORAL of IV_0_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_0_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0_1;

architecture SYN_STRUCTURAL of MUX21_0_1 is

   component ND2_94_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0_1 port map( A => S, Y => SB);
   UND1 : ND2_0_1 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95_1 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0_1;

architecture SYN_struct of MUX21_GENERIC_N4_0_1 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_0_1 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_31_1 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_30_1 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_0_1;

architecture SYN_STRUCTURAL of carry_select_N4_0_1 is

   component MUX21_GENERIC_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_15_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_15_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_0_1 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_31;

architecture SYN_behav of xor_gate_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_30;

architecture SYN_behav of xor_gate_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_29;

architecture SYN_behav of xor_gate_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_28;

architecture SYN_behav of xor_gate_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_27;

architecture SYN_behav of xor_gate_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_26;

architecture SYN_behav of xor_gate_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_25;

architecture SYN_behav of xor_gate_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_24;

architecture SYN_behav of xor_gate_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_23;

architecture SYN_behav of xor_gate_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_22;

architecture SYN_behav of xor_gate_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_21;

architecture SYN_behav of xor_gate_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_20;

architecture SYN_behav of xor_gate_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_19;

architecture SYN_behav of xor_gate_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_18;

architecture SYN_behav of xor_gate_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_17;

architecture SYN_behav of xor_gate_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_16;

architecture SYN_behav of xor_gate_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_15;

architecture SYN_behav of xor_gate_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_14;

architecture SYN_behav of xor_gate_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_13;

architecture SYN_behav of xor_gate_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_12;

architecture SYN_behav of xor_gate_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_11;

architecture SYN_behav of xor_gate_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_10;

architecture SYN_behav of xor_gate_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_9;

architecture SYN_behav of xor_gate_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_8;

architecture SYN_behav of xor_gate_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_7;

architecture SYN_behav of xor_gate_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_6;

architecture SYN_behav of xor_gate_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_5;

architecture SYN_behav of xor_gate_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_4;

architecture SYN_behav of xor_gate_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_3;

architecture SYN_behav of xor_gate_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_2;

architecture SYN_behav of xor_gate_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_1;

architecture SYN_behav of xor_gate_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity sum_generator_Nbits32_Nblocks8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Carry : in std_logic_vector
         (8 downto 0);  S : out std_logic_vector (31 downto 0);  Cout : out 
         std_logic);

end sum_generator_Nbits32_Nblocks8_1;

architecture SYN_STRUCTURAL of sum_generator_Nbits32_Nblocks8_1 is

   component carry_select_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(8);
   
   CS_0 : carry_select_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Carry(0), S(3) => S(3),
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4_7_1 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Carry(1), S(3) => S(7),
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4_6_1 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Carry(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Carry(3), S(3) 
                           => S(15), S(2) => S(14), S(1) => S(13), S(0) => 
                           S(12));
   CS_4 : carry_select_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Carry(4), S(3) 
                           => S(19), S(2) => S(18), S(1) => S(17), S(0) => 
                           S(16));
   CS_5 : carry_select_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Carry(5), S(3) 
                           => S(23), S(2) => S(22), S(1) => S(21), S(0) => 
                           S(20));
   CS_6 : carry_select_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Carry(6), S(3) 
                           => S(27), S(2) => S(26), S(1) => S(25), S(0) => 
                           S(24));
   CS_7 : carry_select_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Carry(7), S(3) 
                           => S(31), S(2) => S(30), S(1) => S(29), S(0) => 
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_generator_N32_Nblocks8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_Nblocks8_1;

architecture SYN_STRUCTURAL of carry_generator_N32_Nblocks8_1 is

   component G_3
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_4
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_7
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_9
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_2
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_5_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_6_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_3
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_4_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_13
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_5
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_6
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_14
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_15
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_16
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_17
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_19
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_8_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_7
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_8
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_9
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_10
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_20
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_18_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_11
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_23
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_21_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_22_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_12
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_24_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_25_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_26_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_0_1
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_2
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_2
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_3
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_4
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_5
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_6
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_7
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_8
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_9
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_10
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_11
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_12
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_13
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_14
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_15
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_16
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_17
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_18
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_19
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_20
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_21
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_22
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_23
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_24
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_25
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_26
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_27
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_28
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_29
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_30_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_31_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_0_1
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_0_1
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   signal Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_3_port, 
      g_cin, p_cin, Gsignal_1_31_port, Gsignal_1_30_port, Gsignal_1_29_port, 
      Gsignal_1_28_port, Gsignal_1_27_port, Gsignal_1_26_port, 
      Gsignal_1_25_port, Gsignal_1_24_port, Gsignal_1_23_port, 
      Gsignal_1_22_port, Gsignal_1_21_port, Gsignal_1_20_port, 
      Gsignal_1_19_port, Gsignal_1_18_port, Gsignal_1_17_port, 
      Gsignal_1_16_port, Gsignal_1_15_port, Gsignal_1_14_port, 
      Gsignal_1_13_port, Gsignal_1_12_port, Gsignal_1_11_port, 
      Gsignal_1_10_port, Gsignal_1_9_port, Gsignal_1_8_port, Gsignal_1_7_port, 
      Gsignal_1_6_port, Gsignal_1_5_port, Gsignal_1_4_port, Gsignal_1_3_port, 
      Gsignal_1_2_port, Gsignal_1_1_port, Gsignal_1_0_port, Gsignal_2_31_port, 
      Gsignal_2_29_port, Gsignal_2_27_port, Gsignal_2_25_port, 
      Gsignal_2_23_port, Gsignal_2_21_port, Gsignal_2_19_port, 
      Gsignal_2_17_port, Gsignal_2_15_port, Gsignal_2_13_port, 
      Gsignal_2_11_port, Gsignal_2_9_port, Gsignal_2_7_port, Gsignal_2_5_port, 
      Gsignal_2_3_port, Gsignal_2_1_port, Gsignal_3_31_port, Gsignal_3_23_port,
      Gsignal_3_15_port, Gsignal_3_7_port, Gsignal_4_31_port, Gsignal_4_15_port
      , Gsignal_5_31_port, Gsignal_5_27_port, Psignal_1_31_port, 
      Psignal_1_30_port, Psignal_1_29_port, Psignal_1_28_port, 
      Psignal_1_27_port, Psignal_1_26_port, Psignal_1_25_port, 
      Psignal_1_24_port, Psignal_1_23_port, Psignal_1_22_port, 
      Psignal_1_21_port, Psignal_1_20_port, Psignal_1_19_port, 
      Psignal_1_18_port, Psignal_1_17_port, Psignal_1_16_port, 
      Psignal_1_15_port, Psignal_1_14_port, Psignal_1_13_port, 
      Psignal_1_12_port, Psignal_1_11_port, Psignal_1_10_port, Psignal_1_9_port
      , Psignal_1_8_port, Psignal_1_7_port, Psignal_1_6_port, Psignal_1_5_port,
      Psignal_1_4_port, Psignal_1_3_port, Psignal_1_2_port, Psignal_1_1_port, 
      Psignal_2_31_port, Psignal_2_29_port, Psignal_2_27_port, 
      Psignal_2_25_port, Psignal_2_23_port, Psignal_2_21_port, 
      Psignal_2_19_port, Psignal_2_17_port, Psignal_2_15_port, 
      Psignal_2_13_port, Psignal_2_11_port, Psignal_2_9_port, Psignal_2_7_port,
      Psignal_2_5_port, Psignal_2_3_port, Psignal_3_31_port, Psignal_3_27_port,
      Psignal_3_23_port, Psignal_3_19_port, Psignal_3_15_port, Psignal_3_7_port
      , Psignal_4_31_port, Psignal_4_23_port, Psignal_4_15_port, 
      Psignal_5_31_port, Psignal_5_27_port, n8, Cout_1_port, n10, Cout_2_port, 
      n12, n13, n15, Cout_4_port : std_logic;

begin
   Cout <= ( Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, Ci );
   
   PGnet_Cin_0 : PGnet_block_0_1 port map( A => A(0), B => B(0), pout => p_cin,
                           gout => g_cin);
   GCin_0 : G_0_1 port map( gleft => g_cin, gright => Ci, pleft => p_cin, gout 
                           => Gsignal_1_0_port);
   PGnet_1 : PGnet_block_31_1 port map( A => A(1), B => B(1), pout => 
                           Psignal_1_1_port, gout => Gsignal_1_1_port);
   PGnet_2 : PGnet_block_30_1 port map( A => A(2), B => B(2), pout => 
                           Psignal_1_2_port, gout => Gsignal_1_2_port);
   PGnet_3 : PGnet_block_29 port map( A => A(3), B => B(3), pout => 
                           Psignal_1_3_port, gout => Gsignal_1_3_port);
   PGnet_4 : PGnet_block_28 port map( A => A(4), B => B(4), pout => 
                           Psignal_1_4_port, gout => Gsignal_1_4_port);
   PGnet_5 : PGnet_block_27 port map( A => A(5), B => B(5), pout => 
                           Psignal_1_5_port, gout => Gsignal_1_5_port);
   PGnet_6 : PGnet_block_26 port map( A => A(6), B => B(6), pout => 
                           Psignal_1_6_port, gout => Gsignal_1_6_port);
   PGnet_7 : PGnet_block_25 port map( A => A(7), B => B(7), pout => 
                           Psignal_1_7_port, gout => Gsignal_1_7_port);
   PGnet_8 : PGnet_block_24 port map( A => A(8), B => B(8), pout => 
                           Psignal_1_8_port, gout => Gsignal_1_8_port);
   PGnet_9 : PGnet_block_23 port map( A => A(9), B => B(9), pout => 
                           Psignal_1_9_port, gout => Gsignal_1_9_port);
   PGnet_10 : PGnet_block_22 port map( A => A(10), B => B(10), pout => 
                           Psignal_1_10_port, gout => Gsignal_1_10_port);
   PGnet_11 : PGnet_block_21 port map( A => A(11), B => B(11), pout => 
                           Psignal_1_11_port, gout => Gsignal_1_11_port);
   PGnet_12 : PGnet_block_20 port map( A => A(12), B => B(12), pout => 
                           Psignal_1_12_port, gout => Gsignal_1_12_port);
   PGnet_13 : PGnet_block_19 port map( A => A(13), B => B(13), pout => 
                           Psignal_1_13_port, gout => Gsignal_1_13_port);
   PGnet_14 : PGnet_block_18 port map( A => A(14), B => B(14), pout => 
                           Psignal_1_14_port, gout => Gsignal_1_14_port);
   PGnet_15 : PGnet_block_17 port map( A => A(15), B => B(15), pout => 
                           Psignal_1_15_port, gout => Gsignal_1_15_port);
   PGnet_16 : PGnet_block_16 port map( A => A(16), B => B(16), pout => 
                           Psignal_1_16_port, gout => Gsignal_1_16_port);
   PGnet_17 : PGnet_block_15 port map( A => A(17), B => B(17), pout => 
                           Psignal_1_17_port, gout => Gsignal_1_17_port);
   PGnet_18 : PGnet_block_14 port map( A => A(18), B => B(18), pout => 
                           Psignal_1_18_port, gout => Gsignal_1_18_port);
   PGnet_19 : PGnet_block_13 port map( A => A(19), B => B(19), pout => 
                           Psignal_1_19_port, gout => Gsignal_1_19_port);
   PGnet_20 : PGnet_block_12 port map( A => A(20), B => B(20), pout => 
                           Psignal_1_20_port, gout => Gsignal_1_20_port);
   PGnet_21 : PGnet_block_11 port map( A => A(21), B => B(21), pout => 
                           Psignal_1_21_port, gout => Gsignal_1_21_port);
   PGnet_22 : PGnet_block_10 port map( A => A(22), B => B(22), pout => 
                           Psignal_1_22_port, gout => Gsignal_1_22_port);
   PGnet_23 : PGnet_block_9 port map( A => A(23), B => B(23), pout => 
                           Psignal_1_23_port, gout => Gsignal_1_23_port);
   PGnet_24 : PGnet_block_8 port map( A => A(24), B => B(24), pout => 
                           Psignal_1_24_port, gout => Gsignal_1_24_port);
   PGnet_25 : PGnet_block_7 port map( A => A(25), B => B(25), pout => 
                           Psignal_1_25_port, gout => Gsignal_1_25_port);
   PGnet_26 : PGnet_block_6 port map( A => A(26), B => B(26), pout => 
                           Psignal_1_26_port, gout => Gsignal_1_26_port);
   PGnet_27 : PGnet_block_5 port map( A => A(27), B => B(27), pout => 
                           Psignal_1_27_port, gout => Gsignal_1_27_port);
   PGnet_28 : PGnet_block_4 port map( A => A(28), B => B(28), pout => 
                           Psignal_1_28_port, gout => Gsignal_1_28_port);
   PGnet_29 : PGnet_block_3 port map( A => A(29), B => B(29), pout => 
                           Psignal_1_29_port, gout => Gsignal_1_29_port);
   PGnet_30 : PGnet_block_2 port map( A => A(30), B => B(30), pout => 
                           Psignal_1_30_port, gout => Gsignal_1_30_port);
   PGnet_31 : PGnet_block_1 port map( A => A(31), B => B(31), pout => 
                           Psignal_1_31_port, gout => Gsignal_1_31_port);
   Gblock_1_1 : G_2 port map( gleft => Gsignal_1_1_port, gright => 
                           Gsignal_1_0_port, pleft => Psignal_1_1_port, gout =>
                           Gsignal_2_1_port);
   PGblock_1_3 : PG_0_1 port map( gleft => Gsignal_1_3_port, gright => 
                           Gsignal_1_2_port, pleft => Psignal_1_3_port, pright 
                           => Psignal_1_2_port, pout => Psignal_2_3_port, gout 
                           => Gsignal_2_3_port);
   PGblock_1_5 : PG_26_1 port map( gleft => Gsignal_1_5_port, gright => 
                           Gsignal_1_4_port, pleft => Psignal_1_5_port, pright 
                           => Psignal_1_4_port, pout => Psignal_2_5_port, gout 
                           => Gsignal_2_5_port);
   PGblock_1_7 : PG_25_1 port map( gleft => Gsignal_1_7_port, gright => 
                           Gsignal_1_6_port, pleft => Psignal_1_7_port, pright 
                           => Psignal_1_6_port, pout => Psignal_2_7_port, gout 
                           => Gsignal_2_7_port);
   PGblock_1_9 : PG_24_1 port map( gleft => Gsignal_1_9_port, gright => 
                           Gsignal_1_8_port, pleft => Psignal_1_9_port, pright 
                           => Psignal_1_8_port, pout => Psignal_2_9_port, gout 
                           => Gsignal_2_9_port);
   PGblock_1_11 : PG_12 port map( gleft => Gsignal_1_11_port, gright => 
                           Gsignal_1_10_port, pleft => Psignal_1_11_port, 
                           pright => Psignal_1_10_port, pout => 
                           Psignal_2_11_port, gout => Gsignal_2_11_port);
   PGblock_1_13 : PG_22_1 port map( gleft => Gsignal_1_13_port, gright => 
                           Gsignal_1_12_port, pleft => Psignal_1_13_port, 
                           pright => Psignal_1_12_port, pout => 
                           Psignal_2_13_port, gout => Gsignal_2_13_port);
   PGblock_1_15 : PG_21_1 port map( gleft => Gsignal_1_15_port, gright => 
                           Gsignal_1_14_port, pleft => Psignal_1_15_port, 
                           pright => Psignal_1_14_port, pout => 
                           Psignal_2_15_port, gout => Gsignal_2_15_port);
   PGblock_1_17 : PG_23 port map( gleft => Gsignal_1_17_port, gright => 
                           Gsignal_1_16_port, pleft => Psignal_1_17_port, 
                           pright => Psignal_1_16_port, pout => 
                           Psignal_2_17_port, gout => Gsignal_2_17_port);
   PGblock_1_19 : PG_11 port map( gleft => Gsignal_1_19_port, gright => 
                           Gsignal_1_18_port, pleft => Psignal_1_19_port, 
                           pright => Psignal_1_18_port, pout => 
                           Psignal_2_19_port, gout => Gsignal_2_19_port);
   PGblock_1_21 : PG_18_1 port map( gleft => Gsignal_1_21_port, gright => 
                           Gsignal_1_20_port, pleft => Psignal_1_21_port, 
                           pright => Psignal_1_20_port, pout => 
                           Psignal_2_21_port, gout => Gsignal_2_21_port);
   PGblock_1_23 : PG_20 port map( gleft => Gsignal_1_23_port, gright => 
                           Gsignal_1_22_port, pleft => Psignal_1_23_port, 
                           pright => Psignal_1_22_port, pout => 
                           Psignal_2_23_port, gout => Gsignal_2_23_port);
   PGblock_1_25 : PG_10 port map( gleft => Gsignal_1_25_port, gright => 
                           Gsignal_1_24_port, pleft => Psignal_1_25_port, 
                           pright => Psignal_1_24_port, pout => 
                           Psignal_2_25_port, gout => Gsignal_2_25_port);
   PGblock_1_27 : PG_9 port map( gleft => Gsignal_1_27_port, gright => 
                           Gsignal_1_26_port, pleft => Psignal_1_27_port, 
                           pright => Psignal_1_26_port, pout => 
                           Psignal_2_27_port, gout => Gsignal_2_27_port);
   PGblock_1_29 : PG_8 port map( gleft => Gsignal_1_29_port, gright => 
                           Gsignal_1_28_port, pleft => Psignal_1_29_port, 
                           pright => Psignal_1_28_port, pout => 
                           Psignal_2_29_port, gout => Gsignal_2_29_port);
   PGblock_1_31 : PG_7 port map( gleft => Gsignal_1_31_port, gright => 
                           Gsignal_1_30_port, pleft => Psignal_1_31_port, 
                           pright => Psignal_1_30_port, pout => 
                           Psignal_2_31_port, gout => Gsignal_2_31_port);
   Gblock_2_3 : G_8_1 port map( gleft => Gsignal_2_3_port, gright => 
                           Gsignal_2_1_port, pleft => Psignal_2_3_port, gout =>
                           Cout_1_port);
   PGblock_2_7 : PG_19 port map( gleft => Gsignal_2_7_port, gright => 
                           Gsignal_2_5_port, pleft => Psignal_2_7_port, pright 
                           => Psignal_2_5_port, pout => Psignal_3_7_port, gout 
                           => Gsignal_3_7_port);
   PGblock_2_11 : PG_17 port map( gleft => Gsignal_2_11_port, gright => 
                           Gsignal_2_9_port, pleft => Psignal_2_11_port, pright
                           => Psignal_2_9_port, pout => n8, gout => n10);
   PGblock_2_15 : PG_16 port map( gleft => Gsignal_2_15_port, gright => 
                           Gsignal_2_13_port, pleft => Psignal_2_15_port, 
                           pright => Psignal_2_13_port, pout => 
                           Psignal_3_15_port, gout => Gsignal_3_15_port);
   PGblock_2_19 : PG_15 port map( gleft => Gsignal_2_19_port, gright => 
                           Gsignal_2_17_port, pleft => Psignal_2_19_port, 
                           pright => Psignal_2_17_port, pout => 
                           Psignal_3_19_port, gout => n13);
   PGblock_2_23 : PG_14 port map( gleft => Gsignal_2_23_port, gright => 
                           Gsignal_2_21_port, pleft => Psignal_2_23_port, 
                           pright => Psignal_2_21_port, pout => 
                           Psignal_3_23_port, gout => Gsignal_3_23_port);
   PGblock_2_27 : PG_6 port map( gleft => Gsignal_2_27_port, gright => 
                           Gsignal_2_25_port, pleft => Psignal_2_27_port, 
                           pright => Psignal_2_25_port, pout => 
                           Psignal_3_27_port, gout => n12);
   PGblock_2_31 : PG_5 port map( gleft => Gsignal_2_31_port, gright => 
                           Gsignal_2_29_port, pleft => Psignal_2_31_port, 
                           pright => Psignal_2_29_port, pout => 
                           Psignal_3_31_port, gout => Gsignal_3_31_port);
   Gblock_3_7 : G_1 port map( gleft => Gsignal_3_7_port, gright => Cout_1_port,
                           pleft => Psignal_3_7_port, gout => Cout_2_port);
   PGblock_3_15 : PG_13 port map( gleft => Gsignal_3_15_port, gright => n10, 
                           pleft => Psignal_3_15_port, pright => n8, pout => 
                           Psignal_4_15_port, gout => Gsignal_4_15_port);
   PGblock_3_23 : PG_4_1 port map( gleft => Gsignal_3_23_port, gright => n13, 
                           pleft => Psignal_3_23_port, pright => 
                           Psignal_3_19_port, pout => Psignal_4_23_port, gout 
                           => n15);
   PGblock_3_31 : PG_3 port map( gleft => Gsignal_3_31_port, gright => n12, 
                           pleft => Psignal_3_31_port, pright => 
                           Psignal_3_27_port, pout => Psignal_4_31_port, gout 
                           => Gsignal_4_31_port);
   Gblock_4_11 : G_6_1 port map( gleft => n10, gright => Cout_2_port, pleft => 
                           n8, gout => Cout_3_port);
   Gblock_4_15 : G_5_1 port map( gleft => Gsignal_4_15_port, gright => 
                           Cout_2_port, pleft => Psignal_4_15_port, gout => 
                           Cout_4_port);
   PGblock_4_27 : PG_1 port map( gleft => n12, gright => n15, pleft => 
                           Psignal_3_27_port, pright => Psignal_4_23_port, pout
                           => Psignal_5_27_port, gout => Gsignal_5_27_port);
   PGblock_4_31 : PG_2 port map( gleft => Gsignal_4_31_port, gright => n15, 
                           pleft => Psignal_4_31_port, pright => 
                           Psignal_4_23_port, pout => Psignal_5_31_port, gout 
                           => Gsignal_5_31_port);
   Gblock_5_19 : G_9 port map( gleft => n13, gright => Cout_4_port, pleft => 
                           Psignal_3_19_port, gout => Cout_5_port);
   Gblock_5_23 : G_7 port map( gleft => n15, gright => Cout_4_port, pleft => 
                           Psignal_4_23_port, gout => Cout_6_port);
   Gblock_5_27 : G_4 port map( gleft => Gsignal_5_27_port, gright => 
                           Cout_4_port, pleft => Psignal_5_27_port, gout => 
                           Cout_7_port);
   Gblock_5_31 : G_3 port map( gleft => Gsignal_5_31_port, gright => 
                           Cout_4_port, pleft => Psignal_5_31_port, gout => 
                           Cout_8_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity cla_adder_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end cla_adder_N32_1;

architecture SYN_struct of cla_adder_N32_1 is

   component sum_generator_Nbits32_Nblocks8_1
      port( A, B : in std_logic_vector (31 downto 0);  Carry : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_Nblocks8_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal Carry_8_port, Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port,
      Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port : std_logic;

begin
   
   CG : carry_generator_N32_Nblocks8_1 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci, Cout(8) => 
                           Carry_8_port, Cout(7) => Carry_7_port, Cout(6) => 
                           Carry_6_port, Cout(5) => Carry_5_port, Cout(4) => 
                           Carry_4_port, Cout(3) => Carry_3_port, Cout(2) => 
                           Carry_2_port, Cout(1) => Carry_1_port, Cout(0) => 
                           Carry_0_port);
   SG : sum_generator_Nbits32_Nblocks8_1 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Carry(8) => Carry_8_port, 
                           Carry(7) => Carry_7_port, Carry(6) => Carry_6_port, 
                           Carry(5) => Carry_5_port, Carry(4) => Carry_4_port, 
                           Carry(3) => Carry_3_port, Carry(2) => Carry_2_port, 
                           Carry(1) => Carry_1_port, Carry(0) => Carry_0_port, 
                           S(31) => Sum(31), S(30) => Sum(30), S(29) => Sum(29)
                           , S(28) => Sum(28), S(27) => Sum(27), S(26) => 
                           Sum(26), S(25) => Sum(25), S(24) => Sum(24), S(23) 
                           => Sum(23), S(22) => Sum(22), S(21) => Sum(21), 
                           S(20) => Sum(20), S(19) => Sum(19), S(18) => Sum(18)
                           , S(17) => Sum(17), S(16) => Sum(16), S(15) => 
                           Sum(15), S(14) => Sum(14), S(13) => Sum(13), S(12) 
                           => Sum(12), S(11) => Sum(11), S(10) => Sum(10), S(9)
                           => Sum(9), S(8) => Sum(8), S(7) => Sum(7), S(6) => 
                           Sum(6), S(5) => Sum(5), S(4) => Sum(4), S(3) => 
                           Sum(3), S(2) => Sum(2), S(1) => Sum(1), S(0) => 
                           Sum(0), Cout => Cout);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n16, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n16);
   U1 : INV_X1 port map( A => n15, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n16, B2 => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n16, n17 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n17, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n17);
   U1 : INV_X1 port map( A => n16, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n17, B2 => Ci, ZN => n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n13, n14 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n14, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U1 : INV_X1 port map( A => n13, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n14, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n13, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n13);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n13, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n14, n15 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n15, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n15);
   U1 : INV_X1 port map( A => n14, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n15, B2 => Ci, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);
   U1 : INV_X1 port map( A => n11, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n10, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : INV_X1 port map( A => n9, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_30_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30_0;

architecture SYN_BEHAVIORAL of IV_30_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH1 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_31_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31_0;

architecture SYN_BEHAVIORAL of IV_31_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_94_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94_0;

architecture SYN_ARCH1 of ND2_94_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_95_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95_0;

architecture SYN_ARCH1 of ND2_95_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity ND2_0_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0_0;

architecture SYN_ARCH1 of ND2_0_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity IV_0_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0_0;

architecture SYN_BEHAVIORAL of IV_0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_182 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_181 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_180 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_30_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30_0;

architecture SYN_STRUCTURAL of MUX21_30_0 is

   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30_0 port map( A => S, Y => SB);
   UND1 : ND2_185 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_184 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_183 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_31_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31_0;

architecture SYN_STRUCTURAL of MUX21_31_0 is

   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31_0 port map( A => S, Y => SB);
   UND1 : ND2_188 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_187 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_186 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_0_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0_0;

architecture SYN_STRUCTURAL of MUX21_0_0 is

   component ND2_94_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0_0 port map( A => S, Y => SB);
   UND1 : ND2_0_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95_0 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94_0 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_62_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62_0;

architecture SYN_BEHAVIORAL of FA_62_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_63_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63_0;

architecture SYN_BEHAVIORAL of FA_63_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_0_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_0;

architecture SYN_BEHAVIORAL of FA_0_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_16;

architecture SYN_STRUCTURAL of rca_generic_N4_16 is

   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_259 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_258 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_257 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_256 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_17;

architecture SYN_STRUCTURAL of rca_generic_N4_17 is

   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_263 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_262 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_261 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_260 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_18;

architecture SYN_STRUCTURAL of rca_generic_N4_18 is

   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_267 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_266 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_265 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_264 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_19;

architecture SYN_STRUCTURAL of rca_generic_N4_19 is

   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_271 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_270 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_269 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_268 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_12;

architecture SYN_struct of MUX21_GENERIC_N4_12 is

   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_51 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_50 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_49 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_48 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_24;

architecture SYN_STRUCTURAL of rca_generic_N4_24 is

   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_291 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_290 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_289 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_288 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_6_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6_0;

architecture SYN_struct of MUX21_GENERIC_N4_6_0 is

   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_55 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_54 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_53 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_52 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_7_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7_0;

architecture SYN_struct of MUX21_GENERIC_N4_7_0 is

   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_59 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_58 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_57 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_56 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_28;

architecture SYN_STRUCTURAL of rca_generic_N4_28 is

   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_307 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_306 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_305 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_304 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_14_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_14_0;

architecture SYN_STRUCTURAL of rca_generic_N4_14_0 is

   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_311 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_310 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_309 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_308 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity MUX21_GENERIC_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0_0;

architecture SYN_struct of MUX21_GENERIC_N4_0_0 is

   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   M_0 : MUX21_0_0 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   M_1 : MUX21_31_0 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   M_2 : MUX21_30_0 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   M_3 : MUX21_60 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_15_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_15_0;

architecture SYN_STRUCTURAL of rca_generic_N4_15_0 is

   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_315 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_314 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_313 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_312 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity rca_generic_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end rca_generic_N4_0_0;

architecture SYN_STRUCTURAL of rca_generic_N4_0_0 is

   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63_0 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_62_0 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_316 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_8;

architecture SYN_STRUCTURAL of carry_select_N4_8 is

   component MUX21_GENERIC_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_8 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_9;

architecture SYN_STRUCTURAL of carry_select_N4_9 is

   component MUX21_GENERIC_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_9 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_10;

architecture SYN_STRUCTURAL of carry_select_N4_10 is

   component MUX21_GENERIC_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_10 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_11;

architecture SYN_STRUCTURAL of carry_select_N4_11 is

   component MUX21_GENERIC_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_11 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_12;

architecture SYN_STRUCTURAL of carry_select_N4_12 is

   component MUX21_GENERIC_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_12 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_6_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_6_0;

architecture SYN_STRUCTURAL of carry_select_N4_6_0 is

   component MUX21_GENERIC_N4_6_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_6_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_7_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_7_0;

architecture SYN_STRUCTURAL of carry_select_N4_7_0 is

   component MUX21_GENERIC_N4_7_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_14_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_14_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_7_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_select_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_0_0;

architecture SYN_STRUCTURAL of carry_select_N4_0_0 is

   component MUX21_GENERIC_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component rca_generic_N4_15_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component rca_generic_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum_carry0_3_port, sum_carry0_2_port, 
      sum_carry0_1_port, sum_carry0_0_port, sum_carry1_3_port, 
      sum_carry1_2_port, sum_carry1_1_port, sum_carry1_0_port, net6204, net6205
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : rca_generic_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum_carry0_3_port, S(2) => sum_carry0_2_port, S(1) 
                           => sum_carry0_1_port, S(0) => sum_carry0_0_port, Co 
                           => net6205);
   RCA1 : rca_generic_N4_15_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum_carry1_3_port, S(2) => sum_carry1_2_port, S(1) 
                           => sum_carry1_1_port, S(0) => sum_carry1_0_port, Co 
                           => net6204);
   MUX : MUX21_GENERIC_N4_0_0 port map( A(3) => sum_carry1_3_port, A(2) => 
                           sum_carry1_2_port, A(1) => sum_carry1_1_port, A(0) 
                           => sum_carry1_0_port, B(3) => sum_carry0_3_port, 
                           B(2) => sum_carry0_2_port, B(1) => sum_carry0_1_port
                           , B(0) => sum_carry0_0_port, SEL => Ci, Y(3) => S(3)
                           , Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_13 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_13;

architecture SYN_STRUCTURAL of G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_5_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_5_0;

architecture SYN_STRUCTURAL of G_5_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_6_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_6_0;

architecture SYN_STRUCTURAL of G_6_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_4_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_4_0;

architecture SYN_STRUCTURAL of PG_4_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_14 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_14;

architecture SYN_STRUCTURAL of G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_36 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_36;

architecture SYN_STRUCTURAL of PG_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_8_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_8_0;

architecture SYN_STRUCTURAL of G_8_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_42 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_42;

architecture SYN_STRUCTURAL of PG_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_18_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_18_0;

architecture SYN_STRUCTURAL of PG_18_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_44 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_44;

architecture SYN_STRUCTURAL of PG_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_21_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_21_0;

architecture SYN_STRUCTURAL of PG_21_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);
   U2 : INV_X1 port map( A => n2, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_22_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_22_0;

architecture SYN_STRUCTURAL of PG_22_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_45 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_45;

architecture SYN_STRUCTURAL of PG_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_24_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_24_0;

architecture SYN_STRUCTURAL of PG_24_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_25_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_25_0;

architecture SYN_STRUCTURAL of PG_25_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_26_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_26_0;

architecture SYN_STRUCTURAL of PG_26_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PG_0_0 is

   port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
         std_logic);

end PG_0_0;

architecture SYN_STRUCTURAL of PG_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gright, B2 => pleft, A => gleft, ZN => n2);
   U3 : AND2_X1 port map( A1 => pright, A2 => pleft, ZN => pout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_15 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_15;

architecture SYN_STRUCTURAL of G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_60 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_60;

architecture SYN_STRUCTURAL of PGnet_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_30_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_30_0;

architecture SYN_STRUCTURAL of PGnet_block_30_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_31_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_31_0;

architecture SYN_STRUCTURAL of PGnet_block_31_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity G_0_0 is

   port( gleft, gright, pleft : in std_logic;  gout : out std_logic);

end G_0_0;

architecture SYN_STRUCTURAL of G_0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => pleft, B2 => gright, A => gleft, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity PGnet_block_0_0 is

   port( A, B : in std_logic;  pout, gout : out std_logic);

end PGnet_block_0_0;

architecture SYN_STRUCTURAL of PGnet_block_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => pout);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => gout);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => A, A2 => B, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity sum_generator_Nbits32_Nblocks8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Carry : in std_logic_vector
         (8 downto 0);  S : out std_logic_vector (31 downto 0);  Cout : out 
         std_logic);

end sum_generator_Nbits32_Nblocks8_0;

architecture SYN_STRUCTURAL of sum_generator_Nbits32_Nblocks8_0 is

   component carry_select_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(8);
   
   CS_0 : carry_select_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Carry(0), S(3) => S(3),
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4_7_0 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Carry(1), S(3) => S(7),
                           S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4_6_0 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Carry(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4_12 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Carry(3), S(3) 
                           => S(15), S(2) => S(14), S(1) => S(13), S(0) => 
                           S(12));
   CS_4 : carry_select_N4_11 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Carry(4), S(3) 
                           => S(19), S(2) => S(18), S(1) => S(17), S(0) => 
                           S(16));
   CS_5 : carry_select_N4_10 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Carry(5), S(3) 
                           => S(23), S(2) => S(22), S(1) => S(21), S(0) => 
                           S(20));
   CS_6 : carry_select_N4_9 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Carry(6), S(3) 
                           => S(27), S(2) => S(26), S(1) => S(25), S(0) => 
                           S(24));
   CS_7 : carry_select_N4_8 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Carry(7), S(3) 
                           => S(31), S(2) => S(30), S(1) => S(29), S(0) => 
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity carry_generator_N32_Nblocks8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_Nblocks8_0;

architecture SYN_STRUCTURAL of carry_generator_N32_Nblocks8_0 is

   component G_10
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_11
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_12
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_13
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_27
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_28
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_5_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component G_6_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_29
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_4_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_30
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_14
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_31
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_32
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_33
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_34
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_35
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_36
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_37
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_8_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_38
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_39
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_40
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_41
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_42
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_18_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_43
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_44
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_21_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_22_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_45
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_24_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_25_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_26_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component PG_0_0
      port( gleft, gright, pleft, pright : in std_logic;  pout, gout : out 
            std_logic);
   end component;
   
   component G_15
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_32
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_33
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_34
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_35
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_36
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_37
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_38
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_39
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_40
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_41
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_42
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_43
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_44
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_45
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_46
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_47
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_48
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_49
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_50
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_51
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_52
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_53
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_54
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_55
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_56
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_57
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_58
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_59
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_60
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_30_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PGnet_block_31_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_0_0
      port( gleft, gright, pleft : in std_logic;  gout : out std_logic);
   end component;
   
   component PGnet_block_0_0
      port( A, B : in std_logic;  pout, gout : out std_logic);
   end component;
   
   signal Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_3_port, 
      g_cin, p_cin, Gsignal_1_31_port, Gsignal_1_30_port, Gsignal_1_29_port, 
      Gsignal_1_28_port, Gsignal_1_27_port, Gsignal_1_26_port, 
      Gsignal_1_25_port, Gsignal_1_24_port, Gsignal_1_23_port, 
      Gsignal_1_22_port, Gsignal_1_21_port, Gsignal_1_20_port, 
      Gsignal_1_19_port, Gsignal_1_18_port, Gsignal_1_17_port, 
      Gsignal_1_16_port, Gsignal_1_15_port, Gsignal_1_14_port, 
      Gsignal_1_13_port, Gsignal_1_12_port, Gsignal_1_11_port, 
      Gsignal_1_10_port, Gsignal_1_9_port, Gsignal_1_8_port, Gsignal_1_7_port, 
      Gsignal_1_6_port, Gsignal_1_5_port, Gsignal_1_4_port, Gsignal_1_3_port, 
      Gsignal_1_2_port, Gsignal_1_1_port, Gsignal_1_0_port, Gsignal_2_31_port, 
      Gsignal_2_29_port, Gsignal_2_27_port, Gsignal_2_25_port, 
      Gsignal_2_23_port, Gsignal_2_21_port, Gsignal_2_19_port, 
      Gsignal_2_17_port, Gsignal_2_15_port, Gsignal_2_13_port, 
      Gsignal_2_11_port, Gsignal_2_9_port, Gsignal_2_7_port, Gsignal_2_5_port, 
      Gsignal_2_3_port, Gsignal_2_1_port, Gsignal_3_31_port, Gsignal_3_23_port,
      Gsignal_3_15_port, Gsignal_3_7_port, Gsignal_4_31_port, Gsignal_4_15_port
      , Gsignal_5_31_port, Gsignal_5_27_port, Psignal_1_31_port, 
      Psignal_1_30_port, Psignal_1_29_port, Psignal_1_28_port, 
      Psignal_1_27_port, Psignal_1_26_port, Psignal_1_25_port, 
      Psignal_1_24_port, Psignal_1_23_port, Psignal_1_22_port, 
      Psignal_1_21_port, Psignal_1_20_port, Psignal_1_19_port, 
      Psignal_1_18_port, Psignal_1_17_port, Psignal_1_16_port, 
      Psignal_1_15_port, Psignal_1_14_port, Psignal_1_13_port, 
      Psignal_1_12_port, Psignal_1_11_port, Psignal_1_10_port, Psignal_1_9_port
      , Psignal_1_8_port, Psignal_1_7_port, Psignal_1_6_port, Psignal_1_5_port,
      Psignal_1_4_port, Psignal_1_3_port, Psignal_1_2_port, Psignal_1_1_port, 
      Psignal_2_31_port, Psignal_2_29_port, Psignal_2_27_port, 
      Psignal_2_25_port, Psignal_2_23_port, Psignal_2_21_port, 
      Psignal_2_19_port, Psignal_2_17_port, Psignal_2_15_port, 
      Psignal_2_13_port, Psignal_2_11_port, Psignal_2_9_port, Psignal_2_7_port,
      Psignal_2_5_port, Psignal_2_3_port, Psignal_3_31_port, Psignal_3_27_port,
      Psignal_3_23_port, Psignal_3_19_port, Psignal_3_15_port, Psignal_3_7_port
      , Psignal_4_31_port, Psignal_4_23_port, Psignal_4_15_port, 
      Psignal_5_31_port, Psignal_5_27_port, n8, Cout_1_port, n10, Cout_2_port, 
      n12, n13, n15, Cout_4_port : std_logic;

begin
   Cout <= ( Cout_8_port, Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, 
      Cout_3_port, Cout_2_port, Cout_1_port, Ci );
   
   PGnet_Cin_0 : PGnet_block_0_0 port map( A => A(0), B => B(0), pout => p_cin,
                           gout => g_cin);
   GCin_0 : G_0_0 port map( gleft => g_cin, gright => Ci, pleft => p_cin, gout 
                           => Gsignal_1_0_port);
   PGnet_1 : PGnet_block_31_0 port map( A => A(1), B => B(1), pout => 
                           Psignal_1_1_port, gout => Gsignal_1_1_port);
   PGnet_2 : PGnet_block_30_0 port map( A => A(2), B => B(2), pout => 
                           Psignal_1_2_port, gout => Gsignal_1_2_port);
   PGnet_3 : PGnet_block_60 port map( A => A(3), B => B(3), pout => 
                           Psignal_1_3_port, gout => Gsignal_1_3_port);
   PGnet_4 : PGnet_block_59 port map( A => A(4), B => B(4), pout => 
                           Psignal_1_4_port, gout => Gsignal_1_4_port);
   PGnet_5 : PGnet_block_58 port map( A => A(5), B => B(5), pout => 
                           Psignal_1_5_port, gout => Gsignal_1_5_port);
   PGnet_6 : PGnet_block_57 port map( A => A(6), B => B(6), pout => 
                           Psignal_1_6_port, gout => Gsignal_1_6_port);
   PGnet_7 : PGnet_block_56 port map( A => A(7), B => B(7), pout => 
                           Psignal_1_7_port, gout => Gsignal_1_7_port);
   PGnet_8 : PGnet_block_55 port map( A => A(8), B => B(8), pout => 
                           Psignal_1_8_port, gout => Gsignal_1_8_port);
   PGnet_9 : PGnet_block_54 port map( A => A(9), B => B(9), pout => 
                           Psignal_1_9_port, gout => Gsignal_1_9_port);
   PGnet_10 : PGnet_block_53 port map( A => A(10), B => B(10), pout => 
                           Psignal_1_10_port, gout => Gsignal_1_10_port);
   PGnet_11 : PGnet_block_52 port map( A => A(11), B => B(11), pout => 
                           Psignal_1_11_port, gout => Gsignal_1_11_port);
   PGnet_12 : PGnet_block_51 port map( A => A(12), B => B(12), pout => 
                           Psignal_1_12_port, gout => Gsignal_1_12_port);
   PGnet_13 : PGnet_block_50 port map( A => A(13), B => B(13), pout => 
                           Psignal_1_13_port, gout => Gsignal_1_13_port);
   PGnet_14 : PGnet_block_49 port map( A => A(14), B => B(14), pout => 
                           Psignal_1_14_port, gout => Gsignal_1_14_port);
   PGnet_15 : PGnet_block_48 port map( A => A(15), B => B(15), pout => 
                           Psignal_1_15_port, gout => Gsignal_1_15_port);
   PGnet_16 : PGnet_block_47 port map( A => A(16), B => B(16), pout => 
                           Psignal_1_16_port, gout => Gsignal_1_16_port);
   PGnet_17 : PGnet_block_46 port map( A => A(17), B => B(17), pout => 
                           Psignal_1_17_port, gout => Gsignal_1_17_port);
   PGnet_18 : PGnet_block_45 port map( A => A(18), B => B(18), pout => 
                           Psignal_1_18_port, gout => Gsignal_1_18_port);
   PGnet_19 : PGnet_block_44 port map( A => A(19), B => B(19), pout => 
                           Psignal_1_19_port, gout => Gsignal_1_19_port);
   PGnet_20 : PGnet_block_43 port map( A => A(20), B => B(20), pout => 
                           Psignal_1_20_port, gout => Gsignal_1_20_port);
   PGnet_21 : PGnet_block_42 port map( A => A(21), B => B(21), pout => 
                           Psignal_1_21_port, gout => Gsignal_1_21_port);
   PGnet_22 : PGnet_block_41 port map( A => A(22), B => B(22), pout => 
                           Psignal_1_22_port, gout => Gsignal_1_22_port);
   PGnet_23 : PGnet_block_40 port map( A => A(23), B => B(23), pout => 
                           Psignal_1_23_port, gout => Gsignal_1_23_port);
   PGnet_24 : PGnet_block_39 port map( A => A(24), B => B(24), pout => 
                           Psignal_1_24_port, gout => Gsignal_1_24_port);
   PGnet_25 : PGnet_block_38 port map( A => A(25), B => B(25), pout => 
                           Psignal_1_25_port, gout => Gsignal_1_25_port);
   PGnet_26 : PGnet_block_37 port map( A => A(26), B => B(26), pout => 
                           Psignal_1_26_port, gout => Gsignal_1_26_port);
   PGnet_27 : PGnet_block_36 port map( A => A(27), B => B(27), pout => 
                           Psignal_1_27_port, gout => Gsignal_1_27_port);
   PGnet_28 : PGnet_block_35 port map( A => A(28), B => B(28), pout => 
                           Psignal_1_28_port, gout => Gsignal_1_28_port);
   PGnet_29 : PGnet_block_34 port map( A => A(29), B => B(29), pout => 
                           Psignal_1_29_port, gout => Gsignal_1_29_port);
   PGnet_30 : PGnet_block_33 port map( A => A(30), B => B(30), pout => 
                           Psignal_1_30_port, gout => Gsignal_1_30_port);
   PGnet_31 : PGnet_block_32 port map( A => A(31), B => B(31), pout => 
                           Psignal_1_31_port, gout => Gsignal_1_31_port);
   Gblock_1_1 : G_15 port map( gleft => Gsignal_1_1_port, gright => 
                           Gsignal_1_0_port, pleft => Psignal_1_1_port, gout =>
                           Gsignal_2_1_port);
   PGblock_1_3 : PG_0_0 port map( gleft => Gsignal_1_3_port, gright => 
                           Gsignal_1_2_port, pleft => Psignal_1_3_port, pright 
                           => Psignal_1_2_port, pout => Psignal_2_3_port, gout 
                           => Gsignal_2_3_port);
   PGblock_1_5 : PG_26_0 port map( gleft => Gsignal_1_5_port, gright => 
                           Gsignal_1_4_port, pleft => Psignal_1_5_port, pright 
                           => Psignal_1_4_port, pout => Psignal_2_5_port, gout 
                           => Gsignal_2_5_port);
   PGblock_1_7 : PG_25_0 port map( gleft => Gsignal_1_7_port, gright => 
                           Gsignal_1_6_port, pleft => Psignal_1_7_port, pright 
                           => Psignal_1_6_port, pout => Psignal_2_7_port, gout 
                           => Gsignal_2_7_port);
   PGblock_1_9 : PG_24_0 port map( gleft => Gsignal_1_9_port, gright => 
                           Gsignal_1_8_port, pleft => Psignal_1_9_port, pright 
                           => Psignal_1_8_port, pout => Psignal_2_9_port, gout 
                           => Gsignal_2_9_port);
   PGblock_1_11 : PG_45 port map( gleft => Gsignal_1_11_port, gright => 
                           Gsignal_1_10_port, pleft => Psignal_1_11_port, 
                           pright => Psignal_1_10_port, pout => 
                           Psignal_2_11_port, gout => Gsignal_2_11_port);
   PGblock_1_13 : PG_22_0 port map( gleft => Gsignal_1_13_port, gright => 
                           Gsignal_1_12_port, pleft => Psignal_1_13_port, 
                           pright => Psignal_1_12_port, pout => 
                           Psignal_2_13_port, gout => Gsignal_2_13_port);
   PGblock_1_15 : PG_21_0 port map( gleft => Gsignal_1_15_port, gright => 
                           Gsignal_1_14_port, pleft => Psignal_1_15_port, 
                           pright => Psignal_1_14_port, pout => 
                           Psignal_2_15_port, gout => Gsignal_2_15_port);
   PGblock_1_17 : PG_44 port map( gleft => Gsignal_1_17_port, gright => 
                           Gsignal_1_16_port, pleft => Psignal_1_17_port, 
                           pright => Psignal_1_16_port, pout => 
                           Psignal_2_17_port, gout => Gsignal_2_17_port);
   PGblock_1_19 : PG_43 port map( gleft => Gsignal_1_19_port, gright => 
                           Gsignal_1_18_port, pleft => Psignal_1_19_port, 
                           pright => Psignal_1_18_port, pout => 
                           Psignal_2_19_port, gout => Gsignal_2_19_port);
   PGblock_1_21 : PG_18_0 port map( gleft => Gsignal_1_21_port, gright => 
                           Gsignal_1_20_port, pleft => Psignal_1_21_port, 
                           pright => Psignal_1_20_port, pout => 
                           Psignal_2_21_port, gout => Gsignal_2_21_port);
   PGblock_1_23 : PG_42 port map( gleft => Gsignal_1_23_port, gright => 
                           Gsignal_1_22_port, pleft => Psignal_1_23_port, 
                           pright => Psignal_1_22_port, pout => 
                           Psignal_2_23_port, gout => Gsignal_2_23_port);
   PGblock_1_25 : PG_41 port map( gleft => Gsignal_1_25_port, gright => 
                           Gsignal_1_24_port, pleft => Psignal_1_25_port, 
                           pright => Psignal_1_24_port, pout => 
                           Psignal_2_25_port, gout => Gsignal_2_25_port);
   PGblock_1_27 : PG_40 port map( gleft => Gsignal_1_27_port, gright => 
                           Gsignal_1_26_port, pleft => Psignal_1_27_port, 
                           pright => Psignal_1_26_port, pout => 
                           Psignal_2_27_port, gout => Gsignal_2_27_port);
   PGblock_1_29 : PG_39 port map( gleft => Gsignal_1_29_port, gright => 
                           Gsignal_1_28_port, pleft => Psignal_1_29_port, 
                           pright => Psignal_1_28_port, pout => 
                           Psignal_2_29_port, gout => Gsignal_2_29_port);
   PGblock_1_31 : PG_38 port map( gleft => Gsignal_1_31_port, gright => 
                           Gsignal_1_30_port, pleft => Psignal_1_31_port, 
                           pright => Psignal_1_30_port, pout => 
                           Psignal_2_31_port, gout => Gsignal_2_31_port);
   Gblock_2_3 : G_8_0 port map( gleft => Gsignal_2_3_port, gright => 
                           Gsignal_2_1_port, pleft => Psignal_2_3_port, gout =>
                           Cout_1_port);
   PGblock_2_7 : PG_37 port map( gleft => Gsignal_2_7_port, gright => 
                           Gsignal_2_5_port, pleft => Psignal_2_7_port, pright 
                           => Psignal_2_5_port, pout => Psignal_3_7_port, gout 
                           => Gsignal_3_7_port);
   PGblock_2_11 : PG_36 port map( gleft => Gsignal_2_11_port, gright => 
                           Gsignal_2_9_port, pleft => Psignal_2_11_port, pright
                           => Psignal_2_9_port, pout => n8, gout => n10);
   PGblock_2_15 : PG_35 port map( gleft => Gsignal_2_15_port, gright => 
                           Gsignal_2_13_port, pleft => Psignal_2_15_port, 
                           pright => Psignal_2_13_port, pout => 
                           Psignal_3_15_port, gout => Gsignal_3_15_port);
   PGblock_2_19 : PG_34 port map( gleft => Gsignal_2_19_port, gright => 
                           Gsignal_2_17_port, pleft => Psignal_2_19_port, 
                           pright => Psignal_2_17_port, pout => 
                           Psignal_3_19_port, gout => n13);
   PGblock_2_23 : PG_33 port map( gleft => Gsignal_2_23_port, gright => 
                           Gsignal_2_21_port, pleft => Psignal_2_23_port, 
                           pright => Psignal_2_21_port, pout => 
                           Psignal_3_23_port, gout => Gsignal_3_23_port);
   PGblock_2_27 : PG_32 port map( gleft => Gsignal_2_27_port, gright => 
                           Gsignal_2_25_port, pleft => Psignal_2_27_port, 
                           pright => Psignal_2_25_port, pout => 
                           Psignal_3_27_port, gout => n12);
   PGblock_2_31 : PG_31 port map( gleft => Gsignal_2_31_port, gright => 
                           Gsignal_2_29_port, pleft => Psignal_2_31_port, 
                           pright => Psignal_2_29_port, pout => 
                           Psignal_3_31_port, gout => Gsignal_3_31_port);
   Gblock_3_7 : G_14 port map( gleft => Gsignal_3_7_port, gright => Cout_1_port
                           , pleft => Psignal_3_7_port, gout => Cout_2_port);
   PGblock_3_15 : PG_30 port map( gleft => Gsignal_3_15_port, gright => n10, 
                           pleft => Psignal_3_15_port, pright => n8, pout => 
                           Psignal_4_15_port, gout => Gsignal_4_15_port);
   PGblock_3_23 : PG_4_0 port map( gleft => Gsignal_3_23_port, gright => n13, 
                           pleft => Psignal_3_23_port, pright => 
                           Psignal_3_19_port, pout => Psignal_4_23_port, gout 
                           => n15);
   PGblock_3_31 : PG_29 port map( gleft => Gsignal_3_31_port, gright => n12, 
                           pleft => Psignal_3_31_port, pright => 
                           Psignal_3_27_port, pout => Psignal_4_31_port, gout 
                           => Gsignal_4_31_port);
   Gblock_4_11 : G_6_0 port map( gleft => n10, gright => Cout_2_port, pleft => 
                           n8, gout => Cout_3_port);
   Gblock_4_15 : G_5_0 port map( gleft => Gsignal_4_15_port, gright => 
                           Cout_2_port, pleft => Psignal_4_15_port, gout => 
                           Cout_4_port);
   PGblock_4_27 : PG_28 port map( gleft => n12, gright => n15, pleft => 
                           Psignal_3_27_port, pright => Psignal_4_23_port, pout
                           => Psignal_5_27_port, gout => Gsignal_5_27_port);
   PGblock_4_31 : PG_27 port map( gleft => Gsignal_4_31_port, gright => n15, 
                           pleft => Psignal_4_31_port, pright => 
                           Psignal_4_23_port, pout => Psignal_5_31_port, gout 
                           => Gsignal_5_31_port);
   Gblock_5_19 : G_13 port map( gleft => n13, gright => Cout_4_port, pleft => 
                           Psignal_3_19_port, gout => Cout_5_port);
   Gblock_5_23 : G_12 port map( gleft => n15, gright => Cout_4_port, pleft => 
                           Psignal_4_23_port, gout => Cout_6_port);
   Gblock_5_27 : G_11 port map( gleft => Gsignal_5_27_port, gright => 
                           Cout_4_port, pleft => Psignal_5_27_port, gout => 
                           Cout_7_port);
   Gblock_5_31 : G_10 port map( gleft => Gsignal_5_31_port, gright => 
                           Cout_4_port, pleft => Psignal_5_31_port, gout => 
                           Cout_8_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity xor_gate_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end xor_gate_0;

architecture SYN_behav of xor_gate_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => Y);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_thirdLevel is

   port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector (38 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end shift_thirdLevel;

architecture SYN_behav of shift_thirdLevel is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n40, n41, n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
      n56, n57, n58, n59, n60, n61, n62, n63, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(2), A2 => n148, ZN => n149);
   U2 : INV_X1 port map( A => n157, ZN => n156);
   U3 : INV_X1 port map( A => n149, ZN => n154);
   U4 : INV_X1 port map( A => n161, ZN => n158);
   U5 : INV_X1 port map( A => n153, ZN => n152);
   U6 : INV_X1 port map( A => n149, ZN => n155);
   U7 : OAI22_X1 port map( A1 => n165, A2 => n126, B1 => sel(0), B2 => n123, ZN
                           => Y(15));
   U8 : OAI22_X1 port map( A1 => n166, A2 => n129, B1 => sel(0), B2 => n126, ZN
                           => Y(14));
   U9 : OAI22_X1 port map( A1 => n166, A2 => n132, B1 => sel(0), B2 => n129, ZN
                           => Y(13));
   U10 : OAI22_X1 port map( A1 => n166, A2 => n135, B1 => sel(0), B2 => n132, 
                           ZN => Y(12));
   U11 : OAI22_X1 port map( A1 => n166, A2 => n138, B1 => sel(0), B2 => n135, 
                           ZN => Y(11));
   U12 : INV_X1 port map( A => n151, ZN => n150);
   U13 : OAI22_X1 port map( A1 => sel(0), A2 => n40, B1 => n41, B2 => n159, ZN 
                           => Y(9));
   U14 : OAI22_X1 port map( A1 => n161, A2 => n83, B1 => n158, B2 => n74, ZN =>
                           Y(29));
   U15 : OAI22_X1 port map( A1 => n162, A2 => n86, B1 => n158, B2 => n83, ZN =>
                           Y(28));
   U16 : OAI22_X1 port map( A1 => n162, A2 => n89, B1 => n158, B2 => n86, ZN =>
                           Y(27));
   U17 : OAI22_X1 port map( A1 => n162, A2 => n91, B1 => n158, B2 => n89, ZN =>
                           Y(26));
   U18 : OAI22_X1 port map( A1 => n162, A2 => n93, B1 => n158, B2 => n91, ZN =>
                           Y(25));
   U19 : OAI22_X1 port map( A1 => n163, A2 => n96, B1 => n158, B2 => n93, ZN =>
                           Y(24));
   U20 : OAI22_X1 port map( A1 => n163, A2 => n99, B1 => n158, B2 => n96, ZN =>
                           Y(23));
   U21 : OAI22_X1 port map( A1 => n163, A2 => n102, B1 => n158, B2 => n99, ZN 
                           => Y(22));
   U22 : OAI22_X1 port map( A1 => n164, A2 => n105, B1 => n158, B2 => n102, ZN 
                           => Y(21));
   U23 : OAI22_X1 port map( A1 => n164, A2 => n108, B1 => n158, B2 => n105, ZN 
                           => Y(20));
   U24 : OAI22_X1 port map( A1 => n164, A2 => n114, B1 => n158, B2 => n108, ZN 
                           => Y(19));
   U25 : OAI22_X1 port map( A1 => n165, A2 => n117, B1 => n158, B2 => n114, ZN 
                           => Y(18));
   U26 : OAI22_X1 port map( A1 => n165, A2 => n120, B1 => n158, B2 => n117, ZN 
                           => Y(17));
   U27 : OAI22_X1 port map( A1 => n165, A2 => n123, B1 => n158, B2 => n120, ZN 
                           => Y(16));
   U28 : OAI22_X1 port map( A1 => n159, A2 => n43, B1 => n158, B2 => n41, ZN =>
                           Y(8));
   U29 : OAI22_X1 port map( A1 => sel(0), A2 => n138, B1 => n159, B2 => n40, ZN
                           => Y(10));
   U30 : OAI221_X1 port map( B1 => A(13), B2 => n154, C1 => A(11), C2 => n44, A
                           => n142, ZN => n138);
   U31 : AOI22_X1 port map( A1 => n47, A2 => n50, B1 => n150, B2 => n137, ZN =>
                           n142);
   U32 : OAI221_X1 port map( B1 => A(20), B2 => n155, C1 => A(18), C2 => n156, 
                           A => n121, ZN => n117);
   U33 : AOI22_X1 port map( A1 => n152, A2 => n122, B1 => n150, B2 => n116, ZN 
                           => n121);
   U34 : OAI221_X1 port map( B1 => A(19), B2 => n154, C1 => A(17), C2 => n156, 
                           A => n124, ZN => n120);
   U35 : AOI22_X1 port map( A1 => n152, A2 => n125, B1 => n150, B2 => n119, ZN 
                           => n124);
   U36 : OAI221_X1 port map( B1 => A(18), B2 => n155, C1 => A(16), C2 => n156, 
                           A => n127, ZN => n123);
   U37 : AOI22_X1 port map( A1 => n152, A2 => n128, B1 => n150, B2 => n122, ZN 
                           => n127);
   U38 : OAI221_X1 port map( B1 => A(16), B2 => n154, C1 => A(14), C2 => n156, 
                           A => n133, ZN => n129);
   U39 : AOI22_X1 port map( A1 => n152, A2 => n134, B1 => n150, B2 => n128, ZN 
                           => n133);
   U40 : OAI221_X1 port map( B1 => A(15), B2 => n155, C1 => A(13), C2 => n156, 
                           A => n136, ZN => n132);
   U41 : AOI22_X1 port map( A1 => n152, A2 => n137, B1 => n150, B2 => n131, ZN 
                           => n136);
   U42 : OAI221_X1 port map( B1 => A(14), B2 => n154, C1 => A(12), C2 => n156, 
                           A => n139, ZN => n135);
   U43 : AOI22_X1 port map( A1 => n152, A2 => n140, B1 => n150, B2 => n134, ZN 
                           => n139);
   U44 : OAI221_X1 port map( B1 => A(12), B2 => n154, C1 => A(10), C2 => n156, 
                           A => n141, ZN => n40);
   U45 : AOI22_X1 port map( A1 => n152, A2 => n54, B1 => n150, B2 => n140, ZN 
                           => n141);
   U46 : OAI221_X1 port map( B1 => A(8), B2 => n44, C1 => A(10), C2 => n154, A 
                           => n52, ZN => n43);
   U47 : AOI22_X1 port map( A1 => n152, A2 => n53, B1 => n49, B2 => n54, ZN => 
                           n52);
   U48 : OAI221_X1 port map( B1 => A(32), B2 => n154, C1 => A(30), C2 => n156, 
                           A => n84, ZN => n74);
   U49 : AOI22_X1 port map( A1 => n152, A2 => n72, B1 => n49, B2 => n85, ZN => 
                           n84);
   U50 : INV_X1 port map( A => A(36), ZN => n85);
   U51 : OAI221_X1 port map( B1 => A(31), B2 => n155, C1 => A(29), C2 => n44, A
                           => n87, ZN => n83);
   U52 : AOI22_X1 port map( A1 => n152, A2 => n79, B1 => n49, B2 => n88, ZN => 
                           n87);
   U53 : INV_X1 port map( A => A(35), ZN => n88);
   U54 : OAI221_X1 port map( B1 => A(30), B2 => n155, C1 => A(28), C2 => n156, 
                           A => n90, ZN => n86);
   U55 : AOI22_X1 port map( A1 => n47, A2 => n73, B1 => n49, B2 => n72, ZN => 
                           n90);
   U56 : OAI221_X1 port map( B1 => A(29), B2 => n155, C1 => A(27), C2 => n44, A
                           => n92, ZN => n89);
   U57 : AOI22_X1 port map( A1 => n47, A2 => n77, B1 => n49, B2 => n79, ZN => 
                           n92);
   U58 : OAI221_X1 port map( B1 => A(28), B2 => n155, C1 => A(26), C2 => n156, 
                           A => n94, ZN => n91);
   U59 : AOI22_X1 port map( A1 => n47, A2 => n95, B1 => n49, B2 => n73, ZN => 
                           n94);
   U60 : OAI221_X1 port map( B1 => A(27), B2 => n155, C1 => A(25), C2 => n44, A
                           => n97, ZN => n93);
   U61 : AOI22_X1 port map( A1 => n47, A2 => n98, B1 => n49, B2 => n77, ZN => 
                           n97);
   U62 : OAI221_X1 port map( B1 => A(26), B2 => n155, C1 => A(24), C2 => n156, 
                           A => n100, ZN => n96);
   U63 : AOI22_X1 port map( A1 => n47, A2 => n101, B1 => n49, B2 => n95, ZN => 
                           n100);
   U64 : OAI221_X1 port map( B1 => A(25), B2 => n155, C1 => A(23), C2 => n44, A
                           => n103, ZN => n99);
   U65 : AOI22_X1 port map( A1 => n47, A2 => n104, B1 => n150, B2 => n98, ZN =>
                           n103);
   U66 : OAI221_X1 port map( B1 => A(24), B2 => n155, C1 => A(22), C2 => n156, 
                           A => n106, ZN => n102);
   U67 : AOI22_X1 port map( A1 => n47, A2 => n107, B1 => n150, B2 => n101, ZN 
                           => n106);
   U68 : OAI221_X1 port map( B1 => A(23), B2 => n155, C1 => A(21), C2 => n156, 
                           A => n109, ZN => n105);
   U69 : AOI22_X1 port map( A1 => n152, A2 => n110, B1 => n150, B2 => n104, ZN 
                           => n109);
   U70 : OAI221_X1 port map( B1 => A(22), B2 => n155, C1 => A(20), C2 => n156, 
                           A => n115, ZN => n108);
   U71 : AOI22_X1 port map( A1 => n152, A2 => n116, B1 => n150, B2 => n107, ZN 
                           => n115);
   U72 : OAI221_X1 port map( B1 => A(21), B2 => n155, C1 => A(19), C2 => n156, 
                           A => n118, ZN => n114);
   U73 : AOI22_X1 port map( A1 => n152, A2 => n119, B1 => n150, B2 => n110, ZN 
                           => n118);
   U74 : OAI221_X1 port map( B1 => A(17), B2 => n155, C1 => A(15), C2 => n156, 
                           A => n130, ZN => n126);
   U75 : AOI22_X1 port map( A1 => n152, A2 => n131, B1 => n150, B2 => n125, ZN 
                           => n130);
   U76 : OAI221_X1 port map( B1 => A(9), B2 => n44, C1 => A(11), C2 => n154, A 
                           => n46, ZN => n41);
   U77 : AOI22_X1 port map( A1 => n152, A2 => n48, B1 => n150, B2 => n50, ZN =>
                           n46);
   U78 : OAI22_X1 port map( A1 => n163, A2 => n74, B1 => n158, B2 => n69, ZN =>
                           Y(30));
   U79 : OAI22_X1 port map( A1 => n160, A2 => n51, B1 => n158, B2 => n43, ZN =>
                           Y(7));
   U80 : OAI22_X1 port map( A1 => n160, A2 => n55, B1 => n158, B2 => n51, ZN =>
                           Y(6));
   U81 : OAI22_X1 port map( A1 => n160, A2 => n58, B1 => n158, B2 => n55, ZN =>
                           Y(5));
   U82 : OAI22_X1 port map( A1 => n160, A2 => n61, B1 => n158, B2 => n58, ZN =>
                           Y(4));
   U83 : OAI22_X1 port map( A1 => n161, A2 => n66, B1 => sel(0), B2 => n61, ZN 
                           => Y(3));
   U84 : OAI22_X1 port map( A1 => n161, A2 => n80, B1 => sel(0), B2 => n66, ZN 
                           => Y(2));
   U85 : OAI22_X1 port map( A1 => n164, A2 => n111, B1 => n158, B2 => n80, ZN 
                           => Y(1));
   U86 : BUF_X1 port map( A => n167, Z => n160);
   U87 : BUF_X1 port map( A => n167, Z => n161);
   U88 : BUF_X1 port map( A => n165, Z => n162);
   U89 : INV_X1 port map( A => A(31), ZN => n77);
   U90 : INV_X1 port map( A => A(32), ZN => n73);
   U91 : BUF_X1 port map( A => n167, Z => n159);
   U92 : BUF_X1 port map( A => n166, Z => n163);
   U93 : BUF_X1 port map( A => n167, Z => n165);
   U94 : BUF_X1 port map( A => n167, Z => n166);
   U95 : BUF_X1 port map( A => n167, Z => n164);
   U96 : INV_X1 port map( A => A(30), ZN => n95);
   U97 : INV_X1 port map( A => A(29), ZN => n98);
   U98 : INV_X1 port map( A => A(28), ZN => n101);
   U99 : INV_X1 port map( A => A(27), ZN => n104);
   U100 : INV_X1 port map( A => A(26), ZN => n107);
   U101 : INV_X1 port map( A => A(25), ZN => n110);
   U102 : INV_X1 port map( A => A(24), ZN => n116);
   U103 : INV_X1 port map( A => A(23), ZN => n119);
   U104 : INV_X1 port map( A => A(22), ZN => n122);
   U105 : INV_X1 port map( A => A(21), ZN => n125);
   U106 : INV_X1 port map( A => A(20), ZN => n128);
   U107 : INV_X1 port map( A => A(19), ZN => n131);
   U108 : INV_X1 port map( A => A(18), ZN => n134);
   U109 : INV_X1 port map( A => A(17), ZN => n137);
   U110 : INV_X1 port map( A => A(16), ZN => n140);
   U111 : INV_X1 port map( A => A(15), ZN => n50);
   U112 : INV_X1 port map( A => A(14), ZN => n54);
   U113 : INV_X1 port map( A => A(13), ZN => n48);
   U114 : INV_X1 port map( A => A(12), ZN => n53);
   U115 : OAI221_X1 port map( B1 => A(1), B2 => n44, C1 => A(3), C2 => n154, A 
                           => n146, ZN => n111);
   U116 : INV_X1 port map( A => n147, ZN => n146);
   U117 : OAI22_X1 port map( A1 => n153, A2 => A(5), B1 => n151, B2 => A(7), ZN
                           => n147);
   U118 : OAI221_X1 port map( B1 => A(3), B2 => n44, C1 => A(5), C2 => n154, A 
                           => n81, ZN => n66);
   U119 : INV_X1 port map( A => n82, ZN => n81);
   U120 : OAI22_X1 port map( A1 => n153, A2 => A(7), B1 => n151, B2 => A(9), ZN
                           => n82);
   U121 : OAI221_X1 port map( B1 => A(2), B2 => n44, C1 => A(4), C2 => n154, A 
                           => n112, ZN => n80);
   U122 : INV_X1 port map( A => n113, ZN => n112);
   U123 : OAI22_X1 port map( A1 => n153, A2 => A(6), B1 => n151, B2 => A(8), ZN
                           => n113);
   U124 : OAI221_X1 port map( B1 => A(9), B2 => n154, C1 => A(7), C2 => n44, A 
                           => n56, ZN => n51);
   U125 : AOI22_X1 port map( A1 => n47, A2 => n57, B1 => n49, B2 => n48, ZN => 
                           n56);
   U126 : INV_X1 port map( A => A(11), ZN => n57);
   U127 : OAI221_X1 port map( B1 => A(8), B2 => n154, C1 => A(6), C2 => n44, A 
                           => n59, ZN => n55);
   U128 : AOI22_X1 port map( A1 => n152, A2 => n60, B1 => n150, B2 => n53, ZN 
                           => n59);
   U129 : INV_X1 port map( A => A(10), ZN => n60);
   U130 : OAI221_X1 port map( B1 => A(7), B2 => n154, C1 => A(5), C2 => n44, A 
                           => n62, ZN => n58);
   U131 : INV_X1 port map( A => n63, ZN => n62);
   U132 : OAI22_X1 port map( A1 => n153, A2 => A(9), B1 => n151, B2 => A(11), 
                           ZN => n63);
   U133 : OAI221_X1 port map( B1 => A(6), B2 => n154, C1 => A(4), C2 => n44, A 
                           => n67, ZN => n61);
   U134 : INV_X1 port map( A => n68, ZN => n67);
   U135 : OAI22_X1 port map( A1 => n153, A2 => A(8), B1 => n151, B2 => A(10), 
                           ZN => n68);
   U136 : OAI221_X1 port map( B1 => A(35), B2 => n153, C1 => A(37), C2 => n151,
                           A => n75, ZN => n69);
   U137 : AOI22_X1 port map( A1 => n157, A2 => n77, B1 => n149, B2 => n79, ZN 
                           => n75);
   U138 : OAI22_X1 port map( A1 => n161, A2 => n69, B1 => n158, B2 => n70, ZN 
                           => Y(31));
   U139 : AOI221_X1 port map( B1 => A(36), B2 => n47, C1 => A(38), C2 => n49, A
                           => n71, ZN => n70);
   U140 : OAI22_X1 port map( A1 => n154, A2 => n72, B1 => n44, B2 => n73, ZN =>
                           n71);
   U141 : OAI22_X1 port map( A1 => sel(0), A2 => n111, B1 => n143, B2 => n159, 
                           ZN => Y(0));
   U142 : AOI221_X1 port map( B1 => A(0), B2 => n157, C1 => A(2), C2 => n149, A
                           => n144, ZN => n143);
   U143 : INV_X1 port map( A => n145, ZN => n144);
   U144 : NOR2_X1 port map( A1 => sel(1), A2 => sel(2), ZN => n49);
   U145 : NOR2_X1 port map( A1 => n148, A2 => sel(2), ZN => n47);
   U146 : AOI22_X1 port map( A1 => n49, A2 => A(6), B1 => n47, B2 => A(4), ZN 
                           => n145);
   U147 : NAND2_X1 port map( A1 => sel(2), A2 => sel(1), ZN => n44);
   U148 : INV_X1 port map( A => A(33), ZN => n79);
   U149 : INV_X1 port map( A => A(34), ZN => n72);
   U150 : INV_X1 port map( A => sel(1), ZN => n148);
   U151 : INV_X1 port map( A => sel(0), ZN => n167);
   U152 : INV_X1 port map( A => n49, ZN => n151);
   U153 : INV_X1 port map( A => n47, ZN => n153);
   U154 : INV_X1 port map( A => n44, ZN => n157);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_secondLevel is

   port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : in 
         std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 downto 
         0));

end shift_secondLevel;

architecture SYN_behav of shift_secondLevel is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
      n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n90, Z => n93);
   U3 : BUF_X1 port map( A => n91, Z => n94);
   U4 : BUF_X1 port map( A => n90, Z => n92);
   U5 : BUF_X1 port map( A => n84, Z => n87);
   U6 : BUF_X1 port map( A => n85, Z => n88);
   U7 : BUF_X1 port map( A => n84, Z => n86);
   U8 : BUF_X1 port map( A => n96, Z => n99);
   U9 : BUF_X1 port map( A => n97, Z => n100);
   U10 : BUF_X1 port map( A => n96, Z => n98);
   U11 : BUF_X1 port map( A => n91, Z => n95);
   U12 : BUF_X1 port map( A => n85, Z => n89);
   U13 : BUF_X1 port map( A => n97, Z => n101);
   U14 : INV_X1 port map( A => n71, ZN => Y(1));
   U15 : INV_X1 port map( A => n52, ZN => Y(37));
   U16 : AOI222_X1 port map( A1 => mask00(37), A2 => n100, B1 => mask16(37), B2
                           => n94, C1 => mask08(37), C2 => n88, ZN => n52);
   U17 : INV_X1 port map( A => n51, ZN => Y(38));
   U18 : INV_X1 port map( A => n82, ZN => Y(0));
   U19 : INV_X1 port map( A => n41, ZN => Y(9));
   U20 : AOI222_X1 port map( A1 => mask00(9), A2 => n101, B1 => mask16(9), B2 
                           => n95, C1 => mask08(9), C2 => n89, ZN => n41);
   U21 : INV_X1 port map( A => n45, ZN => Y(8));
   U22 : AOI222_X1 port map( A1 => mask00(8), A2 => n101, B1 => mask16(8), B2 
                           => n95, C1 => mask08(8), C2 => n89, ZN => n45);
   U23 : INV_X1 port map( A => n80, ZN => Y(11));
   U24 : AOI222_X1 port map( A1 => mask00(11), A2 => n98, B1 => mask16(11), B2 
                           => n92, C1 => mask08(11), C2 => n86, ZN => n80);
   U25 : INV_X1 port map( A => n81, ZN => Y(10));
   U26 : AOI222_X1 port map( A1 => mask00(10), A2 => n98, B1 => mask16(10), B2 
                           => n92, C1 => mask08(10), C2 => n86, ZN => n81);
   U27 : INV_X1 port map( A => n59, ZN => Y(30));
   U28 : AOI222_X1 port map( A1 => mask00(30), A2 => n99, B1 => mask16(30), B2 
                           => n93, C1 => mask08(30), C2 => n87, ZN => n59);
   U29 : INV_X1 port map( A => n61, ZN => Y(29));
   U30 : AOI222_X1 port map( A1 => mask00(29), A2 => n99, B1 => mask16(29), B2 
                           => n93, C1 => mask08(29), C2 => n87, ZN => n61);
   U31 : INV_X1 port map( A => n62, ZN => Y(28));
   U32 : AOI222_X1 port map( A1 => mask00(28), A2 => n99, B1 => mask16(28), B2 
                           => n93, C1 => mask08(28), C2 => n87, ZN => n62);
   U33 : INV_X1 port map( A => n63, ZN => Y(27));
   U34 : AOI222_X1 port map( A1 => mask00(27), A2 => n99, B1 => mask16(27), B2 
                           => n93, C1 => mask08(27), C2 => n87, ZN => n63);
   U35 : INV_X1 port map( A => n64, ZN => Y(26));
   U36 : AOI222_X1 port map( A1 => mask00(26), A2 => n99, B1 => mask16(26), B2 
                           => n93, C1 => mask08(26), C2 => n87, ZN => n64);
   U37 : INV_X1 port map( A => n65, ZN => Y(25));
   U38 : AOI222_X1 port map( A1 => mask00(25), A2 => n99, B1 => mask16(25), B2 
                           => n93, C1 => mask08(25), C2 => n87, ZN => n65);
   U39 : INV_X1 port map( A => n66, ZN => Y(24));
   U40 : AOI222_X1 port map( A1 => mask00(24), A2 => n99, B1 => mask16(24), B2 
                           => n93, C1 => mask08(24), C2 => n87, ZN => n66);
   U41 : INV_X1 port map( A => n67, ZN => Y(23));
   U42 : AOI222_X1 port map( A1 => mask00(23), A2 => n99, B1 => mask16(23), B2 
                           => n93, C1 => mask08(23), C2 => n87, ZN => n67);
   U43 : INV_X1 port map( A => n68, ZN => Y(22));
   U44 : AOI222_X1 port map( A1 => mask00(22), A2 => n99, B1 => mask16(22), B2 
                           => n93, C1 => mask08(22), C2 => n87, ZN => n68);
   U45 : INV_X1 port map( A => n69, ZN => Y(21));
   U46 : AOI222_X1 port map( A1 => mask00(21), A2 => n99, B1 => mask16(21), B2 
                           => n93, C1 => mask08(21), C2 => n87, ZN => n69);
   U47 : INV_X1 port map( A => n70, ZN => Y(20));
   U48 : AOI222_X1 port map( A1 => mask00(20), A2 => n99, B1 => mask16(20), B2 
                           => n93, C1 => mask08(20), C2 => n87, ZN => n70);
   U49 : INV_X1 port map( A => n72, ZN => Y(19));
   U50 : AOI222_X1 port map( A1 => mask00(19), A2 => n98, B1 => mask16(19), B2 
                           => n92, C1 => mask08(19), C2 => n86, ZN => n72);
   U51 : INV_X1 port map( A => n73, ZN => Y(18));
   U52 : AOI222_X1 port map( A1 => mask00(18), A2 => n98, B1 => mask16(18), B2 
                           => n92, C1 => mask08(18), C2 => n86, ZN => n73);
   U53 : INV_X1 port map( A => n74, ZN => Y(17));
   U54 : AOI222_X1 port map( A1 => mask00(17), A2 => n98, B1 => mask16(17), B2 
                           => n92, C1 => mask08(17), C2 => n86, ZN => n74);
   U55 : INV_X1 port map( A => n75, ZN => Y(16));
   U56 : AOI222_X1 port map( A1 => mask00(16), A2 => n98, B1 => mask16(16), B2 
                           => n92, C1 => mask08(16), C2 => n86, ZN => n75);
   U57 : INV_X1 port map( A => n76, ZN => Y(15));
   U58 : AOI222_X1 port map( A1 => mask00(15), A2 => n98, B1 => mask16(15), B2 
                           => n92, C1 => mask08(15), C2 => n86, ZN => n76);
   U59 : INV_X1 port map( A => n77, ZN => Y(14));
   U60 : AOI222_X1 port map( A1 => mask00(14), A2 => n98, B1 => mask16(14), B2 
                           => n92, C1 => mask08(14), C2 => n86, ZN => n77);
   U61 : INV_X1 port map( A => n78, ZN => Y(13));
   U62 : AOI222_X1 port map( A1 => mask00(13), A2 => n98, B1 => mask16(13), B2 
                           => n92, C1 => mask08(13), C2 => n86, ZN => n78);
   U63 : INV_X1 port map( A => n79, ZN => Y(12));
   U64 : AOI222_X1 port map( A1 => mask00(12), A2 => n98, B1 => mask16(12), B2 
                           => n92, C1 => mask08(12), C2 => n86, ZN => n79);
   U65 : INV_X1 port map( A => n56, ZN => Y(33));
   U66 : AOI222_X1 port map( A1 => mask00(33), A2 => n100, B1 => mask16(33), B2
                           => n94, C1 => mask08(33), C2 => n88, ZN => n56);
   U67 : INV_X1 port map( A => n55, ZN => Y(34));
   U68 : AOI222_X1 port map( A1 => mask00(34), A2 => n100, B1 => mask16(34), B2
                           => n94, C1 => mask08(34), C2 => n88, ZN => n55);
   U69 : INV_X1 port map( A => n54, ZN => Y(35));
   U70 : AOI222_X1 port map( A1 => mask00(35), A2 => n100, B1 => mask16(35), B2
                           => n94, C1 => mask08(35), C2 => n88, ZN => n54);
   U71 : INV_X1 port map( A => n57, ZN => Y(32));
   U72 : AOI222_X1 port map( A1 => mask00(32), A2 => n100, B1 => mask16(32), B2
                           => n94, C1 => mask08(32), C2 => n88, ZN => n57);
   U73 : INV_X1 port map( A => n58, ZN => Y(31));
   U74 : AOI222_X1 port map( A1 => mask00(31), A2 => n100, B1 => mask16(31), B2
                           => n94, C1 => mask08(31), C2 => n88, ZN => n58);
   U75 : INV_X1 port map( A => n53, ZN => Y(36));
   U76 : AOI222_X1 port map( A1 => mask00(36), A2 => n100, B1 => mask16(36), B2
                           => n94, C1 => mask08(36), C2 => n88, ZN => n53);
   U77 : BUF_X1 port map( A => n42, Z => n96);
   U78 : BUF_X1 port map( A => n43, Z => n90);
   U79 : BUF_X1 port map( A => n44, Z => n84);
   U80 : BUF_X1 port map( A => n42, Z => n97);
   U81 : BUF_X1 port map( A => n43, Z => n91);
   U82 : BUF_X1 port map( A => n44, Z => n85);
   U83 : AOI222_X1 port map( A1 => mask00(38), A2 => n100, B1 => mask16(38), B2
                           => n94, C1 => mask08(38), C2 => n88, ZN => n51);
   U84 : AOI222_X1 port map( A1 => mask00(1), A2 => n98, B1 => mask16(1), B2 =>
                           n92, C1 => mask08(1), C2 => n86, ZN => n71);
   U85 : AOI222_X1 port map( A1 => mask00(0), A2 => n98, B1 => mask16(0), B2 =>
                           n92, C1 => mask08(0), C2 => n86, ZN => n82);
   U86 : INV_X1 port map( A => n47, ZN => Y(6));
   U87 : AOI222_X1 port map( A1 => mask00(6), A2 => n100, B1 => mask16(6), B2 
                           => n94, C1 => mask08(6), C2 => n88, ZN => n47);
   U88 : INV_X1 port map( A => n46, ZN => Y(7));
   U89 : AOI222_X1 port map( A1 => mask00(7), A2 => n101, B1 => mask16(7), B2 
                           => n95, C1 => mask08(7), C2 => n89, ZN => n46);
   U90 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n42);
   U91 : NOR2_X1 port map( A1 => n83, A2 => sel(0), ZN => n43);
   U92 : INV_X1 port map( A => n49, ZN => Y(4));
   U93 : AOI222_X1 port map( A1 => mask00(4), A2 => n100, B1 => mask16(4), B2 
                           => n94, C1 => mask08(4), C2 => n88, ZN => n49);
   U94 : INV_X1 port map( A => n48, ZN => Y(5));
   U95 : AOI222_X1 port map( A1 => mask00(5), A2 => n100, B1 => mask16(5), B2 
                           => n94, C1 => mask08(5), C2 => n88, ZN => n48);
   U96 : INV_X1 port map( A => n60, ZN => Y(2));
   U97 : AOI222_X1 port map( A1 => mask00(2), A2 => n99, B1 => mask16(2), B2 =>
                           n93, C1 => mask08(2), C2 => n87, ZN => n60);
   U98 : INV_X1 port map( A => n50, ZN => Y(3));
   U99 : AOI222_X1 port map( A1 => mask00(3), A2 => n100, B1 => mask16(3), B2 
                           => n94, C1 => mask08(3), C2 => n88, ZN => n50);
   U100 : INV_X1 port map( A => sel(1), ZN => n83);
   U101 : AND2_X1 port map( A1 => sel(0), A2 => n83, ZN => n44);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_firstLevel is

   port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector (1 
         downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 downto 
         0));

end shift_firstLevel;

architecture SYN_behav of shift_firstLevel is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask08_23_port, mask08_22_port, mask08_21_port, mask08_20_port, 
      mask08_19_port, mask08_18_port, mask08_17_port, mask08_16_port, 
      mask08_15_port, mask08_7_port, mask08_6_port, mask08_5_port, 
      mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port, mask08_0_port
      , mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n98, n116, n117, mask16_22_port, n119, n120, n121 : std_logic
      ;

begin
   mask08 <= ( mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask08_23_port, 
      mask08_22_port, mask08_21_port, mask08_20_port, mask08_19_port, 
      mask08_18_port, mask08_17_port, mask08_16_port, mask08_15_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port, mask08_7_port, mask08_6_port, 
      mask08_5_port, mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port
      , mask08_0_port );
   mask16 <= ( mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_22_port, mask16_22_port, mask16_22_port, mask16_22_port, 
      mask16_22_port, mask16_22_port, mask16_22_port, mask16_15_port, 
      mask16_14_port, mask16_13_port, mask16_12_port, mask16_11_port, 
      mask16_10_port, mask16_9_port, mask16_8_port, mask16_7_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port );
   
   U161 : NAND3_X1 port map( A1 => sel(1), A2 => n108, A3 => A(31), ZN => n61);
   U2 : INV_X1 port map( A => n116, ZN => n98);
   U3 : INV_X1 port map( A => mask16_22_port, ZN => n117);
   U4 : BUF_X1 port map( A => n59, Z => n121);
   U5 : BUF_X1 port map( A => n59, Z => n120);
   U6 : BUF_X1 port map( A => n59, Z => n119);
   U7 : INV_X1 port map( A => mask16_7_port, ZN => n94);
   U8 : INV_X1 port map( A => mask08_6_port, ZN => n111);
   U9 : INV_X1 port map( A => mask08_1_port, ZN => n96);
   U10 : INV_X1 port map( A => mask08_5_port, ZN => n112);
   U11 : INV_X1 port map( A => mask08_4_port, ZN => n113);
   U12 : INV_X1 port map( A => mask08_3_port, ZN => n114);
   U13 : INV_X1 port map( A => mask08_2_port, ZN => n115);
   U14 : OAI21_X1 port map( B1 => n120, B2 => n60, A => n117, ZN => 
                           mask16_38_port);
   U15 : OAI21_X1 port map( B1 => n120, B2 => n63, A => n117, ZN => 
                           mask16_36_port);
   U16 : OAI21_X1 port map( B1 => n120, B2 => n64, A => n117, ZN => 
                           mask16_35_port);
   U17 : OAI21_X1 port map( B1 => n120, B2 => n65, A => n117, ZN => 
                           mask16_34_port);
   U18 : OAI21_X1 port map( B1 => n120, B2 => n66, A => n117, ZN => 
                           mask16_33_port);
   U19 : OAI21_X1 port map( B1 => n120, B2 => n67, A => n117, ZN => 
                           mask16_32_port);
   U20 : OAI21_X1 port map( B1 => n120, B2 => n62, A => n117, ZN => 
                           mask16_37_port);
   U21 : NOR2_X1 port map( A1 => n86, A2 => n116, ZN => mask16_7_port);
   U22 : NOR2_X1 port map( A1 => n60, A2 => n116, ZN => mask08_7_port);
   U23 : NOR2_X1 port map( A1 => n62, A2 => n116, ZN => mask08_6_port);
   U24 : NOR2_X1 port map( A1 => n67, A2 => n116, ZN => mask08_1_port);
   U25 : NOR2_X1 port map( A1 => n65, A2 => n116, ZN => mask08_3_port);
   U26 : NOR2_X1 port map( A1 => n66, A2 => n116, ZN => mask08_2_port);
   U27 : NOR2_X1 port map( A1 => n63, A2 => n116, ZN => mask08_5_port);
   U28 : NOR2_X1 port map( A1 => n64, A2 => n116, ZN => mask08_4_port);
   U29 : INV_X1 port map( A => n61, ZN => mask16_22_port);
   U30 : INV_X1 port map( A => n53, ZN => mask16_9_port);
   U31 : NAND2_X1 port map( A1 => n96, A2 => n75, ZN => mask00(9));
   U32 : INV_X1 port map( A => n54, ZN => mask16_8_port);
   U33 : NAND2_X1 port map( A1 => n95, A2 => n76, ZN => mask00(8));
   U34 : INV_X1 port map( A => n83, ZN => mask16_11_port);
   U35 : NAND2_X1 port map( A1 => n114, A2 => n73, ZN => mask00(11));
   U36 : INV_X1 port map( A => n84, ZN => mask16_10_port);
   U37 : NAND2_X1 port map( A1 => n115, A2 => n74, ZN => mask00(10));
   U38 : OAI21_X1 port map( B1 => n121, B2 => n93, A => n94, ZN => mask00(23));
   U39 : OAI21_X1 port map( B1 => n87, B2 => n119, A => n117, ZN => 
                           mask08_37_port);
   U40 : INV_X1 port map( A => n97, ZN => n59);
   U41 : NAND2_X1 port map( A1 => n61, A2 => n69, ZN => mask16_30_port);
   U42 : OAI21_X1 port map( B1 => n86, B2 => n119, A => n80, ZN => mask00(30));
   U43 : NAND2_X1 port map( A1 => n61, A2 => n71, ZN => mask16_29_port);
   U44 : OAI21_X1 port map( B1 => n87, B2 => n119, A => n81, ZN => mask00(29));
   U45 : NAND2_X1 port map( A1 => n61, A2 => n72, ZN => mask16_28_port);
   U46 : OAI21_X1 port map( B1 => n88, B2 => n119, A => n82, ZN => mask00(28));
   U47 : NAND2_X1 port map( A1 => n61, A2 => n73, ZN => mask16_27_port);
   U48 : OAI21_X1 port map( B1 => n89, B2 => n119, A => n83, ZN => mask00(27));
   U49 : NAND2_X1 port map( A1 => n61, A2 => n74, ZN => mask16_26_port);
   U50 : OAI21_X1 port map( B1 => n90, B2 => n119, A => n84, ZN => mask00(26));
   U51 : NAND2_X1 port map( A1 => n61, A2 => n75, ZN => mask16_25_port);
   U52 : OAI21_X1 port map( B1 => n121, B2 => n91, A => n53, ZN => mask00(25));
   U53 : NAND2_X1 port map( A1 => n117, A2 => n76, ZN => mask16_24_port);
   U54 : OAI21_X1 port map( B1 => n121, B2 => n92, A => n54, ZN => mask00(24));
   U55 : NAND2_X1 port map( A1 => n79, A2 => n68, ZN => mask08_23_port);
   U56 : NAND2_X1 port map( A1 => n61, A2 => n77, ZN => mask16_23_port);
   U57 : NAND2_X1 port map( A1 => n80, A2 => n69, ZN => mask08_22_port);
   U58 : OAI21_X1 port map( B1 => n121, B2 => n60, A => n55, ZN => mask00(22));
   U59 : NAND2_X1 port map( A1 => n81, A2 => n71, ZN => mask08_21_port);
   U60 : OAI21_X1 port map( B1 => n121, B2 => n62, A => n56, ZN => mask00(21));
   U61 : NAND2_X1 port map( A1 => n82, A2 => n72, ZN => mask08_20_port);
   U62 : OAI21_X1 port map( B1 => n121, B2 => n63, A => n57, ZN => mask00(20));
   U63 : NAND2_X1 port map( A1 => n83, A2 => n73, ZN => mask08_19_port);
   U64 : OAI21_X1 port map( B1 => n121, B2 => n64, A => n58, ZN => mask00(19));
   U65 : NAND2_X1 port map( A1 => n84, A2 => n74, ZN => mask08_18_port);
   U66 : OAI21_X1 port map( B1 => n121, B2 => n65, A => n70, ZN => mask00(18));
   U67 : NAND2_X1 port map( A1 => n53, A2 => n75, ZN => mask08_17_port);
   U68 : OAI21_X1 port map( B1 => n121, B2 => n66, A => n78, ZN => mask00(17));
   U69 : NAND2_X1 port map( A1 => n54, A2 => n76, ZN => mask08_16_port);
   U70 : OAI21_X1 port map( B1 => n120, B2 => n67, A => n85, ZN => mask00(16));
   U71 : INV_X1 port map( A => n79, ZN => mask16_15_port);
   U72 : NAND2_X1 port map( A1 => n94, A2 => n77, ZN => mask08_15_port);
   U73 : INV_X1 port map( A => n80, ZN => mask16_14_port);
   U74 : NAND2_X1 port map( A1 => n111, A2 => n69, ZN => mask00(14));
   U75 : INV_X1 port map( A => n81, ZN => mask16_13_port);
   U76 : NAND2_X1 port map( A1 => n112, A2 => n71, ZN => mask00(13));
   U77 : INV_X1 port map( A => n82, ZN => mask16_12_port);
   U78 : NAND2_X1 port map( A1 => n113, A2 => n72, ZN => mask00(12));
   U79 : OAI21_X1 port map( B1 => n120, B2 => n91, A => n61, ZN => 
                           mask08_33_port);
   U80 : OAI21_X1 port map( B1 => n90, B2 => n119, A => n117, ZN => 
                           mask08_34_port);
   U81 : OAI21_X1 port map( B1 => n89, B2 => n119, A => n117, ZN => 
                           mask08_35_port);
   U82 : OAI21_X1 port map( B1 => n121, B2 => n104, A => n61, ZN => mask00(35))
                           ;
   U83 : OAI21_X1 port map( B1 => n120, B2 => n92, A => n117, ZN => 
                           mask08_32_port);
   U84 : OAI21_X1 port map( B1 => n107, B2 => n119, A => n117, ZN => mask00(32)
                           );
   U85 : NAND2_X1 port map( A1 => n61, A2 => n68, ZN => mask16_31_port);
   U86 : OAI21_X1 port map( B1 => n120, B2 => n93, A => n61, ZN => 
                           mask08_31_port);
   U87 : OAI21_X1 port map( B1 => n88, B2 => n119, A => n117, ZN => 
                           mask08_36_port);
   U88 : OAI21_X1 port map( B1 => n121, B2 => n103, A => n117, ZN => mask00(36)
                           );
   U89 : INV_X1 port map( A => n55, ZN => mask16_6_port);
   U90 : INV_X1 port map( A => n56, ZN => mask16_5_port);
   U91 : INV_X1 port map( A => n57, ZN => mask16_4_port);
   U92 : INV_X1 port map( A => n58, ZN => mask16_3_port);
   U93 : INV_X1 port map( A => n78, ZN => mask16_1_port);
   U94 : INV_X1 port map( A => n85, ZN => mask16_0_port);
   U95 : INV_X1 port map( A => n70, ZN => mask16_2_port);
   U96 : NAND2_X1 port map( A1 => n110, A2 => n68, ZN => mask00(15));
   U97 : INV_X1 port map( A => mask08_7_port, ZN => n110);
   U98 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n97);
   U99 : OAI21_X1 port map( B1 => n86, B2 => n119, A => n117, ZN => 
                           mask08_38_port);
   U100 : OAI21_X1 port map( B1 => n120, B2 => n101, A => n61, ZN => mask00(38)
                           );
   U101 : INV_X1 port map( A => A(31), ZN => n101);
   U102 : AND2_X1 port map( A1 => n99, A2 => A(1), ZN => mask00(1));
   U103 : INV_X1 port map( A => n95, ZN => mask08_0_port);
   U104 : AND2_X1 port map( A1 => n99, A2 => A(0), ZN => mask00(0));
   U105 : INV_X1 port map( A => sel(0), ZN => n108);
   U106 : AOI21_X1 port map( B1 => sel(0), B2 => sel(1), A => n97, ZN => n99);
   U107 : NAND2_X1 port map( A1 => A(8), A2 => n97, ZN => n68);
   U108 : NAND2_X1 port map( A1 => A(7), A2 => n97, ZN => n69);
   U109 : NAND2_X1 port map( A1 => A(2), A2 => n97, ZN => n75);
   U110 : NAND2_X1 port map( A1 => A(1), A2 => n97, ZN => n76);
   U111 : NAND2_X1 port map( A1 => A(6), A2 => n97, ZN => n71);
   U112 : NAND2_X1 port map( A1 => A(5), A2 => n97, ZN => n72);
   U113 : NAND2_X1 port map( A1 => A(4), A2 => n97, ZN => n73);
   U114 : NAND2_X1 port map( A1 => A(3), A2 => n97, ZN => n74);
   U115 : AND2_X1 port map( A1 => n99, A2 => A(6), ZN => mask00(6));
   U116 : NAND2_X1 port map( A1 => A(0), A2 => n97, ZN => n77);
   U117 : OAI21_X1 port map( B1 => n116, B2 => n100, A => n77, ZN => mask00(7))
                           ;
   U118 : INV_X1 port map( A => A(7), ZN => n100);
   U119 : NAND2_X1 port map( A1 => A(31), A2 => n98, ZN => n79);
   U120 : NAND2_X1 port map( A1 => A(30), A2 => n98, ZN => n80);
   U121 : NAND2_X1 port map( A1 => A(25), A2 => n98, ZN => n53);
   U122 : NAND2_X1 port map( A1 => A(24), A2 => n98, ZN => n54);
   U123 : NAND2_X1 port map( A1 => A(29), A2 => n98, ZN => n81);
   U124 : NAND2_X1 port map( A1 => A(28), A2 => n98, ZN => n82);
   U125 : NAND2_X1 port map( A1 => A(27), A2 => n98, ZN => n83);
   U126 : NAND2_X1 port map( A1 => A(26), A2 => n98, ZN => n84);
   U127 : OAI21_X1 port map( B1 => n109, B2 => n119, A => n79, ZN => mask00(31)
                           );
   U128 : INV_X1 port map( A => A(24), ZN => n109);
   U129 : OAI21_X1 port map( B1 => n121, B2 => n105, A => n61, ZN => mask00(34)
                           );
   U130 : INV_X1 port map( A => A(27), ZN => n105);
   U131 : OAI21_X1 port map( B1 => n121, B2 => n106, A => n61, ZN => mask00(33)
                           );
   U132 : INV_X1 port map( A => A(26), ZN => n106);
   U133 : OAI21_X1 port map( B1 => n120, B2 => n102, A => n61, ZN => mask00(37)
                           );
   U134 : INV_X1 port map( A => A(30), ZN => n102);
   U135 : NAND2_X1 port map( A1 => A(21), A2 => n98, ZN => n56);
   U136 : NAND2_X1 port map( A1 => A(20), A2 => n98, ZN => n57);
   U137 : NAND2_X1 port map( A1 => A(19), A2 => n98, ZN => n58);
   U138 : NAND2_X1 port map( A1 => A(22), A2 => n98, ZN => n55);
   U139 : AND2_X1 port map( A1 => n99, A2 => A(4), ZN => mask00(4));
   U140 : AND2_X1 port map( A1 => n99, A2 => A(5), ZN => mask00(5));
   U141 : INV_X1 port map( A => A(15), ZN => n60);
   U142 : INV_X1 port map( A => A(14), ZN => n62);
   U143 : INV_X1 port map( A => A(9), ZN => n67);
   U144 : INV_X1 port map( A => A(11), ZN => n65);
   U145 : INV_X1 port map( A => A(10), ZN => n66);
   U146 : INV_X1 port map( A => A(13), ZN => n63);
   U147 : INV_X1 port map( A => A(12), ZN => n64);
   U148 : INV_X1 port map( A => A(23), ZN => n86);
   U149 : NAND2_X1 port map( A1 => A(18), A2 => n99, ZN => n70);
   U150 : NAND2_X1 port map( A1 => A(17), A2 => n99, ZN => n78);
   U151 : NAND2_X1 port map( A1 => A(16), A2 => n99, ZN => n85);
   U152 : NAND2_X1 port map( A1 => A(8), A2 => n99, ZN => n95);
   U153 : AND2_X1 port map( A1 => n99, A2 => A(2), ZN => mask00(2));
   U154 : AND2_X1 port map( A1 => n99, A2 => A(3), ZN => mask00(3));
   U155 : INV_X1 port map( A => A(18), ZN => n91);
   U156 : INV_X1 port map( A => A(17), ZN => n92);
   U157 : INV_X1 port map( A => A(16), ZN => n93);
   U158 : INV_X1 port map( A => A(22), ZN => n87);
   U159 : INV_X1 port map( A => A(21), ZN => n88);
   U160 : INV_X1 port map( A => A(20), ZN => n89);
   U162 : INV_X1 port map( A => A(19), ZN => n90);
   U163 : INV_X1 port map( A => A(29), ZN => n103);
   U164 : INV_X1 port map( A => A(28), ZN => n104);
   U165 : INV_X1 port map( A => A(25), ZN => n107);
   U166 : INV_X1 port map( A => n99, ZN => n116);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_1;

architecture SYN_struct of CSA_Nbits32_1 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_96 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co 
                           => Cout(1));
   FullAdd_1 : FA_95 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co 
                           => Cout(2));
   FullAdd_2 : FA_94 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co 
                           => Cout(3));
   FullAdd_3 : FA_93 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co 
                           => Cout(4));
   FullAdd_4 : FA_92 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co 
                           => Cout(5));
   FullAdd_5 : FA_91 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co 
                           => Cout(6));
   FullAdd_6 : FA_90 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co 
                           => Cout(7));
   FullAdd_7 : FA_89 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co 
                           => Cout(8));
   FullAdd_8 : FA_88 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co 
                           => Cout(9));
   FullAdd_9 : FA_87 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co 
                           => Cout(10));
   FullAdd_10 : FA_86 port map( A => A(10), B => B(10), Ci => C(10), S => S(10)
                           , Co => Cout(11));
   FullAdd_11 : FA_85 port map( A => A(11), B => B(11), Ci => C(11), S => S(11)
                           , Co => Cout(12));
   FullAdd_12 : FA_84 port map( A => A(12), B => B(12), Ci => C(12), S => S(12)
                           , Co => Cout(13));
   FullAdd_13 : FA_83 port map( A => A(13), B => B(13), Ci => C(13), S => S(13)
                           , Co => Cout(14));
   FullAdd_14 : FA_82 port map( A => A(14), B => B(14), Ci => C(14), S => S(14)
                           , Co => Cout(15));
   FullAdd_15 : FA_81 port map( A => A(15), B => B(15), Ci => C(15), S => S(15)
                           , Co => Cout(16));
   FullAdd_16 : FA_80 port map( A => A(16), B => B(16), Ci => C(16), S => S(16)
                           , Co => Cout(17));
   FullAdd_17 : FA_79 port map( A => A(17), B => B(17), Ci => C(17), S => S(17)
                           , Co => Cout(18));
   FullAdd_18 : FA_78 port map( A => A(18), B => B(18), Ci => C(18), S => S(18)
                           , Co => Cout(19));
   FullAdd_19 : FA_77 port map( A => A(19), B => B(19), Ci => C(19), S => S(19)
                           , Co => Cout(20));
   FullAdd_20 : FA_76 port map( A => A(20), B => B(20), Ci => C(20), S => S(20)
                           , Co => Cout(21));
   FullAdd_21 : FA_75 port map( A => A(21), B => B(21), Ci => C(21), S => S(21)
                           , Co => Cout(22));
   FullAdd_22 : FA_74 port map( A => A(22), B => B(22), Ci => C(22), S => S(22)
                           , Co => Cout(23));
   FullAdd_23 : FA_73 port map( A => A(23), B => B(23), Ci => C(23), S => S(23)
                           , Co => Cout(24));
   FullAdd_24 : FA_72 port map( A => A(24), B => B(24), Ci => C(24), S => S(24)
                           , Co => Cout(25));
   FullAdd_25 : FA_71 port map( A => A(25), B => B(25), Ci => C(25), S => S(25)
                           , Co => Cout(26));
   FullAdd_26 : FA_70 port map( A => A(26), B => B(26), Ci => C(26), S => S(26)
                           , Co => Cout(27));
   FullAdd_27 : FA_69 port map( A => A(27), B => B(27), Ci => C(27), S => S(27)
                           , Co => Cout(28));
   FullAdd_28 : FA_68 port map( A => A(28), B => B(28), Ci => C(28), S => S(28)
                           , Co => Cout(29));
   FullAdd_29 : FA_67 port map( A => A(29), B => B(29), Ci => C(29), S => S(29)
                           , Co => Cout(30));
   FullAdd_30 : FA_66 port map( A => A(30), B => B(30), Ci => C(30), S => S(30)
                           , Co => Cout(31));
   LastFA : FA_65 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), Co
                           => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_2;

architecture SYN_struct of CSA_Nbits32_2 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_128 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_127 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_126 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_125 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_124 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_123 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_122 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_121 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_120 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_119 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_118 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_117 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_116 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_115 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_114 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_113 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_112 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_111 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_110 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_109 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_108 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_107 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_106 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_105 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_104 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_103 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_102 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_101 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_100 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_99 port map( A => A(29), B => B(29), Ci => C(29), S => S(29)
                           , Co => Cout(30));
   FullAdd_30 : FA_98 port map( A => A(30), B => B(30), Ci => C(30), S => S(30)
                           , Co => Cout(31));
   LastFA : FA_97 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), Co
                           => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_3;

architecture SYN_struct of CSA_Nbits32_3 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_160 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_159 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_158 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_157 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_156 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_155 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_154 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_153 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_152 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_151 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_150 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_149 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_148 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_147 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_146 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_145 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_144 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_143 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_142 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_141 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_140 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_139 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_138 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_137 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_136 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_135 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_134 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_133 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_132 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_131 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_130 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_129 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_4 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_4;

architecture SYN_struct of CSA_Nbits32_4 is

   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_192 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_191 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_190 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_189 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_188 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_187 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_186 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_185 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_184 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_183 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_182 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_181 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_180 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_179 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_178 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_177 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_176 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_175 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_174 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_173 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_172 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_171 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_170 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_169 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_168 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_167 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_166 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_165 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_164 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_163 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_162 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_161 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_5 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_5;

architecture SYN_struct of CSA_Nbits32_5 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_224 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co
                           => Cout(1));
   FullAdd_1 : FA_223 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_222 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_221 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_220 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_219 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_218 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_217 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_216 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_215 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_214 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_213 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_212 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_211 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_210 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_209 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_208 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_207 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_206 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_205 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_204 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_203 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_202 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_201 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_200 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_199 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_198 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_197 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_196 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_195 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_194 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_193 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity CSA_Nbits32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
         std_logic_vector (31 downto 0));

end CSA_Nbits32_0;

architecture SYN_struct of CSA_Nbits32_0 is

   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal net6198 : std_logic;

begin
   
   Cout(0) <= '0';
   FullAdd_0 : FA_64 port map( A => A(0), B => B(0), Ci => C(0), S => S(0), Co 
                           => Cout(1));
   FullAdd_1 : FA_255 port map( A => A(1), B => B(1), Ci => C(1), S => S(1), Co
                           => Cout(2));
   FullAdd_2 : FA_254 port map( A => A(2), B => B(2), Ci => C(2), S => S(2), Co
                           => Cout(3));
   FullAdd_3 : FA_253 port map( A => A(3), B => B(3), Ci => C(3), S => S(3), Co
                           => Cout(4));
   FullAdd_4 : FA_252 port map( A => A(4), B => B(4), Ci => C(4), S => S(4), Co
                           => Cout(5));
   FullAdd_5 : FA_251 port map( A => A(5), B => B(5), Ci => C(5), S => S(5), Co
                           => Cout(6));
   FullAdd_6 : FA_250 port map( A => A(6), B => B(6), Ci => C(6), S => S(6), Co
                           => Cout(7));
   FullAdd_7 : FA_249 port map( A => A(7), B => B(7), Ci => C(7), S => S(7), Co
                           => Cout(8));
   FullAdd_8 : FA_248 port map( A => A(8), B => B(8), Ci => C(8), S => S(8), Co
                           => Cout(9));
   FullAdd_9 : FA_247 port map( A => A(9), B => B(9), Ci => C(9), S => S(9), Co
                           => Cout(10));
   FullAdd_10 : FA_246 port map( A => A(10), B => B(10), Ci => C(10), S => 
                           S(10), Co => Cout(11));
   FullAdd_11 : FA_245 port map( A => A(11), B => B(11), Ci => C(11), S => 
                           S(11), Co => Cout(12));
   FullAdd_12 : FA_244 port map( A => A(12), B => B(12), Ci => C(12), S => 
                           S(12), Co => Cout(13));
   FullAdd_13 : FA_243 port map( A => A(13), B => B(13), Ci => C(13), S => 
                           S(13), Co => Cout(14));
   FullAdd_14 : FA_242 port map( A => A(14), B => B(14), Ci => C(14), S => 
                           S(14), Co => Cout(15));
   FullAdd_15 : FA_241 port map( A => A(15), B => B(15), Ci => C(15), S => 
                           S(15), Co => Cout(16));
   FullAdd_16 : FA_240 port map( A => A(16), B => B(16), Ci => C(16), S => 
                           S(16), Co => Cout(17));
   FullAdd_17 : FA_239 port map( A => A(17), B => B(17), Ci => C(17), S => 
                           S(17), Co => Cout(18));
   FullAdd_18 : FA_238 port map( A => A(18), B => B(18), Ci => C(18), S => 
                           S(18), Co => Cout(19));
   FullAdd_19 : FA_237 port map( A => A(19), B => B(19), Ci => C(19), S => 
                           S(19), Co => Cout(20));
   FullAdd_20 : FA_236 port map( A => A(20), B => B(20), Ci => C(20), S => 
                           S(20), Co => Cout(21));
   FullAdd_21 : FA_235 port map( A => A(21), B => B(21), Ci => C(21), S => 
                           S(21), Co => Cout(22));
   FullAdd_22 : FA_234 port map( A => A(22), B => B(22), Ci => C(22), S => 
                           S(22), Co => Cout(23));
   FullAdd_23 : FA_233 port map( A => A(23), B => B(23), Ci => C(23), S => 
                           S(23), Co => Cout(24));
   FullAdd_24 : FA_232 port map( A => A(24), B => B(24), Ci => C(24), S => 
                           S(24), Co => Cout(25));
   FullAdd_25 : FA_231 port map( A => A(25), B => B(25), Ci => C(25), S => 
                           S(25), Co => Cout(26));
   FullAdd_26 : FA_230 port map( A => A(26), B => B(26), Ci => C(26), S => 
                           S(26), Co => Cout(27));
   FullAdd_27 : FA_229 port map( A => A(27), B => B(27), Ci => C(27), S => 
                           S(27), Co => Cout(28));
   FullAdd_28 : FA_228 port map( A => A(28), B => B(28), Ci => C(28), S => 
                           S(28), Co => Cout(29));
   FullAdd_29 : FA_227 port map( A => A(29), B => B(29), Ci => C(29), S => 
                           S(29), Co => Cout(30));
   FullAdd_30 : FA_226 port map( A => A(30), B => B(30), Ci => C(30), S => 
                           S(30), Co => Cout(31));
   LastFA : FA_225 port map( A => A(31), B => B(31), Ci => C(31), S => S(31), 
                           Co => net6198);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_1 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_1;

architecture SYN_behav of mux_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n257);
   U2 : BUF_X1 port map( A => n10, Z => n256);
   U3 : BUF_X1 port map( A => n10, Z => n258);
   U4 : BUF_X1 port map( A => n6, Z => n269);
   U5 : BUF_X1 port map( A => n6, Z => n268);
   U6 : BUF_X1 port map( A => n9, Z => n260);
   U7 : BUF_X1 port map( A => n9, Z => n259);
   U8 : BUF_X1 port map( A => n7, Z => n266);
   U9 : BUF_X1 port map( A => n7, Z => n265);
   U10 : BUF_X1 port map( A => n8, Z => n263);
   U11 : BUF_X1 port map( A => n8, Z => n262);
   U12 : BUF_X1 port map( A => n9, Z => n261);
   U13 : BUF_X1 port map( A => n7, Z => n267);
   U14 : BUF_X1 port map( A => n8, Z => n264);
   U15 : BUF_X1 port map( A => n6, Z => n270);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U23 : AOI22_X1 port map( A1 => A(28), A2 => n260, B1 => B(28), B2 => n257, 
                           ZN => n31);
   U24 : AOI222_X1 port map( A1 => D(28), A2 => n269, B1 => E(28), B2 => n266, 
                           C1 => C(28), C2 => n263, ZN => n32);
   U25 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U26 : AOI22_X1 port map( A1 => A(14), A2 => n259, B1 => B(14), B2 => n256, 
                           ZN => n61);
   U27 : AOI222_X1 port map( A1 => D(14), A2 => n268, B1 => E(14), B2 => n265, 
                           C1 => C(14), C2 => n262, ZN => n62);
   U28 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U29 : AOI22_X1 port map( A1 => A(24), A2 => n260, B1 => B(24), B2 => n257, 
                           ZN => n39);
   U30 : AOI222_X1 port map( A1 => D(24), A2 => n269, B1 => E(24), B2 => n266, 
                           C1 => C(24), C2 => n263, ZN => n40);
   U31 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U32 : AOI22_X1 port map( A1 => A(18), A2 => n259, B1 => B(18), B2 => n256, 
                           ZN => n53);
   U33 : AOI222_X1 port map( A1 => D(18), A2 => n268, B1 => E(18), B2 => n265, 
                           C1 => C(18), C2 => n262, ZN => n54);
   U34 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n259, B1 => B(15), B2 => n256, 
                           ZN => n59);
   U36 : AOI222_X1 port map( A1 => D(15), A2 => n268, B1 => E(15), B2 => n265, 
                           C1 => C(15), C2 => n262, ZN => n60);
   U37 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U38 : AOI22_X1 port map( A1 => A(22), A2 => n260, B1 => B(22), B2 => n257, 
                           ZN => n43);
   U39 : AOI222_X1 port map( A1 => D(22), A2 => n269, B1 => E(22), B2 => n266, 
                           C1 => C(22), C2 => n263, ZN => n44);
   U40 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U41 : AOI22_X1 port map( A1 => A(16), A2 => n259, B1 => B(16), B2 => n256, 
                           ZN => n57);
   U42 : AOI222_X1 port map( A1 => D(16), A2 => n268, B1 => E(16), B2 => n265, 
                           C1 => C(16), C2 => n262, ZN => n58);
   U43 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U44 : AOI22_X1 port map( A1 => A(20), A2 => n260, B1 => B(20), B2 => n257, 
                           ZN => n47);
   U45 : AOI222_X1 port map( A1 => D(20), A2 => n269, B1 => E(20), B2 => n266, 
                           C1 => C(20), C2 => n263, ZN => n48);
   U46 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U47 : AOI22_X1 port map( A1 => A(27), A2 => n260, B1 => B(27), B2 => n257, 
                           ZN => n33);
   U48 : AOI222_X1 port map( A1 => D(27), A2 => n269, B1 => E(27), B2 => n266, 
                           C1 => C(27), C2 => n263, ZN => n34);
   U49 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U50 : AOI22_X1 port map( A1 => A(23), A2 => n260, B1 => B(23), B2 => n257, 
                           ZN => n41);
   U51 : AOI222_X1 port map( A1 => D(23), A2 => n269, B1 => E(23), B2 => n266, 
                           C1 => C(23), C2 => n263, ZN => n42);
   U52 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U53 : AOI22_X1 port map( A1 => A(17), A2 => n259, B1 => B(17), B2 => n256, 
                           ZN => n55);
   U54 : AOI222_X1 port map( A1 => D(17), A2 => n268, B1 => E(17), B2 => n265, 
                           C1 => C(17), C2 => n262, ZN => n56);
   U55 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U56 : AOI22_X1 port map( A1 => A(21), A2 => n260, B1 => B(21), B2 => n257, 
                           ZN => n45);
   U57 : AOI222_X1 port map( A1 => D(21), A2 => n269, B1 => E(21), B2 => n266, 
                           C1 => C(21), C2 => n263, ZN => n46);
   U58 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U59 : AOI22_X1 port map( A1 => A(19), A2 => n259, B1 => B(19), B2 => n256, 
                           ZN => n51);
   U60 : AOI222_X1 port map( A1 => D(19), A2 => n268, B1 => E(19), B2 => n265, 
                           C1 => C(19), C2 => n262, ZN => n52);
   U61 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U62 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U63 : AOI22_X1 port map( A1 => A(25), A2 => n260, B1 => B(25), B2 => n257, 
                           ZN => n37);
   U64 : AOI222_X1 port map( A1 => D(25), A2 => n269, B1 => E(25), B2 => n266, 
                           C1 => C(25), C2 => n263, ZN => n38);
   U65 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U66 : AOI22_X1 port map( A1 => A(29), A2 => n260, B1 => B(29), B2 => n257, 
                           ZN => n29);
   U67 : AOI222_X1 port map( A1 => D(29), A2 => n269, B1 => E(29), B2 => n266, 
                           C1 => C(29), C2 => n263, ZN => n30);
   U68 : INV_X1 port map( A => Sel(2), ZN => n74);
   U69 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U70 : AOI22_X1 port map( A1 => A(26), A2 => n260, B1 => B(26), B2 => n257, 
                           ZN => n35);
   U71 : AOI222_X1 port map( A1 => D(26), A2 => n269, B1 => E(26), B2 => n266, 
                           C1 => C(26), C2 => n263, ZN => n36);
   U72 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U73 : AOI22_X1 port map( A1 => A(6), A2 => n261, B1 => B(6), B2 => n258, ZN 
                           => n15);
   U74 : AOI222_X1 port map( A1 => D(6), A2 => n270, B1 => E(6), B2 => n267, C1
                           => C(6), C2 => n264, ZN => n16);
   U75 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U76 : AOI22_X1 port map( A1 => A(3), A2 => n261, B1 => B(3), B2 => n258, ZN 
                           => n21);
   U77 : AOI222_X1 port map( A1 => D(3), A2 => n270, B1 => E(3), B2 => n267, C1
                           => C(3), C2 => n264, ZN => n22);
   U78 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U79 : AOI22_X1 port map( A1 => A(7), A2 => n261, B1 => B(7), B2 => n258, ZN 
                           => n13);
   U80 : AOI222_X1 port map( A1 => D(7), A2 => n270, B1 => E(7), B2 => n267, C1
                           => C(7), C2 => n264, ZN => n14);
   U81 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U82 : AOI22_X1 port map( A1 => A(4), A2 => n261, B1 => B(4), B2 => n258, ZN 
                           => n19);
   U83 : AOI222_X1 port map( A1 => D(4), A2 => n270, B1 => E(4), B2 => n267, C1
                           => C(4), C2 => n264, ZN => n20);
   U84 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U85 : AOI22_X1 port map( A1 => A(8), A2 => n261, B1 => B(8), B2 => n258, ZN 
                           => n11);
   U86 : AOI222_X1 port map( A1 => D(8), A2 => n270, B1 => E(8), B2 => n267, C1
                           => C(8), C2 => n264, ZN => n12);
   U87 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U88 : AOI22_X1 port map( A1 => A(9), A2 => n261, B1 => B(9), B2 => n258, ZN 
                           => n4);
   U89 : AOI222_X1 port map( A1 => D(9), A2 => n270, B1 => E(9), B2 => n267, C1
                           => C(9), C2 => n264, ZN => n5);
   U90 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U91 : AOI22_X1 port map( A1 => A(5), A2 => n261, B1 => B(5), B2 => n258, ZN 
                           => n17);
   U92 : AOI222_X1 port map( A1 => D(5), A2 => n270, B1 => E(5), B2 => n267, C1
                           => C(5), C2 => n264, ZN => n18);
   U93 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U94 : AOI22_X1 port map( A1 => A(31), A2 => n261, B1 => B(31), B2 => n258, 
                           ZN => n23);
   U95 : AOI222_X1 port map( A1 => D(31), A2 => n270, B1 => E(31), B2 => n267, 
                           C1 => C(31), C2 => n264, ZN => n24);
   U96 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U97 : AOI22_X1 port map( A1 => A(2), A2 => n260, B1 => B(2), B2 => n257, ZN 
                           => n27);
   U98 : AOI222_X1 port map( A1 => D(2), A2 => n269, B1 => E(2), B2 => n266, C1
                           => C(2), C2 => n263, ZN => n28);
   U99 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U100 : AOI22_X1 port map( A1 => A(10), A2 => n259, B1 => B(10), B2 => n256, 
                           ZN => n69);
   U101 : AOI222_X1 port map( A1 => D(10), A2 => n268, B1 => E(10), B2 => n265,
                           C1 => C(10), C2 => n262, ZN => n70);
   U102 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U103 : AOI22_X1 port map( A1 => A(11), A2 => n259, B1 => B(11), B2 => n256, 
                           ZN => n67);
   U104 : AOI222_X1 port map( A1 => D(11), A2 => n268, B1 => E(11), B2 => n265,
                           C1 => C(11), C2 => n262, ZN => n68);
   U105 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U106 : AOI22_X1 port map( A1 => A(0), A2 => n259, B1 => B(0), B2 => n256, ZN
                           => n71);
   U107 : AOI222_X1 port map( A1 => D(0), A2 => n268, B1 => E(0), B2 => n265, 
                           C1 => C(0), C2 => n262, ZN => n72);
   U108 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U109 : AOI22_X1 port map( A1 => A(12), A2 => n259, B1 => B(12), B2 => n256, 
                           ZN => n65);
   U110 : AOI222_X1 port map( A1 => D(12), A2 => n268, B1 => E(12), B2 => n265,
                           C1 => C(12), C2 => n262, ZN => n66);
   U111 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U112 : AOI22_X1 port map( A1 => A(13), A2 => n259, B1 => B(13), B2 => n256, 
                           ZN => n63);
   U113 : AOI222_X1 port map( A1 => D(13), A2 => n268, B1 => E(13), B2 => n265,
                           C1 => C(13), C2 => n262, ZN => n64);
   U114 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U115 : AOI22_X1 port map( A1 => A(1), A2 => n259, B1 => B(1), B2 => n256, ZN
                           => n49);
   U116 : AOI222_X1 port map( A1 => D(1), A2 => n268, B1 => E(1), B2 => n265, 
                           C1 => C(1), C2 => n262, ZN => n50);
   U117 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U118 : AOI22_X1 port map( A1 => A(30), A2 => n260, B1 => B(30), B2 => n257, 
                           ZN => n25);
   U119 : AOI222_X1 port map( A1 => D(30), A2 => n269, B1 => E(30), B2 => n266,
                           C1 => C(30), C2 => n263, ZN => n26);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_2 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_2;

architecture SYN_behav of mux_N32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n269);
   U2 : BUF_X1 port map( A => n10, Z => n268);
   U3 : BUF_X1 port map( A => n10, Z => n270);
   U4 : BUF_X1 port map( A => n6, Z => n281);
   U5 : BUF_X1 port map( A => n6, Z => n280);
   U6 : BUF_X1 port map( A => n9, Z => n272);
   U7 : BUF_X1 port map( A => n9, Z => n271);
   U8 : BUF_X1 port map( A => n7, Z => n278);
   U9 : BUF_X1 port map( A => n7, Z => n277);
   U10 : BUF_X1 port map( A => n8, Z => n275);
   U11 : BUF_X1 port map( A => n8, Z => n274);
   U12 : BUF_X1 port map( A => n9, Z => n273);
   U13 : BUF_X1 port map( A => n7, Z => n279);
   U14 : BUF_X1 port map( A => n8, Z => n276);
   U15 : BUF_X1 port map( A => n6, Z => n282);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U24 : AOI22_X1 port map( A1 => A(26), A2 => n272, B1 => B(26), B2 => n269, 
                           ZN => n35);
   U25 : AOI222_X1 port map( A1 => D(26), A2 => n281, B1 => E(26), B2 => n278, 
                           C1 => C(26), C2 => n275, ZN => n36);
   U26 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U27 : AOI22_X1 port map( A1 => A(22), A2 => n272, B1 => B(22), B2 => n269, 
                           ZN => n43);
   U28 : AOI222_X1 port map( A1 => D(22), A2 => n281, B1 => E(22), B2 => n278, 
                           C1 => C(22), C2 => n275, ZN => n44);
   U29 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U30 : AOI22_X1 port map( A1 => A(28), A2 => n272, B1 => B(28), B2 => n269, 
                           ZN => n31);
   U31 : AOI222_X1 port map( A1 => D(28), A2 => n281, B1 => E(28), B2 => n278, 
                           C1 => C(28), C2 => n275, ZN => n32);
   U32 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U33 : AOI22_X1 port map( A1 => A(29), A2 => n272, B1 => B(29), B2 => n269, 
                           ZN => n29);
   U34 : AOI222_X1 port map( A1 => D(29), A2 => n281, B1 => E(29), B2 => n278, 
                           C1 => C(29), C2 => n275, ZN => n30);
   U35 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U36 : AOI22_X1 port map( A1 => A(30), A2 => n272, B1 => B(30), B2 => n269, 
                           ZN => n25);
   U37 : AOI222_X1 port map( A1 => D(30), A2 => n281, B1 => E(30), B2 => n278, 
                           C1 => C(30), C2 => n275, ZN => n26);
   U38 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U39 : AOI22_X1 port map( A1 => A(31), A2 => n273, B1 => B(31), B2 => n270, 
                           ZN => n23);
   U40 : AOI222_X1 port map( A1 => D(31), A2 => n282, B1 => E(31), B2 => n279, 
                           C1 => C(31), C2 => n276, ZN => n24);
   U41 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U42 : AOI22_X1 port map( A1 => A(16), A2 => n271, B1 => B(16), B2 => n268, 
                           ZN => n57);
   U43 : AOI222_X1 port map( A1 => D(16), A2 => n280, B1 => E(16), B2 => n277, 
                           C1 => C(16), C2 => n274, ZN => n58);
   U44 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n272, B1 => B(20), B2 => n269, 
                           ZN => n47);
   U46 : AOI222_X1 port map( A1 => D(20), A2 => n281, B1 => E(20), B2 => n278, 
                           C1 => C(20), C2 => n275, ZN => n48);
   U47 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U48 : AOI22_X1 port map( A1 => A(14), A2 => n271, B1 => B(14), B2 => n268, 
                           ZN => n61);
   U49 : AOI222_X1 port map( A1 => D(14), A2 => n280, B1 => E(14), B2 => n277, 
                           C1 => C(14), C2 => n274, ZN => n62);
   U50 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U51 : AOI22_X1 port map( A1 => A(18), A2 => n271, B1 => B(18), B2 => n268, 
                           ZN => n53);
   U52 : AOI222_X1 port map( A1 => D(18), A2 => n280, B1 => E(18), B2 => n277, 
                           C1 => C(18), C2 => n274, ZN => n54);
   U53 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n272, B1 => B(25), B2 => n269, 
                           ZN => n37);
   U55 : AOI222_X1 port map( A1 => D(25), A2 => n281, B1 => E(25), B2 => n278, 
                           C1 => C(25), C2 => n275, ZN => n38);
   U56 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U57 : AOI22_X1 port map( A1 => A(21), A2 => n272, B1 => B(21), B2 => n269, 
                           ZN => n45);
   U58 : AOI222_X1 port map( A1 => D(21), A2 => n281, B1 => E(21), B2 => n278, 
                           C1 => C(21), C2 => n275, ZN => n46);
   U59 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U60 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U61 : AOI22_X1 port map( A1 => A(15), A2 => n271, B1 => B(15), B2 => n268, 
                           ZN => n59);
   U62 : AOI222_X1 port map( A1 => D(15), A2 => n280, B1 => E(15), B2 => n277, 
                           C1 => C(15), C2 => n274, ZN => n60);
   U63 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U64 : AOI22_X1 port map( A1 => A(19), A2 => n271, B1 => B(19), B2 => n268, 
                           ZN => n51);
   U65 : AOI222_X1 port map( A1 => D(19), A2 => n280, B1 => E(19), B2 => n277, 
                           C1 => C(19), C2 => n274, ZN => n52);
   U66 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U67 : AOI22_X1 port map( A1 => A(17), A2 => n271, B1 => B(17), B2 => n268, 
                           ZN => n55);
   U68 : AOI222_X1 port map( A1 => D(17), A2 => n280, B1 => E(17), B2 => n277, 
                           C1 => C(17), C2 => n274, ZN => n56);
   U69 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U70 : AOI22_X1 port map( A1 => A(12), A2 => n271, B1 => B(12), B2 => n268, 
                           ZN => n65);
   U71 : AOI222_X1 port map( A1 => D(12), A2 => n280, B1 => E(12), B2 => n277, 
                           C1 => C(12), C2 => n274, ZN => n66);
   U72 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U73 : AOI22_X1 port map( A1 => A(13), A2 => n271, B1 => B(13), B2 => n268, 
                           ZN => n63);
   U74 : AOI222_X1 port map( A1 => D(13), A2 => n280, B1 => E(13), B2 => n277, 
                           C1 => C(13), C2 => n274, ZN => n64);
   U75 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U76 : AOI22_X1 port map( A1 => A(23), A2 => n272, B1 => B(23), B2 => n269, 
                           ZN => n41);
   U77 : AOI222_X1 port map( A1 => D(23), A2 => n281, B1 => E(23), B2 => n278, 
                           C1 => C(23), C2 => n275, ZN => n42);
   U78 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U79 : AOI22_X1 port map( A1 => A(27), A2 => n272, B1 => B(27), B2 => n269, 
                           ZN => n33);
   U80 : AOI222_X1 port map( A1 => D(27), A2 => n281, B1 => E(27), B2 => n278, 
                           C1 => C(27), C2 => n275, ZN => n34);
   U81 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U82 : AOI22_X1 port map( A1 => A(24), A2 => n272, B1 => B(24), B2 => n269, 
                           ZN => n39);
   U83 : AOI222_X1 port map( A1 => D(24), A2 => n281, B1 => E(24), B2 => n278, 
                           C1 => C(24), C2 => n275, ZN => n40);
   U84 : INV_X1 port map( A => Sel(1), ZN => n75);
   U85 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U86 : AOI22_X1 port map( A1 => A(6), A2 => n273, B1 => B(6), B2 => n270, ZN 
                           => n15);
   U87 : AOI222_X1 port map( A1 => D(6), A2 => n282, B1 => E(6), B2 => n279, C1
                           => C(6), C2 => n276, ZN => n16);
   U88 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U89 : AOI22_X1 port map( A1 => A(3), A2 => n273, B1 => B(3), B2 => n270, ZN 
                           => n21);
   U90 : AOI222_X1 port map( A1 => D(3), A2 => n282, B1 => E(3), B2 => n279, C1
                           => C(3), C2 => n276, ZN => n22);
   U91 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U92 : AOI22_X1 port map( A1 => A(7), A2 => n273, B1 => B(7), B2 => n270, ZN 
                           => n13);
   U93 : AOI222_X1 port map( A1 => D(7), A2 => n282, B1 => E(7), B2 => n279, C1
                           => C(7), C2 => n276, ZN => n14);
   U94 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U95 : AOI22_X1 port map( A1 => A(4), A2 => n273, B1 => B(4), B2 => n270, ZN 
                           => n19);
   U96 : AOI222_X1 port map( A1 => D(4), A2 => n282, B1 => E(4), B2 => n279, C1
                           => C(4), C2 => n276, ZN => n20);
   U97 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U98 : AOI22_X1 port map( A1 => A(8), A2 => n273, B1 => B(8), B2 => n270, ZN 
                           => n11);
   U99 : AOI222_X1 port map( A1 => D(8), A2 => n282, B1 => E(8), B2 => n279, C1
                           => C(8), C2 => n276, ZN => n12);
   U100 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U101 : AOI22_X1 port map( A1 => A(9), A2 => n273, B1 => B(9), B2 => n270, ZN
                           => n4);
   U102 : AOI222_X1 port map( A1 => D(9), A2 => n282, B1 => E(9), B2 => n279, 
                           C1 => C(9), C2 => n276, ZN => n5);
   U103 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U104 : AOI22_X1 port map( A1 => A(5), A2 => n273, B1 => B(5), B2 => n270, ZN
                           => n17);
   U105 : AOI222_X1 port map( A1 => D(5), A2 => n282, B1 => E(5), B2 => n279, 
                           C1 => C(5), C2 => n276, ZN => n18);
   U106 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U107 : AOI22_X1 port map( A1 => A(2), A2 => n272, B1 => B(2), B2 => n269, ZN
                           => n27);
   U108 : AOI222_X1 port map( A1 => D(2), A2 => n281, B1 => E(2), B2 => n278, 
                           C1 => C(2), C2 => n275, ZN => n28);
   U109 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U110 : AOI22_X1 port map( A1 => A(10), A2 => n271, B1 => B(10), B2 => n268, 
                           ZN => n69);
   U111 : AOI222_X1 port map( A1 => D(10), A2 => n280, B1 => E(10), B2 => n277,
                           C1 => C(10), C2 => n274, ZN => n70);
   U112 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U113 : AOI22_X1 port map( A1 => A(11), A2 => n271, B1 => B(11), B2 => n268, 
                           ZN => n67);
   U114 : AOI222_X1 port map( A1 => D(11), A2 => n280, B1 => E(11), B2 => n277,
                           C1 => C(11), C2 => n274, ZN => n68);
   U115 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U116 : AOI22_X1 port map( A1 => A(0), A2 => n271, B1 => B(0), B2 => n268, ZN
                           => n71);
   U117 : AOI222_X1 port map( A1 => D(0), A2 => n280, B1 => E(0), B2 => n277, 
                           C1 => C(0), C2 => n274, ZN => n72);
   U118 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U119 : AOI22_X1 port map( A1 => A(1), A2 => n271, B1 => B(1), B2 => n268, ZN
                           => n49);
   U120 : AOI222_X1 port map( A1 => D(1), A2 => n280, B1 => E(1), B2 => n277, 
                           C1 => C(1), C2 => n274, ZN => n50);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_3 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_3;

architecture SYN_behav of mux_N32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n265);
   U2 : BUF_X1 port map( A => n10, Z => n266);
   U3 : BUF_X1 port map( A => n10, Z => n267);
   U4 : BUF_X1 port map( A => n6, Z => n277);
   U5 : BUF_X1 port map( A => n6, Z => n278);
   U6 : BUF_X1 port map( A => n9, Z => n268);
   U7 : BUF_X1 port map( A => n9, Z => n269);
   U8 : BUF_X1 port map( A => n7, Z => n274);
   U9 : BUF_X1 port map( A => n7, Z => n275);
   U10 : BUF_X1 port map( A => n8, Z => n271);
   U11 : BUF_X1 port map( A => n8, Z => n272);
   U12 : BUF_X1 port map( A => n9, Z => n270);
   U13 : BUF_X1 port map( A => n7, Z => n276);
   U14 : BUF_X1 port map( A => n8, Z => n273);
   U15 : BUF_X1 port map( A => n6, Z => n279);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U24 : AOI22_X1 port map( A1 => A(24), A2 => n269, B1 => B(24), B2 => n266, 
                           ZN => n39);
   U25 : AOI222_X1 port map( A1 => D(24), A2 => n278, B1 => E(24), B2 => n275, 
                           C1 => C(24), C2 => n272, ZN => n40);
   U26 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U27 : AOI22_X1 port map( A1 => A(20), A2 => n269, B1 => B(20), B2 => n266, 
                           ZN => n47);
   U28 : AOI222_X1 port map( A1 => D(20), A2 => n278, B1 => E(20), B2 => n275, 
                           C1 => C(20), C2 => n272, ZN => n48);
   U29 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U30 : AOI22_X1 port map( A1 => A(14), A2 => n268, B1 => B(14), B2 => n265, 
                           ZN => n61);
   U31 : AOI222_X1 port map( A1 => D(14), A2 => n277, B1 => E(14), B2 => n274, 
                           C1 => C(14), C2 => n271, ZN => n62);
   U32 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U33 : AOI22_X1 port map( A1 => A(18), A2 => n268, B1 => B(18), B2 => n265, 
                           ZN => n53);
   U34 : AOI222_X1 port map( A1 => D(18), A2 => n277, B1 => E(18), B2 => n274, 
                           C1 => C(18), C2 => n271, ZN => n54);
   U35 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U36 : AOI22_X1 port map( A1 => A(12), A2 => n268, B1 => B(12), B2 => n265, 
                           ZN => n65);
   U37 : AOI222_X1 port map( A1 => D(12), A2 => n277, B1 => E(12), B2 => n274, 
                           C1 => C(12), C2 => n271, ZN => n66);
   U38 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U39 : AOI22_X1 port map( A1 => A(16), A2 => n268, B1 => B(16), B2 => n265, 
                           ZN => n57);
   U40 : AOI222_X1 port map( A1 => D(16), A2 => n277, B1 => E(16), B2 => n274, 
                           C1 => C(16), C2 => n271, ZN => n58);
   U41 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U42 : AOI22_X1 port map( A1 => A(23), A2 => n269, B1 => B(23), B2 => n266, 
                           ZN => n41);
   U43 : AOI222_X1 port map( A1 => D(23), A2 => n278, B1 => E(23), B2 => n275, 
                           C1 => C(23), C2 => n272, ZN => n42);
   U44 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U45 : AOI22_X1 port map( A1 => A(19), A2 => n268, B1 => B(19), B2 => n265, 
                           ZN => n51);
   U46 : AOI222_X1 port map( A1 => D(19), A2 => n277, B1 => E(19), B2 => n274, 
                           C1 => C(19), C2 => n271, ZN => n52);
   U47 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U48 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U49 : AOI22_X1 port map( A1 => A(13), A2 => n268, B1 => B(13), B2 => n265, 
                           ZN => n63);
   U50 : AOI222_X1 port map( A1 => D(13), A2 => n277, B1 => E(13), B2 => n274, 
                           C1 => C(13), C2 => n271, ZN => n64);
   U51 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U52 : AOI22_X1 port map( A1 => A(17), A2 => n268, B1 => B(17), B2 => n265, 
                           ZN => n55);
   U53 : AOI222_X1 port map( A1 => D(17), A2 => n277, B1 => E(17), B2 => n274, 
                           C1 => C(17), C2 => n271, ZN => n56);
   U54 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U55 : AOI22_X1 port map( A1 => A(15), A2 => n268, B1 => B(15), B2 => n265, 
                           ZN => n59);
   U56 : AOI222_X1 port map( A1 => D(15), A2 => n277, B1 => E(15), B2 => n274, 
                           C1 => C(15), C2 => n271, ZN => n60);
   U57 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U58 : AOI22_X1 port map( A1 => A(10), A2 => n268, B1 => B(10), B2 => n265, 
                           ZN => n69);
   U59 : AOI222_X1 port map( A1 => D(10), A2 => n277, B1 => E(10), B2 => n274, 
                           C1 => C(10), C2 => n271, ZN => n70);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U61 : AOI22_X1 port map( A1 => A(11), A2 => n268, B1 => B(11), B2 => n265, 
                           ZN => n67);
   U62 : AOI222_X1 port map( A1 => D(11), A2 => n277, B1 => E(11), B2 => n274, 
                           C1 => C(11), C2 => n271, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U64 : AOI22_X1 port map( A1 => A(21), A2 => n269, B1 => B(21), B2 => n266, 
                           ZN => n45);
   U65 : AOI222_X1 port map( A1 => D(21), A2 => n278, B1 => E(21), B2 => n275, 
                           C1 => C(21), C2 => n272, ZN => n46);
   U66 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U67 : AOI22_X1 port map( A1 => A(25), A2 => n269, B1 => B(25), B2 => n266, 
                           ZN => n37);
   U68 : AOI222_X1 port map( A1 => D(25), A2 => n278, B1 => E(25), B2 => n275, 
                           C1 => C(25), C2 => n272, ZN => n38);
   U69 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U70 : AOI22_X1 port map( A1 => A(26), A2 => n269, B1 => B(26), B2 => n266, 
                           ZN => n35);
   U71 : AOI222_X1 port map( A1 => D(26), A2 => n278, B1 => E(26), B2 => n275, 
                           C1 => C(26), C2 => n272, ZN => n36);
   U72 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U73 : AOI22_X1 port map( A1 => A(27), A2 => n269, B1 => B(27), B2 => n266, 
                           ZN => n33);
   U74 : AOI222_X1 port map( A1 => D(27), A2 => n278, B1 => E(27), B2 => n275, 
                           C1 => C(27), C2 => n272, ZN => n34);
   U75 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U76 : AOI22_X1 port map( A1 => A(28), A2 => n269, B1 => B(28), B2 => n266, 
                           ZN => n31);
   U77 : AOI222_X1 port map( A1 => D(28), A2 => n278, B1 => E(28), B2 => n275, 
                           C1 => C(28), C2 => n272, ZN => n32);
   U78 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U79 : AOI22_X1 port map( A1 => A(29), A2 => n269, B1 => B(29), B2 => n266, 
                           ZN => n29);
   U80 : AOI222_X1 port map( A1 => D(29), A2 => n278, B1 => E(29), B2 => n275, 
                           C1 => C(29), C2 => n272, ZN => n30);
   U81 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U82 : AOI22_X1 port map( A1 => A(30), A2 => n269, B1 => B(30), B2 => n266, 
                           ZN => n25);
   U83 : AOI222_X1 port map( A1 => D(30), A2 => n278, B1 => E(30), B2 => n275, 
                           C1 => C(30), C2 => n272, ZN => n26);
   U84 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U85 : AOI22_X1 port map( A1 => A(31), A2 => n270, B1 => B(31), B2 => n267, 
                           ZN => n23);
   U86 : AOI222_X1 port map( A1 => D(31), A2 => n279, B1 => E(31), B2 => n276, 
                           C1 => C(31), C2 => n273, ZN => n24);
   U87 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U88 : AOI22_X1 port map( A1 => A(22), A2 => n269, B1 => B(22), B2 => n266, 
                           ZN => n43);
   U89 : AOI222_X1 port map( A1 => D(22), A2 => n278, B1 => E(22), B2 => n275, 
                           C1 => C(22), C2 => n272, ZN => n44);
   U90 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U91 : AOI22_X1 port map( A1 => A(9), A2 => n270, B1 => B(9), B2 => n267, ZN 
                           => n4);
   U92 : AOI222_X1 port map( A1 => D(9), A2 => n279, B1 => E(9), B2 => n276, C1
                           => C(9), C2 => n273, ZN => n5);
   U93 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U94 : AOI22_X1 port map( A1 => A(5), A2 => n270, B1 => B(5), B2 => n267, ZN 
                           => n17);
   U95 : AOI222_X1 port map( A1 => D(5), A2 => n279, B1 => E(5), B2 => n276, C1
                           => C(5), C2 => n273, ZN => n18);
   U96 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U97 : AOI22_X1 port map( A1 => A(6), A2 => n270, B1 => B(6), B2 => n267, ZN 
                           => n15);
   U98 : AOI222_X1 port map( A1 => D(6), A2 => n279, B1 => E(6), B2 => n276, C1
                           => C(6), C2 => n273, ZN => n16);
   U99 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U100 : AOI22_X1 port map( A1 => A(3), A2 => n270, B1 => B(3), B2 => n267, ZN
                           => n21);
   U101 : AOI222_X1 port map( A1 => D(3), A2 => n279, B1 => E(3), B2 => n276, 
                           C1 => C(3), C2 => n273, ZN => n22);
   U102 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U103 : AOI22_X1 port map( A1 => A(7), A2 => n270, B1 => B(7), B2 => n267, ZN
                           => n13);
   U104 : AOI222_X1 port map( A1 => D(7), A2 => n279, B1 => E(7), B2 => n276, 
                           C1 => C(7), C2 => n273, ZN => n14);
   U105 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U106 : AOI22_X1 port map( A1 => A(4), A2 => n270, B1 => B(4), B2 => n267, ZN
                           => n19);
   U107 : AOI222_X1 port map( A1 => D(4), A2 => n279, B1 => E(4), B2 => n276, 
                           C1 => C(4), C2 => n273, ZN => n20);
   U108 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U109 : AOI22_X1 port map( A1 => A(8), A2 => n270, B1 => B(8), B2 => n267, ZN
                           => n11);
   U110 : AOI222_X1 port map( A1 => D(8), A2 => n279, B1 => E(8), B2 => n276, 
                           C1 => C(8), C2 => n273, ZN => n12);
   U111 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U112 : AOI22_X1 port map( A1 => A(1), A2 => n268, B1 => B(1), B2 => n265, ZN
                           => n49);
   U113 : AOI222_X1 port map( A1 => D(1), A2 => n277, B1 => E(1), B2 => n274, 
                           C1 => C(1), C2 => n271, ZN => n50);
   U114 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U115 : AOI22_X1 port map( A1 => A(2), A2 => n269, B1 => B(2), B2 => n266, ZN
                           => n27);
   U116 : AOI222_X1 port map( A1 => D(2), A2 => n278, B1 => E(2), B2 => n275, 
                           C1 => C(2), C2 => n272, ZN => n28);
   U117 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U118 : AOI22_X1 port map( A1 => A(0), A2 => n268, B1 => B(0), B2 => n265, ZN
                           => n71);
   U119 : AOI222_X1 port map( A1 => D(0), A2 => n277, B1 => E(0), B2 => n274, 
                           C1 => C(0), C2 => n271, ZN => n72);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_4 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_4;

architecture SYN_behav of mux_N32_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n280);
   U2 : BUF_X1 port map( A => n10, Z => n281);
   U3 : BUF_X1 port map( A => n10, Z => n282);
   U4 : BUF_X1 port map( A => n6, Z => n292);
   U5 : BUF_X1 port map( A => n6, Z => n293);
   U6 : BUF_X1 port map( A => n9, Z => n283);
   U7 : BUF_X1 port map( A => n9, Z => n284);
   U8 : BUF_X1 port map( A => n7, Z => n289);
   U9 : BUF_X1 port map( A => n7, Z => n290);
   U10 : BUF_X1 port map( A => n8, Z => n286);
   U11 : BUF_X1 port map( A => n8, Z => n287);
   U12 : BUF_X1 port map( A => n9, Z => n285);
   U13 : BUF_X1 port map( A => n7, Z => n291);
   U14 : BUF_X1 port map( A => n8, Z => n288);
   U15 : BUF_X1 port map( A => n6, Z => n294);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U24 : AOI22_X1 port map( A1 => A(22), A2 => n284, B1 => B(22), B2 => n281, 
                           ZN => n43);
   U25 : AOI222_X1 port map( A1 => D(22), A2 => n293, B1 => E(22), B2 => n290, 
                           C1 => C(22), C2 => n287, ZN => n44);
   U26 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U27 : AOI22_X1 port map( A1 => A(8), A2 => n285, B1 => B(8), B2 => n282, ZN 
                           => n11);
   U28 : AOI222_X1 port map( A1 => D(8), A2 => n294, B1 => E(8), B2 => n291, C1
                           => C(8), C2 => n288, ZN => n12);
   U29 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U30 : AOI22_X1 port map( A1 => A(18), A2 => n283, B1 => B(18), B2 => n280, 
                           ZN => n53);
   U31 : AOI222_X1 port map( A1 => D(18), A2 => n292, B1 => E(18), B2 => n289, 
                           C1 => C(18), C2 => n286, ZN => n54);
   U32 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U33 : AOI22_X1 port map( A1 => A(25), A2 => n284, B1 => B(25), B2 => n281, 
                           ZN => n37);
   U34 : AOI222_X1 port map( A1 => D(25), A2 => n293, B1 => E(25), B2 => n290, 
                           C1 => C(25), C2 => n287, ZN => n38);
   U35 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U36 : AOI22_X1 port map( A1 => A(26), A2 => n284, B1 => B(26), B2 => n281, 
                           ZN => n35);
   U37 : AOI222_X1 port map( A1 => D(26), A2 => n293, B1 => E(26), B2 => n290, 
                           C1 => C(26), C2 => n287, ZN => n36);
   U38 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U39 : AOI22_X1 port map( A1 => A(27), A2 => n284, B1 => B(27), B2 => n281, 
                           ZN => n33);
   U40 : AOI222_X1 port map( A1 => D(27), A2 => n293, B1 => E(27), B2 => n290, 
                           C1 => C(27), C2 => n287, ZN => n34);
   U41 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U42 : AOI22_X1 port map( A1 => A(28), A2 => n284, B1 => B(28), B2 => n281, 
                           ZN => n31);
   U43 : AOI222_X1 port map( A1 => D(28), A2 => n293, B1 => E(28), B2 => n290, 
                           C1 => C(28), C2 => n287, ZN => n32);
   U44 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U45 : AOI22_X1 port map( A1 => A(24), A2 => n284, B1 => B(24), B2 => n281, 
                           ZN => n39);
   U46 : AOI222_X1 port map( A1 => D(24), A2 => n293, B1 => E(24), B2 => n290, 
                           C1 => C(24), C2 => n287, ZN => n40);
   U47 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U48 : AOI22_X1 port map( A1 => A(29), A2 => n284, B1 => B(29), B2 => n281, 
                           ZN => n29);
   U49 : AOI222_X1 port map( A1 => D(29), A2 => n293, B1 => E(29), B2 => n290, 
                           C1 => C(29), C2 => n287, ZN => n30);
   U50 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U51 : AOI22_X1 port map( A1 => A(30), A2 => n284, B1 => B(30), B2 => n281, 
                           ZN => n25);
   U52 : AOI222_X1 port map( A1 => D(30), A2 => n293, B1 => E(30), B2 => n290, 
                           C1 => C(30), C2 => n287, ZN => n26);
   U53 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U54 : AOI22_X1 port map( A1 => A(31), A2 => n285, B1 => B(31), B2 => n282, 
                           ZN => n23);
   U55 : AOI222_X1 port map( A1 => D(31), A2 => n294, B1 => E(31), B2 => n291, 
                           C1 => C(31), C2 => n288, ZN => n24);
   U56 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U57 : AOI22_X1 port map( A1 => A(12), A2 => n283, B1 => B(12), B2 => n280, 
                           ZN => n65);
   U58 : AOI222_X1 port map( A1 => D(12), A2 => n292, B1 => E(12), B2 => n289, 
                           C1 => C(12), C2 => n286, ZN => n66);
   U59 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U60 : AOI22_X1 port map( A1 => A(9), A2 => n285, B1 => B(9), B2 => n282, ZN 
                           => n4);
   U61 : AOI222_X1 port map( A1 => D(9), A2 => n294, B1 => E(9), B2 => n291, C1
                           => C(9), C2 => n288, ZN => n5);
   U62 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U63 : AOI22_X1 port map( A1 => A(16), A2 => n283, B1 => B(16), B2 => n280, 
                           ZN => n57);
   U64 : AOI222_X1 port map( A1 => D(16), A2 => n292, B1 => E(16), B2 => n289, 
                           C1 => C(16), C2 => n286, ZN => n58);
   U65 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U66 : AOI22_X1 port map( A1 => A(10), A2 => n283, B1 => B(10), B2 => n280, 
                           ZN => n69);
   U67 : AOI222_X1 port map( A1 => D(10), A2 => n292, B1 => E(10), B2 => n289, 
                           C1 => C(10), C2 => n286, ZN => n70);
   U68 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U69 : AOI22_X1 port map( A1 => A(14), A2 => n283, B1 => B(14), B2 => n280, 
                           ZN => n61);
   U70 : AOI222_X1 port map( A1 => D(14), A2 => n292, B1 => E(14), B2 => n289, 
                           C1 => C(14), C2 => n286, ZN => n62);
   U71 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U72 : AOI22_X1 port map( A1 => A(21), A2 => n284, B1 => B(21), B2 => n281, 
                           ZN => n45);
   U73 : AOI222_X1 port map( A1 => D(21), A2 => n293, B1 => E(21), B2 => n290, 
                           C1 => C(21), C2 => n287, ZN => n46);
   U74 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U75 : AOI22_X1 port map( A1 => A(17), A2 => n283, B1 => B(17), B2 => n280, 
                           ZN => n55);
   U76 : AOI222_X1 port map( A1 => D(17), A2 => n292, B1 => E(17), B2 => n289, 
                           C1 => C(17), C2 => n286, ZN => n56);
   U77 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U78 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U79 : AOI22_X1 port map( A1 => A(11), A2 => n283, B1 => B(11), B2 => n280, 
                           ZN => n67);
   U80 : AOI222_X1 port map( A1 => D(11), A2 => n292, B1 => E(11), B2 => n289, 
                           C1 => C(11), C2 => n286, ZN => n68);
   U81 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U82 : AOI22_X1 port map( A1 => A(15), A2 => n283, B1 => B(15), B2 => n280, 
                           ZN => n59);
   U83 : AOI222_X1 port map( A1 => D(15), A2 => n292, B1 => E(15), B2 => n289, 
                           C1 => C(15), C2 => n286, ZN => n60);
   U84 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U85 : AOI22_X1 port map( A1 => A(13), A2 => n283, B1 => B(13), B2 => n280, 
                           ZN => n63);
   U86 : AOI222_X1 port map( A1 => D(13), A2 => n292, B1 => E(13), B2 => n289, 
                           C1 => C(13), C2 => n286, ZN => n64);
   U87 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U88 : AOI22_X1 port map( A1 => A(20), A2 => n284, B1 => B(20), B2 => n281, 
                           ZN => n47);
   U89 : AOI222_X1 port map( A1 => D(20), A2 => n293, B1 => E(20), B2 => n290, 
                           C1 => C(20), C2 => n287, ZN => n48);
   U90 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U91 : AOI22_X1 port map( A1 => A(19), A2 => n283, B1 => B(19), B2 => n280, 
                           ZN => n51);
   U92 : AOI222_X1 port map( A1 => D(19), A2 => n292, B1 => E(19), B2 => n289, 
                           C1 => C(19), C2 => n286, ZN => n52);
   U93 : INV_X1 port map( A => Sel(1), ZN => n75);
   U94 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U95 : AOI22_X1 port map( A1 => A(5), A2 => n285, B1 => B(5), B2 => n282, ZN 
                           => n17);
   U96 : AOI222_X1 port map( A1 => D(5), A2 => n294, B1 => E(5), B2 => n291, C1
                           => C(5), C2 => n288, ZN => n18);
   U97 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U98 : AOI22_X1 port map( A1 => A(6), A2 => n285, B1 => B(6), B2 => n282, ZN 
                           => n15);
   U99 : AOI222_X1 port map( A1 => D(6), A2 => n294, B1 => E(6), B2 => n291, C1
                           => C(6), C2 => n288, ZN => n16);
   U100 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U101 : AOI22_X1 port map( A1 => A(3), A2 => n285, B1 => B(3), B2 => n282, ZN
                           => n21);
   U102 : AOI222_X1 port map( A1 => D(3), A2 => n294, B1 => E(3), B2 => n291, 
                           C1 => C(3), C2 => n288, ZN => n22);
   U103 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U104 : AOI22_X1 port map( A1 => A(7), A2 => n285, B1 => B(7), B2 => n282, ZN
                           => n13);
   U105 : AOI222_X1 port map( A1 => D(7), A2 => n294, B1 => E(7), B2 => n291, 
                           C1 => C(7), C2 => n288, ZN => n14);
   U106 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U107 : AOI22_X1 port map( A1 => A(4), A2 => n285, B1 => B(4), B2 => n282, ZN
                           => n19);
   U108 : AOI222_X1 port map( A1 => D(4), A2 => n294, B1 => E(4), B2 => n291, 
                           C1 => C(4), C2 => n288, ZN => n20);
   U109 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U110 : AOI22_X1 port map( A1 => A(1), A2 => n283, B1 => B(1), B2 => n280, ZN
                           => n49);
   U111 : AOI222_X1 port map( A1 => D(1), A2 => n292, B1 => E(1), B2 => n289, 
                           C1 => C(1), C2 => n286, ZN => n50);
   U112 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U113 : AOI22_X1 port map( A1 => A(2), A2 => n284, B1 => B(2), B2 => n281, ZN
                           => n27);
   U114 : AOI222_X1 port map( A1 => D(2), A2 => n293, B1 => E(2), B2 => n290, 
                           C1 => C(2), C2 => n287, ZN => n28);
   U115 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U116 : AOI22_X1 port map( A1 => A(23), A2 => n284, B1 => B(23), B2 => n281, 
                           ZN => n41);
   U117 : AOI222_X1 port map( A1 => D(23), A2 => n293, B1 => E(23), B2 => n290,
                           C1 => C(23), C2 => n287, ZN => n42);
   U118 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U119 : AOI22_X1 port map( A1 => A(0), A2 => n283, B1 => B(0), B2 => n280, ZN
                           => n71);
   U120 : AOI222_X1 port map( A1 => D(0), A2 => n292, B1 => E(0), B2 => n289, 
                           C1 => C(0), C2 => n286, ZN => n72);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_5 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_5;

architecture SYN_behav of mux_N32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n274);
   U2 : BUF_X1 port map( A => n10, Z => n275);
   U3 : BUF_X1 port map( A => n10, Z => n276);
   U4 : BUF_X1 port map( A => n6, Z => n286);
   U5 : BUF_X1 port map( A => n6, Z => n287);
   U6 : BUF_X1 port map( A => n9, Z => n277);
   U7 : BUF_X1 port map( A => n9, Z => n278);
   U8 : BUF_X1 port map( A => n7, Z => n283);
   U9 : BUF_X1 port map( A => n7, Z => n284);
   U10 : BUF_X1 port map( A => n8, Z => n280);
   U11 : BUF_X1 port map( A => n8, Z => n281);
   U12 : BUF_X1 port map( A => n9, Z => n279);
   U13 : BUF_X1 port map( A => n7, Z => n285);
   U14 : BUF_X1 port map( A => n8, Z => n282);
   U15 : BUF_X1 port map( A => n6, Z => n288);
   U16 : AND2_X1 port map( A1 => n74, A2 => n73, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n73, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n73, ZN => n8);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n74);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n73);
   U23 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U24 : AOI22_X1 port map( A1 => A(20), A2 => n278, B1 => B(20), B2 => n275, 
                           ZN => n47);
   U25 : AOI222_X1 port map( A1 => D(20), A2 => n287, B1 => C(20), B2 => n284, 
                           C1 => E(20), C2 => n281, ZN => n48);
   U26 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U27 : AOI22_X1 port map( A1 => A(16), A2 => n277, B1 => B(16), B2 => n274, 
                           ZN => n57);
   U28 : AOI222_X1 port map( A1 => D(16), A2 => n286, B1 => C(16), B2 => n283, 
                           C1 => E(16), C2 => n280, ZN => n58);
   U29 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n277, B1 => B(10), B2 => n274, 
                           ZN => n69);
   U31 : AOI222_X1 port map( A1 => D(10), A2 => n286, B1 => C(10), B2 => n283, 
                           C1 => E(10), C2 => n280, ZN => n70);
   U32 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n277, B1 => B(14), B2 => n274, 
                           ZN => n61);
   U34 : AOI222_X1 port map( A1 => D(14), A2 => n286, B1 => C(14), B2 => n283, 
                           C1 => E(14), C2 => n280, ZN => n62);
   U35 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n279, B1 => B(8), B2 => n276, ZN 
                           => n11);
   U37 : AOI222_X1 port map( A1 => D(8), A2 => n288, B1 => C(8), B2 => n285, C1
                           => E(8), C2 => n282, ZN => n12);
   U38 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U39 : AOI22_X1 port map( A1 => A(12), A2 => n277, B1 => B(12), B2 => n274, 
                           ZN => n65);
   U40 : AOI222_X1 port map( A1 => D(12), A2 => n286, B1 => C(12), B2 => n283, 
                           C1 => E(12), C2 => n280, ZN => n66);
   U41 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U42 : AOI22_X1 port map( A1 => A(19), A2 => n277, B1 => B(19), B2 => n274, 
                           ZN => n51);
   U43 : AOI222_X1 port map( A1 => D(19), A2 => n286, B1 => C(19), B2 => n283, 
                           C1 => E(19), C2 => n280, ZN => n52);
   U44 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U45 : AOI22_X1 port map( A1 => A(15), A2 => n277, B1 => B(15), B2 => n274, 
                           ZN => n59);
   U46 : AOI222_X1 port map( A1 => D(15), A2 => n286, B1 => C(15), B2 => n283, 
                           C1 => E(15), C2 => n280, ZN => n60);
   U47 : AND2_X1 port map( A1 => Sel(2), A2 => n74, ZN => n7);
   U48 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U49 : AOI22_X1 port map( A1 => A(9), A2 => n279, B1 => B(9), B2 => n276, ZN 
                           => n4);
   U50 : AOI222_X1 port map( A1 => D(9), A2 => n288, B1 => C(9), B2 => n285, C1
                           => E(9), C2 => n282, ZN => n5);
   U51 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U52 : AOI22_X1 port map( A1 => A(13), A2 => n277, B1 => B(13), B2 => n274, 
                           ZN => n63);
   U53 : AOI222_X1 port map( A1 => D(13), A2 => n286, B1 => C(13), B2 => n283, 
                           C1 => E(13), C2 => n280, ZN => n64);
   U54 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U55 : AOI22_X1 port map( A1 => A(7), A2 => n279, B1 => B(7), B2 => n276, ZN 
                           => n13);
   U56 : AOI222_X1 port map( A1 => D(7), A2 => n288, B1 => C(7), B2 => n285, C1
                           => E(7), C2 => n282, ZN => n14);
   U57 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U58 : AOI22_X1 port map( A1 => A(17), A2 => n277, B1 => B(17), B2 => n274, 
                           ZN => n55);
   U59 : AOI222_X1 port map( A1 => D(17), A2 => n286, B1 => C(17), B2 => n283, 
                           C1 => E(17), C2 => n280, ZN => n56);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U61 : AOI22_X1 port map( A1 => A(11), A2 => n277, B1 => B(11), B2 => n274, 
                           ZN => n67);
   U62 : AOI222_X1 port map( A1 => D(11), A2 => n286, B1 => C(11), B2 => n283, 
                           C1 => E(11), C2 => n280, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U64 : AOI22_X1 port map( A1 => A(6), A2 => n279, B1 => B(6), B2 => n276, ZN 
                           => n15);
   U65 : AOI222_X1 port map( A1 => D(6), A2 => n288, B1 => C(6), B2 => n285, C1
                           => E(6), C2 => n282, ZN => n16);
   U66 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U67 : AOI22_X1 port map( A1 => A(18), A2 => n277, B1 => B(18), B2 => n274, 
                           ZN => n53);
   U68 : AOI222_X1 port map( A1 => D(18), A2 => n286, B1 => C(18), B2 => n283, 
                           C1 => E(18), C2 => n280, ZN => n54);
   U69 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U70 : AOI22_X1 port map( A1 => A(21), A2 => n278, B1 => B(21), B2 => n275, 
                           ZN => n45);
   U71 : AOI222_X1 port map( A1 => D(21), A2 => n287, B1 => C(21), B2 => n284, 
                           C1 => E(21), C2 => n281, ZN => n46);
   U72 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U73 : AOI22_X1 port map( A1 => A(5), A2 => n279, B1 => B(5), B2 => n276, ZN 
                           => n17);
   U74 : AOI222_X1 port map( A1 => D(5), A2 => n288, B1 => C(5), B2 => n285, C1
                           => E(5), C2 => n282, ZN => n18);
   U75 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U76 : AOI22_X1 port map( A1 => A(3), A2 => n279, B1 => B(3), B2 => n276, ZN 
                           => n21);
   U77 : AOI222_X1 port map( A1 => D(3), A2 => n288, B1 => C(3), B2 => n285, C1
                           => E(3), C2 => n282, ZN => n22);
   U78 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U79 : AOI22_X1 port map( A1 => A(4), A2 => n279, B1 => B(4), B2 => n276, ZN 
                           => n19);
   U80 : AOI222_X1 port map( A1 => D(4), A2 => n288, B1 => C(4), B2 => n285, C1
                           => E(4), C2 => n282, ZN => n20);
   U81 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U82 : AOI22_X1 port map( A1 => A(31), A2 => n279, B1 => B(31), B2 => n276, 
                           ZN => n23);
   U83 : AOI222_X1 port map( A1 => D(31), A2 => n288, B1 => C(31), B2 => n285, 
                           C1 => E(31), C2 => n282, ZN => n24);
   U84 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U85 : AOI22_X1 port map( A1 => A(1), A2 => n277, B1 => B(1), B2 => n274, ZN 
                           => n49);
   U86 : AOI222_X1 port map( A1 => D(1), A2 => n286, B1 => C(1), B2 => n283, C1
                           => E(1), C2 => n280, ZN => n50);
   U87 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U88 : AOI22_X1 port map( A1 => A(25), A2 => n278, B1 => B(25), B2 => n275, 
                           ZN => n37);
   U89 : AOI222_X1 port map( A1 => D(25), A2 => n287, B1 => C(25), B2 => n284, 
                           C1 => E(25), C2 => n281, ZN => n38);
   U90 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U91 : AOI22_X1 port map( A1 => A(2), A2 => n278, B1 => B(2), B2 => n275, ZN 
                           => n27);
   U92 : AOI222_X1 port map( A1 => D(2), A2 => n287, B1 => C(2), B2 => n284, C1
                           => E(2), C2 => n281, ZN => n28);
   U93 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U94 : AOI22_X1 port map( A1 => A(26), A2 => n278, B1 => B(26), B2 => n275, 
                           ZN => n35);
   U95 : AOI222_X1 port map( A1 => D(26), A2 => n287, B1 => C(26), B2 => n284, 
                           C1 => E(26), C2 => n281, ZN => n36);
   U96 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U97 : AOI22_X1 port map( A1 => A(22), A2 => n278, B1 => B(22), B2 => n275, 
                           ZN => n43);
   U98 : AOI222_X1 port map( A1 => D(22), A2 => n287, B1 => C(22), B2 => n284, 
                           C1 => E(22), C2 => n281, ZN => n44);
   U99 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U100 : AOI22_X1 port map( A1 => A(27), A2 => n278, B1 => B(27), B2 => n275, 
                           ZN => n33);
   U101 : AOI222_X1 port map( A1 => D(27), A2 => n287, B1 => C(27), B2 => n284,
                           C1 => E(27), C2 => n281, ZN => n34);
   U102 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U103 : AOI22_X1 port map( A1 => A(23), A2 => n278, B1 => B(23), B2 => n275, 
                           ZN => n41);
   U104 : AOI222_X1 port map( A1 => D(23), A2 => n287, B1 => C(23), B2 => n284,
                           C1 => E(23), C2 => n281, ZN => n42);
   U105 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U106 : AOI22_X1 port map( A1 => A(0), A2 => n277, B1 => B(0), B2 => n274, ZN
                           => n71);
   U107 : AOI222_X1 port map( A1 => D(0), A2 => n286, B1 => C(0), B2 => n283, 
                           C1 => E(0), C2 => n280, ZN => n72);
   U108 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U109 : AOI22_X1 port map( A1 => A(28), A2 => n278, B1 => B(28), B2 => n275, 
                           ZN => n31);
   U110 : AOI222_X1 port map( A1 => D(28), A2 => n287, B1 => C(28), B2 => n284,
                           C1 => E(28), C2 => n281, ZN => n32);
   U111 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U112 : AOI22_X1 port map( A1 => A(24), A2 => n278, B1 => B(24), B2 => n275, 
                           ZN => n39);
   U113 : AOI222_X1 port map( A1 => D(24), A2 => n287, B1 => C(24), B2 => n284,
                           C1 => E(24), C2 => n281, ZN => n40);
   U114 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U115 : AOI22_X1 port map( A1 => A(29), A2 => n278, B1 => B(29), B2 => n275, 
                           ZN => n29);
   U116 : AOI222_X1 port map( A1 => D(29), A2 => n287, B1 => C(29), B2 => n284,
                           C1 => E(29), C2 => n281, ZN => n30);
   U117 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U118 : AOI22_X1 port map( A1 => A(30), A2 => n278, B1 => B(30), B2 => n275, 
                           ZN => n25);
   U119 : AOI222_X1 port map( A1 => D(30), A2 => n287, B1 => C(30), B2 => n284,
                           C1 => E(30), C2 => n281, ZN => n26);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_6 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_6;

architecture SYN_behav of mux_N32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n277);
   U2 : BUF_X1 port map( A => n10, Z => n278);
   U3 : BUF_X1 port map( A => n10, Z => n279);
   U4 : BUF_X1 port map( A => n6, Z => n289);
   U5 : BUF_X1 port map( A => n6, Z => n290);
   U6 : BUF_X1 port map( A => n9, Z => n280);
   U7 : BUF_X1 port map( A => n9, Z => n281);
   U8 : BUF_X1 port map( A => n7, Z => n286);
   U9 : BUF_X1 port map( A => n7, Z => n287);
   U10 : BUF_X1 port map( A => n8, Z => n283);
   U11 : BUF_X1 port map( A => n8, Z => n284);
   U12 : BUF_X1 port map( A => n9, Z => n282);
   U13 : BUF_X1 port map( A => n7, Z => n288);
   U14 : BUF_X1 port map( A => n8, Z => n285);
   U15 : BUF_X1 port map( A => n6, Z => n291);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U23 : AOI22_X1 port map( A1 => A(24), A2 => n281, B1 => B(24), B2 => n278, 
                           ZN => n39);
   U24 : AOI222_X1 port map( A1 => D(24), A2 => n290, B1 => E(24), B2 => n287, 
                           C1 => C(24), C2 => n284, ZN => n40);
   U25 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U26 : AOI22_X1 port map( A1 => A(25), A2 => n281, B1 => B(25), B2 => n278, 
                           ZN => n37);
   U27 : AOI222_X1 port map( A1 => D(25), A2 => n290, B1 => E(25), B2 => n287, 
                           C1 => C(25), C2 => n284, ZN => n38);
   U28 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U29 : AOI22_X1 port map( A1 => A(28), A2 => n281, B1 => B(28), B2 => n278, 
                           ZN => n31);
   U30 : AOI222_X1 port map( A1 => D(28), A2 => n290, B1 => E(28), B2 => n287, 
                           C1 => C(28), C2 => n284, ZN => n32);
   U31 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U32 : AOI22_X1 port map( A1 => A(29), A2 => n281, B1 => B(29), B2 => n278, 
                           ZN => n29);
   U33 : AOI222_X1 port map( A1 => D(29), A2 => n290, B1 => E(29), B2 => n287, 
                           C1 => C(29), C2 => n284, ZN => n30);
   U34 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U35 : AOI22_X1 port map( A1 => A(30), A2 => n281, B1 => B(30), B2 => n278, 
                           ZN => n25);
   U36 : AOI222_X1 port map( A1 => D(30), A2 => n290, B1 => E(30), B2 => n287, 
                           C1 => C(30), C2 => n284, ZN => n26);
   U37 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U38 : AOI22_X1 port map( A1 => A(31), A2 => n282, B1 => B(31), B2 => n279, 
                           ZN => n23);
   U39 : AOI222_X1 port map( A1 => D(31), A2 => n291, B1 => E(31), B2 => n288, 
                           C1 => C(31), C2 => n285, ZN => n24);
   U40 : INV_X1 port map( A => Sel(2), ZN => n74);
   U41 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U42 : AOI22_X1 port map( A1 => A(18), A2 => n280, B1 => B(18), B2 => n277, 
                           ZN => n53);
   U43 : AOI222_X1 port map( A1 => D(18), A2 => n289, B1 => E(18), B2 => n286, 
                           C1 => C(18), C2 => n283, ZN => n54);
   U44 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n282, B1 => B(4), B2 => n279, ZN 
                           => n19);
   U46 : AOI222_X1 port map( A1 => D(4), A2 => n291, B1 => E(4), B2 => n288, C1
                           => C(4), C2 => n285, ZN => n20);
   U47 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U48 : AOI22_X1 port map( A1 => A(14), A2 => n280, B1 => B(14), B2 => n277, 
                           ZN => n61);
   U49 : AOI222_X1 port map( A1 => D(14), A2 => n289, B1 => E(14), B2 => n286, 
                           C1 => C(14), C2 => n283, ZN => n62);
   U50 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U51 : AOI22_X1 port map( A1 => A(21), A2 => n281, B1 => B(21), B2 => n278, 
                           ZN => n45);
   U52 : AOI222_X1 port map( A1 => D(21), A2 => n290, B1 => E(21), B2 => n287, 
                           C1 => C(21), C2 => n284, ZN => n46);
   U53 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U54 : AOI22_X1 port map( A1 => A(22), A2 => n281, B1 => B(22), B2 => n278, 
                           ZN => n43);
   U55 : AOI222_X1 port map( A1 => D(22), A2 => n290, B1 => E(22), B2 => n287, 
                           C1 => C(22), C2 => n284, ZN => n44);
   U56 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U57 : AOI22_X1 port map( A1 => A(8), A2 => n282, B1 => B(8), B2 => n279, ZN 
                           => n11);
   U58 : AOI222_X1 port map( A1 => D(8), A2 => n291, B1 => E(8), B2 => n288, C1
                           => C(8), C2 => n285, ZN => n12);
   U59 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U60 : AOI22_X1 port map( A1 => A(5), A2 => n282, B1 => B(5), B2 => n279, ZN 
                           => n17);
   U61 : AOI222_X1 port map( A1 => D(5), A2 => n291, B1 => E(5), B2 => n288, C1
                           => C(5), C2 => n285, ZN => n18);
   U62 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U63 : AOI22_X1 port map( A1 => A(20), A2 => n281, B1 => B(20), B2 => n278, 
                           ZN => n47);
   U64 : AOI222_X1 port map( A1 => D(20), A2 => n290, B1 => E(20), B2 => n287, 
                           C1 => C(20), C2 => n284, ZN => n48);
   U65 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U66 : AOI22_X1 port map( A1 => A(26), A2 => n281, B1 => B(26), B2 => n278, 
                           ZN => n35);
   U67 : AOI222_X1 port map( A1 => D(26), A2 => n290, B1 => E(26), B2 => n287, 
                           C1 => C(26), C2 => n284, ZN => n36);
   U68 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U69 : AOI22_X1 port map( A1 => A(27), A2 => n281, B1 => B(27), B2 => n278, 
                           ZN => n33);
   U70 : AOI222_X1 port map( A1 => D(27), A2 => n290, B1 => E(27), B2 => n287, 
                           C1 => C(27), C2 => n284, ZN => n34);
   U71 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U72 : AOI22_X1 port map( A1 => A(23), A2 => n281, B1 => B(23), B2 => n278, 
                           ZN => n41);
   U73 : AOI222_X1 port map( A1 => D(23), A2 => n290, B1 => E(23), B2 => n287, 
                           C1 => C(23), C2 => n284, ZN => n42);
   U74 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U75 : AOI22_X1 port map( A1 => A(6), A2 => n282, B1 => B(6), B2 => n279, ZN 
                           => n15);
   U76 : AOI222_X1 port map( A1 => D(6), A2 => n291, B1 => E(6), B2 => n288, C1
                           => C(6), C2 => n285, ZN => n16);
   U77 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U78 : AOI22_X1 port map( A1 => A(10), A2 => n280, B1 => B(10), B2 => n277, 
                           ZN => n69);
   U79 : AOI222_X1 port map( A1 => D(10), A2 => n289, B1 => E(10), B2 => n286, 
                           C1 => C(10), C2 => n283, ZN => n70);
   U80 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U81 : AOI22_X1 port map( A1 => A(17), A2 => n280, B1 => B(17), B2 => n277, 
                           ZN => n55);
   U82 : AOI222_X1 port map( A1 => D(17), A2 => n289, B1 => E(17), B2 => n286, 
                           C1 => C(17), C2 => n283, ZN => n56);
   U83 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U84 : AOI22_X1 port map( A1 => A(13), A2 => n280, B1 => B(13), B2 => n277, 
                           ZN => n63);
   U85 : AOI222_X1 port map( A1 => D(13), A2 => n289, B1 => E(13), B2 => n286, 
                           C1 => C(13), C2 => n283, ZN => n64);
   U86 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U87 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U88 : AOI22_X1 port map( A1 => A(7), A2 => n282, B1 => B(7), B2 => n279, ZN 
                           => n13);
   U89 : AOI222_X1 port map( A1 => D(7), A2 => n291, B1 => E(7), B2 => n288, C1
                           => C(7), C2 => n285, ZN => n14);
   U90 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U91 : AOI22_X1 port map( A1 => A(9), A2 => n282, B1 => B(9), B2 => n279, ZN 
                           => n4);
   U92 : AOI222_X1 port map( A1 => D(9), A2 => n291, B1 => E(9), B2 => n288, C1
                           => C(9), C2 => n285, ZN => n5);
   U93 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U94 : AOI22_X1 port map( A1 => A(12), A2 => n280, B1 => B(12), B2 => n277, 
                           ZN => n65);
   U95 : AOI222_X1 port map( A1 => D(12), A2 => n289, B1 => E(12), B2 => n286, 
                           C1 => C(12), C2 => n283, ZN => n66);
   U96 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U97 : AOI22_X1 port map( A1 => A(16), A2 => n280, B1 => B(16), B2 => n277, 
                           ZN => n57);
   U98 : AOI222_X1 port map( A1 => D(16), A2 => n289, B1 => E(16), B2 => n286, 
                           C1 => C(16), C2 => n283, ZN => n58);
   U99 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U100 : AOI22_X1 port map( A1 => A(15), A2 => n280, B1 => B(15), B2 => n277, 
                           ZN => n59);
   U101 : AOI222_X1 port map( A1 => D(15), A2 => n289, B1 => E(15), B2 => n286,
                           C1 => C(15), C2 => n283, ZN => n60);
   U102 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U103 : AOI22_X1 port map( A1 => A(11), A2 => n280, B1 => B(11), B2 => n277, 
                           ZN => n67);
   U104 : AOI222_X1 port map( A1 => D(11), A2 => n289, B1 => E(11), B2 => n286,
                           C1 => C(11), C2 => n283, ZN => n68);
   U105 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U106 : AOI22_X1 port map( A1 => A(3), A2 => n282, B1 => B(3), B2 => n279, ZN
                           => n21);
   U107 : AOI222_X1 port map( A1 => D(3), A2 => n291, B1 => E(3), B2 => n288, 
                           C1 => C(3), C2 => n285, ZN => n22);
   U108 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U109 : AOI22_X1 port map( A1 => A(0), A2 => n280, B1 => B(0), B2 => n277, ZN
                           => n71);
   U110 : AOI222_X1 port map( A1 => D(0), A2 => n289, B1 => E(0), B2 => n286, 
                           C1 => C(0), C2 => n283, ZN => n72);
   U111 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U112 : AOI22_X1 port map( A1 => A(1), A2 => n280, B1 => B(1), B2 => n277, ZN
                           => n49);
   U113 : AOI222_X1 port map( A1 => D(1), A2 => n289, B1 => E(1), B2 => n286, 
                           C1 => C(1), C2 => n283, ZN => n50);
   U114 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U115 : AOI22_X1 port map( A1 => A(2), A2 => n281, B1 => B(2), B2 => n278, ZN
                           => n27);
   U116 : AOI222_X1 port map( A1 => D(2), A2 => n290, B1 => E(2), B2 => n287, 
                           C1 => C(2), C2 => n284, ZN => n28);
   U117 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U118 : AOI22_X1 port map( A1 => A(19), A2 => n280, B1 => B(19), B2 => n277, 
                           ZN => n51);
   U119 : AOI222_X1 port map( A1 => D(19), A2 => n289, B1 => E(19), B2 => n286,
                           C1 => C(19), C2 => n283, ZN => n52);
   U120 : INV_X1 port map( A => Sel(1), ZN => n75);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_7 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_7;

architecture SYN_behav of mux_N32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n325);
   U2 : BUF_X1 port map( A => n10, Z => n326);
   U3 : BUF_X1 port map( A => n10, Z => n327);
   U4 : BUF_X1 port map( A => n6, Z => n337);
   U5 : BUF_X1 port map( A => n6, Z => n338);
   U6 : BUF_X1 port map( A => n9, Z => n328);
   U7 : BUF_X1 port map( A => n9, Z => n329);
   U8 : BUF_X1 port map( A => n7, Z => n334);
   U9 : BUF_X1 port map( A => n7, Z => n335);
   U10 : BUF_X1 port map( A => n8, Z => n331);
   U11 : BUF_X1 port map( A => n8, Z => n332);
   U12 : BUF_X1 port map( A => n9, Z => n330);
   U13 : BUF_X1 port map( A => n7, Z => n336);
   U14 : BUF_X1 port map( A => n8, Z => n333);
   U15 : BUF_X1 port map( A => n6, Z => n339);
   U16 : AND2_X1 port map( A1 => n73, A2 => n74, ZN => n10);
   U17 : AOI222_X1 port map( A1 => n75, A2 => Sel(0), B1 => n76, B2 => Sel(2), 
                           C1 => n74, C2 => Sel(1), ZN => n9);
   U18 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n74, ZN => n7);
   U19 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U20 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n73);
   U21 : INV_X1 port map( A => Sel(0), ZN => n76);
   U22 : INV_X1 port map( A => Sel(2), ZN => n74);
   U23 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U24 : AOI22_X1 port map( A1 => A(16), A2 => n328, B1 => B(16), B2 => n325, 
                           ZN => n57);
   U25 : AOI222_X1 port map( A1 => D(16), A2 => n337, B1 => E(16), B2 => n334, 
                           C1 => C(16), C2 => n331, ZN => n58);
   U26 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U27 : AOI22_X1 port map( A1 => A(2), A2 => n329, B1 => B(2), B2 => n326, ZN 
                           => n27);
   U28 : AOI222_X1 port map( A1 => D(2), A2 => n338, B1 => E(2), B2 => n335, C1
                           => C(2), C2 => n332, ZN => n28);
   U29 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U30 : AOI22_X1 port map( A1 => A(12), A2 => n328, B1 => B(12), B2 => n325, 
                           ZN => n65);
   U31 : AOI222_X1 port map( A1 => D(12), A2 => n337, B1 => E(12), B2 => n334, 
                           C1 => C(12), C2 => n331, ZN => n66);
   U32 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U33 : AOI22_X1 port map( A1 => A(6), A2 => n330, B1 => B(6), B2 => n327, ZN 
                           => n15);
   U34 : AOI222_X1 port map( A1 => D(6), A2 => n339, B1 => E(6), B2 => n336, C1
                           => C(6), C2 => n333, ZN => n16);
   U35 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U36 : AOI22_X1 port map( A1 => A(3), A2 => n330, B1 => B(3), B2 => n327, ZN 
                           => n21);
   U37 : AOI222_X1 port map( A1 => D(3), A2 => n339, B1 => E(3), B2 => n336, C1
                           => C(3), C2 => n333, ZN => n22);
   U38 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U39 : AOI22_X1 port map( A1 => A(10), A2 => n328, B1 => B(10), B2 => n325, 
                           ZN => n69);
   U40 : AOI222_X1 port map( A1 => D(10), A2 => n337, B1 => E(10), B2 => n334, 
                           C1 => C(10), C2 => n331, ZN => n70);
   U41 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n330, B1 => B(4), B2 => n327, ZN 
                           => n19);
   U43 : AOI222_X1 port map( A1 => D(4), A2 => n339, B1 => E(4), B2 => n336, C1
                           => C(4), C2 => n333, ZN => n20);
   U44 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U45 : AOI22_X1 port map( A1 => A(8), A2 => n330, B1 => B(8), B2 => n327, ZN 
                           => n11);
   U46 : AOI222_X1 port map( A1 => D(8), A2 => n339, B1 => E(8), B2 => n336, C1
                           => C(8), C2 => n333, ZN => n12);
   U47 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U48 : AOI22_X1 port map( A1 => A(15), A2 => n328, B1 => B(15), B2 => n325, 
                           ZN => n59);
   U49 : AOI222_X1 port map( A1 => D(15), A2 => n337, B1 => E(15), B2 => n334, 
                           C1 => C(15), C2 => n331, ZN => n60);
   U50 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U51 : AOI22_X1 port map( A1 => A(11), A2 => n328, B1 => B(11), B2 => n325, 
                           ZN => n67);
   U52 : AOI222_X1 port map( A1 => D(11), A2 => n337, B1 => E(11), B2 => n334, 
                           C1 => C(11), C2 => n331, ZN => n68);
   U53 : AND2_X1 port map( A1 => Sel(2), A2 => n73, ZN => n8);
   U54 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n329, B1 => B(25), B2 => n326, 
                           ZN => n37);
   U56 : AOI222_X1 port map( A1 => D(25), A2 => n338, B1 => E(25), B2 => n335, 
                           C1 => C(25), C2 => n332, ZN => n38);
   U57 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U58 : AOI22_X1 port map( A1 => A(26), A2 => n329, B1 => B(26), B2 => n326, 
                           ZN => n35);
   U59 : AOI222_X1 port map( A1 => D(26), A2 => n338, B1 => E(26), B2 => n335, 
                           C1 => C(26), C2 => n332, ZN => n36);
   U60 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U61 : AOI22_X1 port map( A1 => A(22), A2 => n329, B1 => B(22), B2 => n326, 
                           ZN => n43);
   U62 : AOI222_X1 port map( A1 => D(22), A2 => n338, B1 => E(22), B2 => n335, 
                           C1 => C(22), C2 => n332, ZN => n44);
   U63 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n329, B1 => B(27), B2 => n326, 
                           ZN => n33);
   U65 : AOI222_X1 port map( A1 => D(27), A2 => n338, B1 => E(27), B2 => n335, 
                           C1 => C(27), C2 => n332, ZN => n34);
   U66 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U67 : AOI22_X1 port map( A1 => A(19), A2 => n328, B1 => B(19), B2 => n325, 
                           ZN => n51);
   U68 : AOI222_X1 port map( A1 => D(19), A2 => n337, B1 => E(19), B2 => n334, 
                           C1 => C(19), C2 => n331, ZN => n52);
   U69 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U70 : AOI22_X1 port map( A1 => A(28), A2 => n329, B1 => B(28), B2 => n326, 
                           ZN => n31);
   U71 : AOI222_X1 port map( A1 => D(28), A2 => n338, B1 => E(28), B2 => n335, 
                           C1 => C(28), C2 => n332, ZN => n32);
   U72 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U73 : AOI22_X1 port map( A1 => A(29), A2 => n329, B1 => B(29), B2 => n326, 
                           ZN => n29);
   U74 : AOI222_X1 port map( A1 => D(29), A2 => n338, B1 => E(29), B2 => n335, 
                           C1 => C(29), C2 => n332, ZN => n30);
   U75 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U76 : AOI22_X1 port map( A1 => A(5), A2 => n330, B1 => B(5), B2 => n327, ZN 
                           => n17);
   U77 : AOI222_X1 port map( A1 => D(5), A2 => n339, B1 => E(5), B2 => n336, C1
                           => C(5), C2 => n333, ZN => n18);
   U78 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U79 : AOI22_X1 port map( A1 => A(9), A2 => n330, B1 => B(9), B2 => n327, ZN 
                           => n4);
   U80 : AOI222_X1 port map( A1 => D(9), A2 => n339, B1 => E(9), B2 => n336, C1
                           => C(9), C2 => n333, ZN => n5);
   U81 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U82 : AOI22_X1 port map( A1 => A(7), A2 => n330, B1 => B(7), B2 => n327, ZN 
                           => n13);
   U83 : AOI222_X1 port map( A1 => D(7), A2 => n339, B1 => E(7), B2 => n336, C1
                           => C(7), C2 => n333, ZN => n14);
   U84 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U85 : AOI22_X1 port map( A1 => A(13), A2 => n328, B1 => B(13), B2 => n325, 
                           ZN => n63);
   U86 : AOI222_X1 port map( A1 => D(13), A2 => n337, B1 => E(13), B2 => n334, 
                           C1 => C(13), C2 => n331, ZN => n64);
   U87 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U88 : AOI22_X1 port map( A1 => A(17), A2 => n328, B1 => B(17), B2 => n325, 
                           ZN => n55);
   U89 : AOI222_X1 port map( A1 => D(17), A2 => n337, B1 => E(17), B2 => n334, 
                           C1 => C(17), C2 => n331, ZN => n56);
   U90 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U91 : AOI22_X1 port map( A1 => A(14), A2 => n328, B1 => B(14), B2 => n325, 
                           ZN => n61);
   U92 : AOI222_X1 port map( A1 => D(14), A2 => n337, B1 => E(14), B2 => n334, 
                           C1 => C(14), C2 => n331, ZN => n62);
   U93 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U94 : AOI22_X1 port map( A1 => A(23), A2 => n329, B1 => B(23), B2 => n326, 
                           ZN => n41);
   U95 : AOI222_X1 port map( A1 => D(23), A2 => n338, B1 => E(23), B2 => n335, 
                           C1 => C(23), C2 => n332, ZN => n42);
   U96 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U97 : AOI22_X1 port map( A1 => A(24), A2 => n329, B1 => B(24), B2 => n326, 
                           ZN => n39);
   U98 : AOI222_X1 port map( A1 => D(24), A2 => n338, B1 => E(24), B2 => n335, 
                           C1 => C(24), C2 => n332, ZN => n40);
   U99 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U100 : AOI22_X1 port map( A1 => A(20), A2 => n329, B1 => B(20), B2 => n326, 
                           ZN => n47);
   U101 : AOI222_X1 port map( A1 => D(20), A2 => n338, B1 => E(20), B2 => n335,
                           C1 => C(20), C2 => n332, ZN => n48);
   U102 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U103 : AOI22_X1 port map( A1 => A(21), A2 => n329, B1 => B(21), B2 => n326, 
                           ZN => n45);
   U104 : AOI222_X1 port map( A1 => D(21), A2 => n338, B1 => E(21), B2 => n335,
                           C1 => C(21), C2 => n332, ZN => n46);
   U105 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U106 : AOI22_X1 port map( A1 => A(18), A2 => n328, B1 => B(18), B2 => n325, 
                           ZN => n53);
   U107 : AOI222_X1 port map( A1 => D(18), A2 => n337, B1 => E(18), B2 => n334,
                           C1 => C(18), C2 => n331, ZN => n54);
   U108 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U109 : AOI22_X1 port map( A1 => A(30), A2 => n329, B1 => B(30), B2 => n326, 
                           ZN => n25);
   U110 : AOI222_X1 port map( A1 => D(30), A2 => n338, B1 => E(30), B2 => n335,
                           C1 => C(30), C2 => n332, ZN => n26);
   U111 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U112 : AOI22_X1 port map( A1 => A(31), A2 => n330, B1 => B(31), B2 => n327, 
                           ZN => n23);
   U113 : AOI222_X1 port map( A1 => D(31), A2 => n339, B1 => E(31), B2 => n336,
                           C1 => C(31), C2 => n333, ZN => n24);
   U114 : INV_X1 port map( A => Sel(1), ZN => n75);
   U115 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U116 : AOI22_X1 port map( A1 => A(0), A2 => n328, B1 => B(0), B2 => n325, ZN
                           => n71);
   U117 : AOI222_X1 port map( A1 => D(0), A2 => n337, B1 => E(0), B2 => n334, 
                           C1 => C(0), C2 => n331, ZN => n72);
   U118 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U119 : AOI22_X1 port map( A1 => A(1), A2 => n328, B1 => B(1), B2 => n325, ZN
                           => n49);
   U120 : AOI222_X1 port map( A1 => D(1), A2 => n337, B1 => E(1), B2 => n334, 
                           C1 => C(1), C2 => n331, ZN => n50);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_N32_0 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto 0)
         );

end mux_N32_0;

architecture SYN_behav of mux_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286 : std_logic;

begin
   
   U105 : OAI33_X1 port map( A1 => n73, A2 => n75, A3 => n76, B1 => Sel(0), B2 
                           => Sel(2), B3 => Sel(1), ZN => n9);
   U1 : BUF_X1 port map( A => n10, Z => n272);
   U2 : BUF_X1 port map( A => n10, Z => n273);
   U3 : BUF_X1 port map( A => n10, Z => n274);
   U4 : BUF_X1 port map( A => n6, Z => n284);
   U5 : BUF_X1 port map( A => n6, Z => n285);
   U6 : BUF_X1 port map( A => n9, Z => n275);
   U7 : BUF_X1 port map( A => n9, Z => n276);
   U8 : BUF_X1 port map( A => n7, Z => n281);
   U9 : BUF_X1 port map( A => n7, Z => n282);
   U10 : BUF_X1 port map( A => n9, Z => n277);
   U11 : BUF_X1 port map( A => n8, Z => n278);
   U12 : BUF_X1 port map( A => n8, Z => n279);
   U13 : BUF_X1 port map( A => n7, Z => n283);
   U14 : BUF_X1 port map( A => n8, Z => n280);
   U15 : BUF_X1 port map( A => n6, Z => n286);
   U16 : AND2_X1 port map( A1 => n74, A2 => n73, ZN => n10);
   U17 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(1), A3 => n73, ZN => n8);
   U18 : NOR3_X1 port map( A1 => n75, A2 => Sel(2), A3 => n76, ZN => n6);
   U19 : XNOR2_X1 port map( A => n76, B => Sel(1), ZN => n74);
   U20 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => O(14));
   U21 : AOI22_X1 port map( A1 => A(14), A2 => n275, B1 => B(14), B2 => n272, 
                           ZN => n61);
   U22 : AOI222_X1 port map( A1 => D(14), A2 => n284, B1 => C(14), B2 => n281, 
                           C1 => E(14), C2 => n278, ZN => n62);
   U23 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => O(1));
   U24 : AOI22_X1 port map( A1 => A(1), A2 => n275, B1 => B(1), B2 => n272, ZN 
                           => n49);
   U25 : AOI222_X1 port map( A1 => D(1), A2 => n284, B1 => C(1), B2 => n281, C1
                           => E(1), C2 => n278, ZN => n50);
   U26 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => O(10));
   U27 : AOI22_X1 port map( A1 => A(10), A2 => n275, B1 => B(10), B2 => n272, 
                           ZN => n69);
   U28 : AOI222_X1 port map( A1 => D(10), A2 => n284, B1 => C(10), B2 => n281, 
                           C1 => E(10), C2 => n278, ZN => n70);
   U29 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => O(4));
   U30 : AOI22_X1 port map( A1 => A(4), A2 => n277, B1 => B(4), B2 => n274, ZN 
                           => n19);
   U31 : AOI222_X1 port map( A1 => D(4), A2 => n286, B1 => C(4), B2 => n283, C1
                           => E(4), C2 => n280, ZN => n20);
   U32 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => O(0));
   U33 : AOI22_X1 port map( A1 => A(0), A2 => n275, B1 => B(0), B2 => n272, ZN 
                           => n71);
   U34 : AOI222_X1 port map( A1 => D(0), A2 => n284, B1 => C(0), B2 => n281, C1
                           => E(0), C2 => n278, ZN => n72);
   U35 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => O(8));
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n277, B1 => B(8), B2 => n274, ZN 
                           => n11);
   U37 : AOI222_X1 port map( A1 => D(8), A2 => n286, B1 => C(8), B2 => n283, C1
                           => E(8), C2 => n280, ZN => n12);
   U38 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => O(2));
   U39 : AOI22_X1 port map( A1 => A(2), A2 => n276, B1 => B(2), B2 => n273, ZN 
                           => n27);
   U40 : AOI222_X1 port map( A1 => D(2), A2 => n285, B1 => C(2), B2 => n282, C1
                           => E(2), C2 => n279, ZN => n28);
   U41 : INV_X1 port map( A => Sel(2), ZN => n73);
   U42 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => O(13));
   U43 : AOI22_X1 port map( A1 => A(13), A2 => n275, B1 => B(13), B2 => n272, 
                           ZN => n63);
   U44 : AOI222_X1 port map( A1 => D(13), A2 => n284, B1 => C(13), B2 => n281, 
                           C1 => E(13), C2 => n278, ZN => n64);
   U45 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => O(9));
   U46 : AOI22_X1 port map( A1 => A(9), A2 => n277, B1 => B(9), B2 => n274, ZN 
                           => n4);
   U47 : AOI222_X1 port map( A1 => D(9), A2 => n286, B1 => C(9), B2 => n283, C1
                           => E(9), C2 => n280, ZN => n5);
   U48 : AND2_X1 port map( A1 => Sel(2), A2 => n74, ZN => n7);
   U49 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => O(3));
   U50 : AOI22_X1 port map( A1 => A(3), A2 => n277, B1 => B(3), B2 => n274, ZN 
                           => n21);
   U51 : AOI222_X1 port map( A1 => D(3), A2 => n286, B1 => C(3), B2 => n283, C1
                           => E(3), C2 => n280, ZN => n22);
   U52 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => O(7));
   U53 : AOI22_X1 port map( A1 => A(7), A2 => n277, B1 => B(7), B2 => n274, ZN 
                           => n13);
   U54 : AOI222_X1 port map( A1 => D(7), A2 => n286, B1 => C(7), B2 => n283, C1
                           => E(7), C2 => n280, ZN => n14);
   U55 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => O(15));
   U56 : AOI22_X1 port map( A1 => A(15), A2 => n275, B1 => B(15), B2 => n272, 
                           ZN => n59);
   U57 : AOI222_X1 port map( A1 => D(15), A2 => n284, B1 => C(15), B2 => n281, 
                           C1 => E(15), C2 => n278, ZN => n60);
   U58 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => O(11));
   U59 : AOI22_X1 port map( A1 => A(11), A2 => n275, B1 => B(11), B2 => n272, 
                           ZN => n67);
   U60 : AOI222_X1 port map( A1 => D(11), A2 => n284, B1 => C(11), B2 => n281, 
                           C1 => E(11), C2 => n278, ZN => n68);
   U61 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => O(12));
   U62 : AOI22_X1 port map( A1 => A(12), A2 => n275, B1 => B(12), B2 => n272, 
                           ZN => n65);
   U63 : AOI222_X1 port map( A1 => D(12), A2 => n284, B1 => C(12), B2 => n281, 
                           C1 => E(12), C2 => n278, ZN => n66);
   U64 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => O(6));
   U65 : AOI22_X1 port map( A1 => A(6), A2 => n277, B1 => B(6), B2 => n274, ZN 
                           => n15);
   U66 : AOI222_X1 port map( A1 => D(6), A2 => n286, B1 => C(6), B2 => n283, C1
                           => E(6), C2 => n280, ZN => n16);
   U67 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => O(24));
   U68 : AOI22_X1 port map( A1 => A(24), A2 => n276, B1 => B(24), B2 => n273, 
                           ZN => n39);
   U69 : AOI222_X1 port map( A1 => D(24), A2 => n285, B1 => C(24), B2 => n282, 
                           C1 => E(24), C2 => n279, ZN => n40);
   U70 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => O(20));
   U71 : AOI22_X1 port map( A1 => A(20), A2 => n276, B1 => B(20), B2 => n273, 
                           ZN => n47);
   U72 : AOI222_X1 port map( A1 => D(20), A2 => n285, B1 => C(20), B2 => n282, 
                           C1 => E(20), C2 => n279, ZN => n48);
   U73 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => O(25));
   U74 : AOI22_X1 port map( A1 => A(25), A2 => n276, B1 => B(25), B2 => n273, 
                           ZN => n37);
   U75 : AOI222_X1 port map( A1 => D(25), A2 => n285, B1 => C(25), B2 => n282, 
                           C1 => E(25), C2 => n279, ZN => n38);
   U76 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => O(21));
   U77 : AOI22_X1 port map( A1 => A(21), A2 => n276, B1 => B(21), B2 => n273, 
                           ZN => n45);
   U78 : AOI222_X1 port map( A1 => D(21), A2 => n285, B1 => C(21), B2 => n282, 
                           C1 => E(21), C2 => n279, ZN => n46);
   U79 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => O(17));
   U80 : AOI22_X1 port map( A1 => A(17), A2 => n275, B1 => B(17), B2 => n272, 
                           ZN => n55);
   U81 : AOI222_X1 port map( A1 => D(17), A2 => n284, B1 => C(17), B2 => n281, 
                           C1 => E(17), C2 => n278, ZN => n56);
   U82 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => O(26));
   U83 : AOI22_X1 port map( A1 => A(26), A2 => n276, B1 => B(26), B2 => n273, 
                           ZN => n35);
   U84 : AOI222_X1 port map( A1 => D(26), A2 => n285, B1 => C(26), B2 => n282, 
                           C1 => E(26), C2 => n279, ZN => n36);
   U85 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => O(22));
   U86 : AOI22_X1 port map( A1 => A(22), A2 => n276, B1 => B(22), B2 => n273, 
                           ZN => n43);
   U87 : AOI222_X1 port map( A1 => D(22), A2 => n285, B1 => C(22), B2 => n282, 
                           C1 => E(22), C2 => n279, ZN => n44);
   U88 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => O(18));
   U89 : AOI22_X1 port map( A1 => A(18), A2 => n275, B1 => B(18), B2 => n272, 
                           ZN => n53);
   U90 : AOI222_X1 port map( A1 => D(18), A2 => n284, B1 => C(18), B2 => n281, 
                           C1 => E(18), C2 => n278, ZN => n54);
   U91 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => O(27));
   U92 : AOI22_X1 port map( A1 => A(27), A2 => n276, B1 => B(27), B2 => n273, 
                           ZN => n33);
   U93 : AOI222_X1 port map( A1 => D(27), A2 => n285, B1 => C(27), B2 => n282, 
                           C1 => E(27), C2 => n279, ZN => n34);
   U94 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => O(23));
   U95 : AOI22_X1 port map( A1 => A(23), A2 => n276, B1 => B(23), B2 => n273, 
                           ZN => n41);
   U96 : AOI222_X1 port map( A1 => D(23), A2 => n285, B1 => C(23), B2 => n282, 
                           C1 => E(23), C2 => n279, ZN => n42);
   U97 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => O(19));
   U98 : AOI22_X1 port map( A1 => A(19), A2 => n275, B1 => B(19), B2 => n272, 
                           ZN => n51);
   U99 : AOI222_X1 port map( A1 => D(19), A2 => n284, B1 => C(19), B2 => n281, 
                           C1 => E(19), C2 => n278, ZN => n52);
   U100 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => O(28));
   U101 : AOI22_X1 port map( A1 => A(28), A2 => n276, B1 => B(28), B2 => n273, 
                           ZN => n31);
   U102 : AOI222_X1 port map( A1 => D(28), A2 => n285, B1 => C(28), B2 => n282,
                           C1 => E(28), C2 => n279, ZN => n32);
   U103 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => O(29));
   U104 : AOI22_X1 port map( A1 => A(29), A2 => n276, B1 => B(29), B2 => n273, 
                           ZN => n29);
   U106 : AOI222_X1 port map( A1 => D(29), A2 => n285, B1 => C(29), B2 => n282,
                           C1 => E(29), C2 => n279, ZN => n30);
   U107 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => O(30));
   U108 : AOI22_X1 port map( A1 => A(30), A2 => n276, B1 => B(30), B2 => n273, 
                           ZN => n25);
   U109 : AOI222_X1 port map( A1 => D(30), A2 => n285, B1 => C(30), B2 => n282,
                           C1 => E(30), C2 => n279, ZN => n26);
   U110 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => O(31));
   U111 : AOI22_X1 port map( A1 => A(31), A2 => n277, B1 => B(31), B2 => n274, 
                           ZN => n23);
   U112 : AOI222_X1 port map( A1 => D(31), A2 => n286, B1 => C(31), B2 => n283,
                           C1 => E(31), C2 => n280, ZN => n24);
   U113 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => O(16));
   U114 : AOI22_X1 port map( A1 => A(16), A2 => n275, B1 => B(16), B2 => n272, 
                           ZN => n57);
   U115 : AOI222_X1 port map( A1 => D(16), A2 => n284, B1 => C(16), B2 => n281,
                           C1 => E(16), C2 => n278, ZN => n58);
   U116 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => O(5));
   U117 : AOI22_X1 port map( A1 => A(5), A2 => n277, B1 => B(5), B2 => n274, ZN
                           => n17);
   U118 : AOI222_X1 port map( A1 => D(5), A2 => n286, B1 => C(5), B2 => n283, 
                           C1 => E(5), C2 => n280, ZN => n18);
   U119 : INV_X1 port map( A => Sel(1), ZN => n75);
   U120 : INV_X1 port map( A => Sel(0), ZN => n76);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S14 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S14;

architecture SYN_struct of shift_mul_N16_S14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_31_port, E_30_port, E_29_port, E_28_port, E_27_port,
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, n9, n10, n12, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n62, n63, 
      D_21_port, n65, D_23_port, n67, D_25_port, n69, D_27_port, n71, n72 : 
      std_logic;

begin
   B <= ( A(15), A(15), A(15), A(14), A(13), D_27_port, A(11), D_25_port, A(9),
      D_23_port, A(7), D_21_port, A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   C <= ( E_31_port, E_31_port, E_30_port, E_29_port, E_28_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   D <= ( A(15), A(15), A(14), A(13), D_27_port, A(11), D_25_port, A(9), 
      D_23_port, A(7), D_21_port, A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port );
   E <= ( E_31_port, E_30_port, E_29_port, E_28_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n12, B => A(13), Z => E_28_port);
   U28 : XOR2_X1 port map( A => n14, B => n71, Z => E_27_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_26_port);
   U30 : XOR2_X1 port map( A => n17, B => n69, Z => E_25_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_24_port);
   U32 : XOR2_X1 port map( A => n20, B => n67, Z => E_23_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_22_port);
   U34 : XOR2_X1 port map( A => n23, B => n65, Z => E_21_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_20_port);
   U36 : XOR2_X1 port map( A => n26, B => n63, Z => E_19_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_18_port);
   U38 : XOR2_X1 port map( A => n29, B => n62, Z => E_17_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_16_port);
   U2 : INV_X1 port map( A => n9, ZN => E_31_port);
   U3 : OAI21_X1 port map( B1 => n10, B2 => n72, A => n9, ZN => E_30_port);
   U4 : NAND2_X1 port map( A1 => n14, A2 => n71, ZN => n12);
   U5 : NAND2_X1 port map( A1 => n17, A2 => n69, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n72, A2 => n10, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n26, A2 => n63, ZN => n25);
   U8 : NAND2_X1 port map( A1 => n20, A2 => n67, ZN => n19);
   U9 : NAND2_X1 port map( A1 => n23, A2 => n65, ZN => n22);
   U10 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U11 : XNOR2_X1 port map( A => A(14), B => n13, ZN => E_29_port);
   U12 : NOR2_X1 port map( A1 => A(13), A2 => n12, ZN => n13);
   U13 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U14 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U15 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U16 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U18 : INV_X1 port map( A => A(8), ZN => n67);
   U19 : INV_X1 port map( A => A(12), ZN => n71);
   U20 : INV_X1 port map( A => A(10), ZN => n69);
   U21 : INV_X1 port map( A => A(6), ZN => n65);
   U22 : INV_X1 port map( A => A(4), ZN => n63);
   U23 : INV_X1 port map( A => A(15), ZN => n72);
   U24 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n12, ZN => n10);
   U25 : NAND2_X1 port map( A1 => n29, A2 => n62, ZN => n28);
   U26 : INV_X1 port map( A => A(2), ZN => n62);
   U40 : INV_X1 port map( A => n65, ZN => D_21_port);
   U41 : INV_X1 port map( A => n67, ZN => D_23_port);
   U42 : INV_X1 port map( A => n69, ZN => D_25_port);
   U43 : INV_X1 port map( A => n71, ZN => D_27_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S12 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S12;

architecture SYN_struct of shift_mul_N16_S12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_28_port, E_27_port, E_26_port, E_25_port, E_24_port,
      E_23_port, E_22_port, E_21_port, E_20_port, E_19_port, E_18_port, 
      E_17_port, E_16_port, E_15_port, E_14_port, E_29_port, n9, n10, n11, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n66, n67, n68, 
      D_21_port, n70, n71, D_25_port, n73, n74, D_28_port : std_logic;

begin
   B <= ( D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), 
      D_25_port, A(11), A(10), A(9), D_21_port, A(7), A(6), A(5), A(4), A(3), 
      A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_29_port, E_29_port, E_29_port, E_29_port, E_28_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), D_25_port, 
      A(11), A(10), A(9), D_21_port, A(7), A(6), A(5), A(4), A(3), A(2), A(1), 
      A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_29_port, E_29_port, E_29_port, E_28_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U25 : NAND3_X1 port map( A1 => n11, A2 => n74, A3 => D_28_port, ZN => n10);
   U26 : XOR2_X1 port map( A => n11, B => n74, Z => E_27_port);
   U27 : XOR2_X1 port map( A => n13, B => A(13), Z => E_26_port);
   U28 : XOR2_X1 port map( A => n14, B => n73, Z => E_25_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_24_port);
   U30 : XOR2_X1 port map( A => n17, B => n71, Z => E_23_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_22_port);
   U32 : XOR2_X1 port map( A => n20, B => n70, Z => E_21_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_20_port);
   U34 : XOR2_X1 port map( A => n23, B => n68, Z => E_19_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_18_port);
   U36 : XOR2_X1 port map( A => n26, B => n67, Z => E_17_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_16_port);
   U38 : XOR2_X1 port map( A => n29, B => n66, Z => E_15_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_14_port);
   U2 : AOI21_X1 port map( B1 => n74, B2 => n11, A => D_28_port, ZN => 
                           E_29_port);
   U3 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => E_28_port);
   U4 : INV_X1 port map( A => E_29_port, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n17, A2 => n71, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n26, A2 => n67, ZN => n25);
   U7 : NAND2_X1 port map( A1 => n20, A2 => n70, ZN => n19);
   U8 : NAND2_X1 port map( A1 => n23, A2 => n68, ZN => n22);
   U9 : NAND2_X1 port map( A1 => n14, A2 => n73, ZN => n13);
   U10 : NOR2_X1 port map( A1 => n13, A2 => A(13), ZN => n11);
   U11 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U12 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U13 : BUF_X1 port map( A => A(15), Z => D_28_port);
   U14 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U15 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U16 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U18 : INV_X1 port map( A => A(8), ZN => n70);
   U19 : INV_X1 port map( A => A(12), ZN => n73);
   U20 : INV_X1 port map( A => A(10), ZN => n71);
   U21 : INV_X1 port map( A => A(6), ZN => n68);
   U22 : INV_X1 port map( A => A(4), ZN => n67);
   U23 : NAND2_X1 port map( A1 => n29, A2 => n66, ZN => n28);
   U24 : INV_X1 port map( A => A(2), ZN => n66);
   U40 : INV_X1 port map( A => n70, ZN => D_21_port);
   U41 : INV_X1 port map( A => n73, ZN => D_25_port);
   U42 : INV_X1 port map( A => A(14), ZN => n74);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S10 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S10;

architecture SYN_struct of shift_mul_N16_S10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port,
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_26_port, E_27_port, n9, n10, n12, n13,
      n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29, n81, n82, n83, n84
      , n85, n86, D_26_port, n88 : std_logic;

begin
   B <= ( D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, 
      D_26_port, A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), 
      A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, 
      E_26_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, D_26_port, 
      A(14), A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), 
      A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_27_port, E_27_port, E_27_port, E_27_port, E_27_port, E_26_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n12, B => A(13), Z => E_24_port);
   U28 : XOR2_X1 port map( A => n14, B => n86, Z => E_23_port);
   U29 : XOR2_X1 port map( A => n16, B => A(11), Z => E_22_port);
   U30 : XOR2_X1 port map( A => n17, B => n85, Z => E_21_port);
   U31 : XOR2_X1 port map( A => n19, B => A(9), Z => E_20_port);
   U32 : XOR2_X1 port map( A => n20, B => n84, Z => E_19_port);
   U33 : XOR2_X1 port map( A => n22, B => A(7), Z => E_18_port);
   U34 : XOR2_X1 port map( A => n23, B => n83, Z => E_17_port);
   U35 : XOR2_X1 port map( A => n25, B => A(5), Z => E_16_port);
   U36 : XOR2_X1 port map( A => n26, B => n82, Z => E_15_port);
   U37 : XOR2_X1 port map( A => n28, B => A(3), Z => E_14_port);
   U38 : XOR2_X1 port map( A => n29, B => n81, Z => E_13_port);
   U39 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_12_port);
   U2 : INV_X1 port map( A => n9, ZN => E_27_port);
   U3 : INV_X1 port map( A => n88, ZN => D_26_port);
   U4 : OAI21_X1 port map( B1 => n10, B2 => n88, A => n9, ZN => E_26_port);
   U5 : NAND2_X1 port map( A1 => n14, A2 => n86, ZN => n12);
   U6 : NAND2_X1 port map( A1 => n17, A2 => n85, ZN => n16);
   U7 : NAND2_X1 port map( A1 => n88, A2 => n10, ZN => n9);
   U8 : NAND2_X1 port map( A1 => n26, A2 => n82, ZN => n25);
   U9 : NAND2_X1 port map( A1 => n20, A2 => n84, ZN => n19);
   U10 : NAND2_X1 port map( A1 => n23, A2 => n83, ZN => n22);
   U11 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n29);
   U12 : XNOR2_X1 port map( A => A(14), B => n13, ZN => E_25_port);
   U13 : NOR2_X1 port map( A1 => A(13), A2 => n12, ZN => n13);
   U14 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n17);
   U15 : NOR2_X1 port map( A1 => n28, A2 => A(3), ZN => n26);
   U16 : NOR2_X1 port map( A1 => n22, A2 => A(7), ZN => n20);
   U17 : NOR2_X1 port map( A1 => n25, A2 => A(5), ZN => n23);
   U18 : NOR2_X1 port map( A1 => n16, A2 => A(11), ZN => n14);
   U19 : INV_X1 port map( A => A(8), ZN => n84);
   U20 : INV_X1 port map( A => A(12), ZN => n86);
   U21 : INV_X1 port map( A => A(10), ZN => n85);
   U22 : INV_X1 port map( A => A(6), ZN => n83);
   U23 : INV_X1 port map( A => A(4), ZN => n82);
   U24 : INV_X1 port map( A => A(15), ZN => n88);
   U25 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n12, ZN => n10);
   U26 : NAND2_X1 port map( A1 => n29, A2 => n81, ZN => n28);
   U40 : INV_X1 port map( A => A(2), ZN => n81);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S8 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S8;

architecture SYN_struct of shift_mul_N16_S8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_23_port, E_22_port, E_21_port, E_20_port, E_19_port,
      E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, E_13_port, 
      E_12_port, E_11_port, E_10_port, E_25_port, E_24_port, n7, n8, n9, n11, 
      n13, n15, n17, n18, n19, n21, n22, n24, n25, n95, n96, D_11_port, n98, 
      D_13_port, n100, D_15_port, n102, D_20_port, n104, D_23_port, n106, 
      D_24_port, B_27_port : std_logic;

begin
   B <= ( B_27_port, B_27_port, B_27_port, B_27_port, B_27_port, D_24_port, 
      D_24_port, D_24_port, D_24_port, D_23_port, A(13), A(12), D_20_port, 
      A(10), A(9), A(8), A(7), D_15_port, A(5), D_13_port, A(3), D_11_port, 
      A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   C <= ( E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, 
      E_25_port, E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   D <= ( D_24_port, D_24_port, D_24_port, D_24_port, D_24_port, D_24_port, 
      D_24_port, D_24_port, D_23_port, A(13), A(12), D_20_port, A(10), A(9), 
      A(8), A(7), D_15_port, A(5), D_13_port, A(3), D_11_port, A(1), A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, E_25_port, 
      E_25_port, E_24_port, E_23_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U29 : NAND3_X1 port map( A1 => n9, A2 => n106, A3 => B_27_port, ZN => n8);
   U31 : XOR2_X1 port map( A => n11, B => A(12), Z => E_21_port);
   U33 : XOR2_X1 port map( A => n15, B => A(9), Z => E_18_port);
   U34 : XOR2_X1 port map( A => n17, B => A(7), Z => E_16_port);
   U35 : XOR2_X1 port map( A => n21, B => A(5), Z => E_14_port);
   U36 : XOR2_X1 port map( A => n24, B => A(3), Z => E_12_port);
   U37 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_10_port);
   U2 : AOI21_X2 port map( B1 => n106, B2 => n9, A => B_27_port, ZN => 
                           E_25_port);
   U3 : XNOR2_X1 port map( A => n9, B => D_23_port, ZN => E_23_port);
   U4 : XNOR2_X1 port map( A => n13, B => D_20_port, ZN => E_20_port);
   U5 : XNOR2_X1 port map( A => n22, B => D_13_port, ZN => E_13_port);
   U6 : XNOR2_X1 port map( A => n25, B => D_11_port, ZN => E_11_port);
   U7 : XNOR2_X1 port map( A => n19, B => D_15_port, ZN => E_15_port);
   U8 : NAND2_X1 port map( A1 => n13, A2 => n104, ZN => n11);
   U9 : NAND2_X1 port map( A1 => n19, A2 => n102, ZN => n17);
   U10 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => E_24_port);
   U11 : INV_X1 port map( A => E_25_port, ZN => n7);
   U12 : NAND2_X1 port map( A1 => n22, A2 => n100, ZN => n21);
   U13 : NOR3_X1 port map( A1 => A(12), A2 => A(13), A3 => n11, ZN => n9);
   U14 : XNOR2_X1 port map( A => n95, B => A(13), ZN => E_22_port);
   U15 : NOR2_X1 port map( A1 => n11, A2 => A(12), ZN => n95);
   U16 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n15, ZN => n13);
   U17 : XNOR2_X1 port map( A => n96, B => A(10), ZN => E_19_port);
   U18 : NOR2_X1 port map( A1 => n15, A2 => A(9), ZN => n96);
   U19 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n25);
   U20 : BUF_X1 port map( A => A(15), Z => D_24_port);
   U21 : XNOR2_X1 port map( A => A(8), B => n18, ZN => E_17_port);
   U22 : NOR2_X1 port map( A1 => A(7), A2 => n17, ZN => n18);
   U23 : NOR2_X1 port map( A1 => n24, A2 => A(3), ZN => n22);
   U24 : NOR2_X1 port map( A1 => n21, A2 => A(5), ZN => n19);
   U25 : BUF_X1 port map( A => A(15), Z => B_27_port);
   U26 : NAND2_X1 port map( A1 => n25, A2 => n98, ZN => n24);
   U27 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n17, ZN => n15);
   U28 : INV_X1 port map( A => n98, ZN => D_11_port);
   U30 : INV_X1 port map( A => A(2), ZN => n98);
   U32 : INV_X1 port map( A => n100, ZN => D_13_port);
   U38 : INV_X1 port map( A => A(4), ZN => n100);
   U39 : INV_X1 port map( A => n102, ZN => D_15_port);
   U40 : INV_X1 port map( A => A(6), ZN => n102);
   U41 : INV_X1 port map( A => n104, ZN => D_20_port);
   U42 : INV_X1 port map( A => A(11), ZN => n104);
   U43 : INV_X1 port map( A => n106, ZN => D_23_port);
   U44 : INV_X1 port map( A => A(14), ZN => n106);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S6 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S6;

architecture SYN_struct of shift_mul_N16_S6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_21_port, E_20_port, E_19_port, E_18_port, E_17_port,
      E_16_port, E_15_port, E_14_port, E_13_port, E_12_port, E_11_port, 
      E_10_port, E_9_port, E_8_port, E_23_port, E_22_port, n4, n6, n7, n9, n10,
      n11, n13, n15, n16, n17, n19, n20, n87, n88, n89, n90, E_26_port, 
      E_30_port, C_31_port, C_30_port, C_24_port, C_28_port, C_22_port, 
      C_26_port, E_27_port, D_18_port, n101, n102, D_22_port, B_23_port : 
      std_logic;

begin
   B <= ( B_23_port, B_23_port, B_23_port, B_23_port, B_23_port, B_23_port, 
      B_23_port, B_23_port, B_23_port, D_22_port, D_22_port, A(14), A(13), 
      A(12), D_18_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), 
      A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   C <= ( C_31_port, C_30_port, C_24_port, C_28_port, C_22_port, C_26_port, 
      E_26_port, C_24_port, C_28_port, C_22_port, E_22_port, E_21_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   D <= ( D_22_port, D_22_port, D_22_port, D_22_port, D_22_port, D_22_port, 
      D_22_port, D_22_port, D_22_port, D_22_port, A(14), A(13), A(12), 
      D_18_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), 
      A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port );
   E <= ( C_26_port, E_30_port, E_26_port, E_27_port, E_27_port, E_26_port, 
      E_30_port, C_31_port, C_30_port, E_22_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, A(0), 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U24 : XOR2_X1 port map( A => n4, B => A(2), Z => E_9_port);
   U25 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_8_port);
   U26 : NAND3_X1 port map( A1 => n7, A2 => n102, A3 => B_23_port, ZN => n6);
   U27 : XOR2_X1 port map( A => n9, B => A(13), Z => E_20_port);
   U28 : XOR2_X1 port map( A => n10, B => A(12), Z => E_19_port);
   U30 : XOR2_X1 port map( A => n13, B => A(9), Z => E_16_port);
   U31 : XOR2_X1 port map( A => n15, B => A(7), Z => E_14_port);
   U33 : XOR2_X1 port map( A => n17, B => A(5), Z => E_12_port);
   U34 : XOR2_X1 port map( A => n19, B => A(3), Z => E_10_port);
   U2 : AOI21_X1 port map( B1 => n102, B2 => n7, A => B_23_port, ZN => 
                           E_23_port);
   U3 : XNOR2_X1 port map( A => n7, B => A(14), ZN => E_21_port);
   U4 : XNOR2_X1 port map( A => n11, B => D_18_port, ZN => E_18_port);
   U5 : NAND2_X1 port map( A1 => n11, A2 => n101, ZN => n10);
   U6 : NAND2_X1 port map( A1 => n90, A2 => n6, ZN => E_22_port);
   U7 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n13, ZN => n11);
   U8 : XNOR2_X1 port map( A => n87, B => A(10), ZN => E_17_port);
   U9 : NOR2_X1 port map( A1 => n13, A2 => A(9), ZN => n87);
   U10 : XNOR2_X1 port map( A => n88, B => A(6), ZN => E_13_port);
   U11 : NOR2_X1 port map( A1 => n17, A2 => A(5), ZN => n88);
   U12 : NOR2_X1 port map( A1 => n9, A2 => A(13), ZN => n7);
   U13 : BUF_X1 port map( A => A(15), Z => D_22_port);
   U14 : XNOR2_X1 port map( A => A(8), B => n16, ZN => E_15_port);
   U15 : NOR2_X1 port map( A1 => A(7), A2 => n15, ZN => n16);
   U16 : BUF_X1 port map( A => A(15), Z => B_23_port);
   U17 : XNOR2_X1 port map( A => A(4), B => n20, ZN => E_11_port);
   U18 : NOR2_X1 port map( A1 => A(3), A2 => n19, ZN => n20);
   U19 : OR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n19, ZN => n17);
   U20 : OR3_X1 port map( A1 => A(5), A2 => A(6), A3 => n17, ZN => n15);
   U21 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n15, ZN => n13);
   U22 : OR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n4);
   U23 : OR2_X1 port map( A1 => n10, A2 => A(12), ZN => n9);
   U29 : OR2_X1 port map( A1 => n4, A2 => A(2), ZN => n19);
   U32 : INV_X1 port map( A => E_23_port, ZN => n89);
   U35 : INV_X1 port map( A => E_23_port, ZN => n90);
   U36 : INV_X1 port map( A => n89, ZN => E_26_port);
   U37 : INV_X1 port map( A => n89, ZN => E_30_port);
   U38 : INV_X1 port map( A => n89, ZN => C_31_port);
   U39 : INV_X1 port map( A => n89, ZN => C_30_port);
   U40 : INV_X1 port map( A => n90, ZN => C_24_port);
   U41 : INV_X1 port map( A => n90, ZN => C_28_port);
   U42 : INV_X1 port map( A => n90, ZN => C_22_port);
   U43 : INV_X1 port map( A => n90, ZN => C_26_port);
   U44 : INV_X1 port map( A => n89, ZN => E_27_port);
   U45 : INV_X1 port map( A => n101, ZN => D_18_port);
   U46 : INV_X1 port map( A => A(11), ZN => n101);
   U47 : INV_X1 port map( A => A(14), ZN => n102);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S4 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S4;

architecture SYN_struct of shift_mul_N16_S4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_20_port, E_19_port, E_18_port, E_17_port, E_16_port,
      E_15_port, E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, 
      E_9_port, E_8_port, E_7_port, E_6_port, E_23_port, E_21_port, n6, n7, n8,
      n10, n12, n13, n14, n15, n16, n19, n21, n22, n24, n25, n105, n106, n107, 
      n108, n109, D_19_port, n111, D_20_port, B_19_port, n114 : std_logic;

begin
   B <= ( B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, 
      B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, B_19_port, 
      B_19_port, D_19_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6),
      A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   C <= ( E_21_port, E_21_port, E_21_port, E_21_port, E_23_port, E_23_port, 
      E_21_port, E_21_port, E_23_port, E_23_port, E_23_port, E_23_port, 
      E_20_port, E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   D <= ( D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, 
      D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, D_20_port, 
      D_19_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4)
      , A(3), A(2), A(1), A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   E <= ( E_23_port, E_23_port, E_23_port, E_21_port, E_23_port, E_23_port, 
      E_23_port, E_23_port, E_23_port, E_21_port, E_21_port, E_20_port, 
      E_19_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, A(0), X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U26 : XOR2_X1 port map( A => n6, B => A(4), Z => E_9_port);
   U27 : XOR2_X1 port map( A => n7, B => A(3), Z => E_8_port);
   U28 : XOR2_X1 port map( A => n8, B => n107, Z => E_7_port);
   U29 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_6_port);
   U30 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n114, ZN => n13);
   U32 : XOR2_X1 port map( A => A(12), B => n16, Z => E_17_port);
   U33 : XOR2_X1 port map( A => n15, B => n109, Z => E_16_port);
   U35 : XOR2_X1 port map( A => n19, B => A(9), Z => E_14_port);
   U36 : XOR2_X1 port map( A => n21, B => A(8), Z => E_13_port);
   U37 : XOR2_X1 port map( A => n22, B => n108, Z => E_12_port);
   U38 : XOR2_X1 port map( A => n24, B => A(5), Z => E_10_port);
   U2 : AOI21_X1 port map( B1 => n15, B2 => n14, A => n114, ZN => E_21_port);
   U3 : AOI21_X2 port map( B1 => n10, B2 => n111, A => n114, ZN => E_23_port);
   U4 : XNOR2_X1 port map( A => n10, B => D_19_port, ZN => E_19_port);
   U5 : NAND2_X1 port map( A1 => n15, A2 => n109, ZN => n16);
   U6 : NAND2_X1 port map( A1 => n22, A2 => n108, ZN => n21);
   U7 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => E_20_port);
   U8 : INV_X1 port map( A => E_21_port, ZN => n12);
   U9 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n19, ZN => n15);
   U10 : NOR3_X1 port map( A1 => A(12), A2 => A(13), A3 => n16, ZN => n10);
   U11 : NOR4_X1 port map( A1 => A(11), A2 => A(12), A3 => A(13), A4 => 
                           D_19_port, ZN => n14);
   U12 : XNOR2_X1 port map( A => n105, B => A(13), ZN => E_18_port);
   U13 : NOR2_X1 port map( A1 => n16, A2 => A(12), ZN => n105);
   U14 : XNOR2_X1 port map( A => n106, B => A(10), ZN => E_15_port);
   U15 : NOR2_X1 port map( A1 => n19, A2 => A(9), ZN => n106);
   U16 : NOR3_X1 port map( A1 => A(5), A2 => A(6), A3 => n24, ZN => n22);
   U17 : BUF_X1 port map( A => A(15), Z => B_19_port);
   U18 : BUF_X1 port map( A => A(15), Z => D_20_port);
   U19 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n8);
   U20 : XNOR2_X1 port map( A => A(6), B => n25, ZN => E_11_port);
   U21 : NOR2_X1 port map( A1 => A(5), A2 => n24, ZN => n25);
   U22 : INV_X1 port map( A => A(7), ZN => n108);
   U23 : INV_X1 port map( A => A(11), ZN => n109);
   U24 : OR2_X1 port map( A1 => n6, A2 => A(4), ZN => n24);
   U25 : OR2_X1 port map( A1 => n21, A2 => A(8), ZN => n19);
   U31 : BUF_X1 port map( A => A(15), Z => n114);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n107, ZN => n7);
   U39 : OR2_X1 port map( A1 => n7, A2 => A(3), ZN => n6);
   U40 : INV_X1 port map( A => A(2), ZN => n107);
   U41 : INV_X1 port map( A => n111, ZN => D_19_port);
   U42 : INV_X1 port map( A => A(14), ZN => n111);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S2 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S2;

architecture SYN_struct of shift_mul_N16_S2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port,
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, C_22_port, n7, n8, n9, n11, n12, n15, n16, 
      n17, n18, n19, n20, n21, n23, n24, n26, n27, n28, E_23_port, n118, n119, 
      n120, D_13_port, n122, D_15_port, n124, D_18_port, D_30_port, B_29_port :
      std_logic;

begin
   B <= ( B_29_port, B_29_port, B_29_port, B_29_port, B_29_port, D_30_port, 
      D_30_port, D_30_port, D_30_port, D_30_port, D_30_port, D_30_port, 
      D_30_port, D_30_port, D_30_port, A(14), A(13), D_15_port, A(11), 
      D_13_port, A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port, X_Logic0_port );
   C <= ( C_22_port, E_23_port, C_22_port, C_22_port, C_22_port, C_22_port, 
      C_22_port, E_23_port, C_22_port, C_22_port, E_23_port, E_23_port, 
      C_22_port, E_23_port, E_18_port, E_17_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, E_5_port, E_4_port, A(0), X_Logic0_port, 
      X_Logic0_port );
   D <= ( D_30_port, D_30_port, D_18_port, D_18_port, D_18_port, D_18_port, 
      D_18_port, D_18_port, D_18_port, D_18_port, D_18_port, D_18_port, 
      D_18_port, D_18_port, A(14), A(13), D_15_port, A(11), D_13_port, A(9), 
      A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   E <= ( C_22_port, C_22_port, E_23_port, C_22_port, E_23_port, E_23_port, 
      E_23_port, E_23_port, E_23_port, E_23_port, E_23_port, E_23_port, 
      E_23_port, E_18_port, E_17_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, A(0), X_Logic0_port, X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U27 : XOR2_X1 port map( A => n7, B => A(6), Z => E_9_port);
   U28 : XOR2_X1 port map( A => n8, B => A(5), Z => E_8_port);
   U29 : XOR2_X1 port map( A => n9, B => n120, Z => E_7_port);
   U30 : XOR2_X1 port map( A => n11, B => A(3), Z => E_6_port);
   U31 : XOR2_X1 port map( A => n12, B => n119, Z => E_5_port);
   U32 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_4_port);
   U33 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => B_29_port, ZN => n15);
   U34 : XOR2_X1 port map( A => n20, B => A(13), Z => E_16_port);
   U35 : XOR2_X1 port map( A => n124, B => n21, Z => E_15_port);
   U36 : XOR2_X1 port map( A => n23, B => A(11), Z => E_14_port);
   U37 : XOR2_X1 port map( A => n122, B => n24, Z => E_13_port);
   U38 : XOR2_X1 port map( A => n26, B => A(9), Z => E_12_port);
   U39 : XOR2_X1 port map( A => n27, B => A(7), Z => E_10_port);
   U2 : INV_X1 port map( A => n118, ZN => E_23_port);
   U3 : INV_X1 port map( A => C_22_port, ZN => n118);
   U4 : AOI21_X1 port map( B1 => n17, B2 => n16, A => B_29_port, ZN => 
                           C_22_port);
   U5 : NAND2_X1 port map( A1 => n118, A2 => n15, ZN => E_18_port);
   U6 : INV_X1 port map( A => n16, ZN => n26);
   U7 : NAND2_X1 port map( A1 => n24, A2 => n122, ZN => n23);
   U8 : NAND2_X1 port map( A1 => n21, A2 => n124, ZN => n20);
   U9 : NAND2_X1 port map( A1 => n9, A2 => n120, ZN => n8);
   U10 : NOR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n27, ZN => n16);
   U11 : NOR4_X1 port map( A1 => A(11), A2 => D_15_port, A3 => D_13_port, A4 =>
                           n18, ZN => n17);
   U12 : OR3_X1 port map( A1 => A(13), A2 => A(9), A3 => A(14), ZN => n18);
   U13 : BUF_X1 port map( A => A(15), Z => D_18_port);
   U14 : BUF_X1 port map( A => A(15), Z => D_30_port);
   U15 : XNOR2_X1 port map( A => A(8), B => n28, ZN => E_11_port);
   U16 : NOR2_X1 port map( A1 => A(7), A2 => n27, ZN => n28);
   U17 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n12);
   U18 : XNOR2_X1 port map( A => A(14), B => n19, ZN => E_17_port);
   U19 : NOR2_X1 port map( A1 => A(13), A2 => n20, ZN => n19);
   U20 : NOR2_X1 port map( A1 => n26, A2 => A(9), ZN => n24);
   U21 : NOR2_X1 port map( A1 => n11, A2 => A(3), ZN => n9);
   U22 : NOR2_X1 port map( A1 => n23, A2 => A(11), ZN => n21);
   U23 : INV_X1 port map( A => A(12), ZN => n124);
   U24 : INV_X1 port map( A => A(10), ZN => n122);
   U25 : BUF_X1 port map( A => A(15), Z => B_29_port);
   U26 : INV_X1 port map( A => A(4), ZN => n120);
   U40 : OR2_X1 port map( A1 => n7, A2 => A(6), ZN => n27);
   U41 : NAND2_X1 port map( A1 => n12, A2 => n119, ZN => n11);
   U42 : OR2_X1 port map( A1 => n8, A2 => A(5), ZN => n7);
   U43 : INV_X1 port map( A => A(2), ZN => n119);
   U44 : INV_X1 port map( A => n122, ZN => D_13_port);
   U45 : INV_X1 port map( A => n124, ZN => D_15_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shift_mul_N16_S0 is

   port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
         std_logic_vector (31 downto 0));

end shift_mul_N16_S0;

architecture SYN_struct of shift_mul_N16_S0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, E_16_port, E_15_port, E_14_port, E_13_port, E_12_port,
      E_11_port, E_10_port, E_9_port, E_8_port, E_7_port, E_6_port, E_5_port, 
      E_3_port, E_2_port, net25272, E_4_port, n6, n8, n9, n10, n11, n12, n13, 
      n14, n16, n18, n19, n21, n22, n99, n100, C_20_port, D_3_port, n103, n104,
      D_12_port, n106, D_28_port, n108 : std_logic;

begin
   B <= ( A(15), D_28_port, D_28_port, D_28_port, A(15), D_28_port, D_28_port, 
      D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, D_28_port, 
      D_28_port, D_28_port, D_28_port, D_28_port, A(14), A(13), A(12), 
      D_12_port, A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), D_3_port, 
      A(1), A(0) );
   C <= ( C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, E_16_port, E_15_port, 
      E_14_port, E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port
      , E_7_port, E_6_port, E_5_port, E_4_port, E_3_port, E_2_port, A(0) );
   D <= ( D_28_port, D_28_port, D_28_port, D_28_port, A(15), D_28_port, A(15), 
      D_28_port, A(15), D_28_port, A(15), D_28_port, A(15), D_28_port, A(15), 
      D_28_port, A(14), A(13), A(12), D_12_port, A(10), A(9), A(8), A(7), A(6),
      A(5), A(4), A(3), D_3_port, A(1), A(0), X_Logic0_port );
   E <= ( C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, C_20_port, 
      C_20_port, C_20_port, C_20_port, E_16_port, E_15_port, E_14_port, 
      E_13_port, E_12_port, E_11_port, E_10_port, E_9_port, E_8_port, E_7_port,
      E_6_port, E_5_port, E_4_port, E_3_port, E_2_port, A(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U29 : XOR2_X1 port map( A => n8, B => A(7), Z => E_8_port);
   U30 : XOR2_X1 port map( A => n9, B => A(6), Z => E_7_port);
   U31 : XOR2_X1 port map( A => n12, B => A(3), Z => E_4_port);
   U32 : XOR2_X1 port map( A => A(1), B => A(0), Z => E_2_port);
   U34 : XOR2_X1 port map( A => n16, B => A(13), Z => E_14_port);
   U35 : XOR2_X1 port map( A => n18, B => A(12), Z => E_13_port);
   U36 : XOR2_X1 port map( A => n21, B => A(9), Z => E_10_port);
   U2 : BUF_X2 port map( A => net25272, Z => C_20_port);
   U3 : INV_X1 port map( A => n6, ZN => net25272);
   U4 : INV_X1 port map( A => n108, ZN => D_28_port);
   U5 : XNOR2_X1 port map( A => n19, B => D_12_port, ZN => E_12_port);
   U6 : XNOR2_X1 port map( A => n10, B => A(5), ZN => E_6_port);
   U7 : XNOR2_X1 port map( A => n13, B => D_3_port, ZN => E_3_port);
   U8 : OAI21_X1 port map( B1 => n14, B2 => n108, A => n6, ZN => E_16_port);
   U9 : NAND2_X1 port map( A1 => n10, A2 => n104, ZN => n9);
   U10 : NAND2_X1 port map( A1 => n19, A2 => n106, ZN => n18);
   U11 : NAND2_X1 port map( A1 => n108, A2 => n14, ZN => n6);
   U12 : NOR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n12, ZN => n10);
   U13 : NOR3_X1 port map( A1 => A(10), A2 => A(9), A3 => n21, ZN => n19);
   U14 : XNOR2_X1 port map( A => n99, B => A(8), ZN => E_9_port);
   U15 : NOR2_X1 port map( A1 => n8, A2 => A(7), ZN => n99);
   U16 : XNOR2_X1 port map( A => n100, B => A(14), ZN => E_15_port);
   U17 : NOR2_X1 port map( A1 => n16, A2 => A(13), ZN => n100);
   U18 : NOR2_X1 port map( A1 => A(1), A2 => A(0), ZN => n13);
   U19 : XNOR2_X1 port map( A => A(10), B => n22, ZN => E_11_port);
   U20 : NOR2_X1 port map( A1 => A(9), A2 => n21, ZN => n22);
   U21 : XNOR2_X1 port map( A => A(4), B => n11, ZN => E_5_port);
   U22 : NOR2_X1 port map( A1 => A(3), A2 => n12, ZN => n11);
   U23 : NAND2_X1 port map( A1 => n13, A2 => n103, ZN => n12);
   U24 : OR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n8, ZN => n21);
   U25 : OR3_X1 port map( A1 => A(13), A2 => A(14), A3 => n16, ZN => n14);
   U26 : OR2_X1 port map( A1 => n18, A2 => A(12), ZN => n16);
   U27 : OR2_X1 port map( A1 => n9, A2 => A(6), ZN => n8);
   U28 : INV_X1 port map( A => n103, ZN => D_3_port);
   U33 : INV_X1 port map( A => A(2), ZN => n103);
   U37 : INV_X1 port map( A => A(5), ZN => n104);
   U38 : INV_X1 port map( A => n106, ZN => D_12_port);
   U39 : INV_X1 port map( A => A(11), ZN => n106);
   U40 : INV_X1 port map( A => A(15), ZN => n108);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity cla_adder_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end cla_adder_N32_0;

architecture SYN_struct of cla_adder_N32_0 is

   component sum_generator_Nbits32_Nblocks8_0
      port( A, B : in std_logic_vector (31 downto 0);  Carry : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_Nblocks8_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic_vector (8 downto 0));
   end component;
   
   signal Carry_8_port, Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port,
      Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port : std_logic;

begin
   
   CG : carry_generator_N32_Nblocks8_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci, Cout(8) => 
                           Carry_8_port, Cout(7) => Carry_7_port, Cout(6) => 
                           Carry_6_port, Cout(5) => Carry_5_port, Cout(4) => 
                           Carry_4_port, Cout(3) => Carry_3_port, Cout(2) => 
                           Carry_2_port, Cout(1) => Carry_1_port, Cout(0) => 
                           Carry_0_port);
   SG : sum_generator_Nbits32_Nblocks8_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Carry(8) => Carry_8_port, 
                           Carry(7) => Carry_7_port, Carry(6) => Carry_6_port, 
                           Carry(5) => Carry_5_port, Carry(4) => Carry_4_port, 
                           Carry(3) => Carry_3_port, Carry(2) => Carry_2_port, 
                           Carry(1) => Carry_1_port, Carry(0) => Carry_0_port, 
                           S(31) => Sum(31), S(30) => Sum(30), S(29) => Sum(29)
                           , S(28) => Sum(28), S(27) => Sum(27), S(26) => 
                           Sum(26), S(25) => Sum(25), S(24) => Sum(24), S(23) 
                           => Sum(23), S(22) => Sum(22), S(21) => Sum(21), 
                           S(20) => Sum(20), S(19) => Sum(19), S(18) => Sum(18)
                           , S(17) => Sum(17), S(16) => Sum(16), S(15) => 
                           Sum(15), S(14) => Sum(14), S(13) => Sum(13), S(12) 
                           => Sum(12), S(11) => Sum(11), S(10) => Sum(10), S(9)
                           => Sum(9), S(8) => Sum(8), S(7) => Sum(7), S(6) => 
                           Sum(6), S(5) => Sum(5), S(4) => Sum(4), S(3) => 
                           Sum(3), S(2) => Sum(2), S(1) => Sum(1), S(0) => 
                           Sum(0), Cout => Cout);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity generic_xor_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end generic_xor_N32;

architecture SYN_struct of generic_xor_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component xor_gate_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component xor_gate_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   X_gate_0 : xor_gate_0 port map( A => A(0), B => n3, Y => Y(0));
   X_gate_1 : xor_gate_31 port map( A => A(1), B => n1, Y => Y(1));
   X_gate_2 : xor_gate_30 port map( A => A(2), B => n1, Y => Y(2));
   X_gate_3 : xor_gate_29 port map( A => A(3), B => n1, Y => Y(3));
   X_gate_4 : xor_gate_28 port map( A => A(4), B => n1, Y => Y(4));
   X_gate_5 : xor_gate_27 port map( A => A(5), B => n1, Y => Y(5));
   X_gate_6 : xor_gate_26 port map( A => A(6), B => n1, Y => Y(6));
   X_gate_7 : xor_gate_25 port map( A => A(7), B => n1, Y => Y(7));
   X_gate_8 : xor_gate_24 port map( A => A(8), B => n1, Y => Y(8));
   X_gate_9 : xor_gate_23 port map( A => A(9), B => n1, Y => Y(9));
   X_gate_10 : xor_gate_22 port map( A => A(10), B => n1, Y => Y(10));
   X_gate_11 : xor_gate_21 port map( A => A(11), B => n1, Y => Y(11));
   X_gate_12 : xor_gate_20 port map( A => A(12), B => n1, Y => Y(12));
   X_gate_13 : xor_gate_19 port map( A => A(13), B => n2, Y => Y(13));
   X_gate_14 : xor_gate_18 port map( A => A(14), B => n2, Y => Y(14));
   X_gate_15 : xor_gate_17 port map( A => A(15), B => n2, Y => Y(15));
   X_gate_16 : xor_gate_16 port map( A => A(16), B => n2, Y => Y(16));
   X_gate_17 : xor_gate_15 port map( A => A(17), B => n2, Y => Y(17));
   X_gate_18 : xor_gate_14 port map( A => A(18), B => n2, Y => Y(18));
   X_gate_19 : xor_gate_13 port map( A => A(19), B => n2, Y => Y(19));
   X_gate_20 : xor_gate_12 port map( A => A(20), B => n2, Y => Y(20));
   X_gate_21 : xor_gate_11 port map( A => A(21), B => n2, Y => Y(21));
   X_gate_22 : xor_gate_10 port map( A => A(22), B => n2, Y => Y(22));
   X_gate_23 : xor_gate_9 port map( A => A(23), B => n2, Y => Y(23));
   X_gate_24 : xor_gate_8 port map( A => A(24), B => n2, Y => Y(24));
   X_gate_25 : xor_gate_7 port map( A => A(25), B => n3, Y => Y(25));
   X_gate_26 : xor_gate_6 port map( A => A(26), B => n3, Y => Y(26));
   X_gate_27 : xor_gate_5 port map( A => A(27), B => n3, Y => Y(27));
   X_gate_28 : xor_gate_4 port map( A => A(28), B => n3, Y => Y(28));
   X_gate_29 : xor_gate_3 port map( A => A(29), B => n3, Y => Y(29));
   X_gate_30 : xor_gate_2 port map( A => A(30), B => n3, Y => Y(30));
   X_gate_31 : xor_gate_1 port map( A => A(31), B => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : BUF_X1 port map( A => B, Z => n2);
   U3 : BUF_X1 port map( A => B, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity mux_alu is

   port( addsub, mul, log, shift, lhi : in std_logic_vector (31 downto 0);  gt,
         get, lt, let, eq, neq : in std_logic;  sel : in std_logic_vector (0 to
         4);  out_mux : out std_logic_vector (31 downto 0));

end mux_alu;

architecture SYN_behav of mux_alu is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n2, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n144 : std_logic;

begin
   
   U128 : OAI33_X1 port map( A1 => n101, A2 => n30, A3 => n102, B1 => n103, B2 
                           => sel(0), B3 => sel(2), ZN => n16);
   out_mux_tri_0_inst : TBUF_X1 port map( A => n153, EN => n119, Z => 
                           out_mux(0));
   out_mux_tri_1_inst : TBUF_X1 port map( A => n152, EN => n119, Z => 
                           out_mux(1));
   out_mux_tri_2_inst : TBUF_X1 port map( A => n151, EN => n119, Z => 
                           out_mux(2));
   out_mux_tri_3_inst : TBUF_X1 port map( A => n150, EN => n119, Z => 
                           out_mux(3));
   out_mux_tri_4_inst : TBUF_X1 port map( A => n149, EN => n119, Z => 
                           out_mux(4));
   out_mux_tri_5_inst : TBUF_X1 port map( A => n148, EN => n119, Z => 
                           out_mux(5));
   out_mux_tri_6_inst : TBUF_X1 port map( A => n147, EN => n119, Z => 
                           out_mux(6));
   out_mux_tri_7_inst : TBUF_X1 port map( A => n146, EN => n119, Z => 
                           out_mux(7));
   out_mux_tri_8_inst : TBUF_X1 port map( A => n145, EN => n119, Z => 
                           out_mux(8));
   out_mux_tri_9_inst : TBUF_X1 port map( A => n143, EN => n119, Z => 
                           out_mux(9));
   out_mux_tri_10_inst : TBUF_X1 port map( A => n142, EN => n119, Z => 
                           out_mux(10));
   out_mux_tri_11_inst : TBUF_X1 port map( A => n141, EN => n119, Z => 
                           out_mux(11));
   out_mux_tri_12_inst : TBUF_X1 port map( A => n140, EN => n120, Z => 
                           out_mux(12));
   out_mux_tri_13_inst : TBUF_X1 port map( A => n139, EN => n120, Z => 
                           out_mux(13));
   out_mux_tri_14_inst : TBUF_X1 port map( A => n138, EN => n120, Z => 
                           out_mux(14));
   out_mux_tri_15_inst : TBUF_X1 port map( A => n137, EN => n120, Z => 
                           out_mux(15));
   out_mux_tri_16_inst : TBUF_X1 port map( A => n136, EN => n120, Z => 
                           out_mux(16));
   out_mux_tri_17_inst : TBUF_X1 port map( A => n135, EN => n120, Z => 
                           out_mux(17));
   out_mux_tri_18_inst : TBUF_X1 port map( A => n134, EN => n120, Z => 
                           out_mux(18));
   out_mux_tri_19_inst : TBUF_X1 port map( A => n133, EN => n120, Z => 
                           out_mux(19));
   out_mux_tri_20_inst : TBUF_X1 port map( A => n132, EN => n120, Z => 
                           out_mux(20));
   out_mux_tri_21_inst : TBUF_X1 port map( A => n131, EN => n120, Z => 
                           out_mux(21));
   out_mux_tri_22_inst : TBUF_X1 port map( A => n130, EN => n120, Z => 
                           out_mux(22));
   out_mux_tri_23_inst : TBUF_X1 port map( A => n129, EN => n120, Z => 
                           out_mux(23));
   out_mux_tri_24_inst : TBUF_X1 port map( A => n128, EN => n144, Z => 
                           out_mux(24));
   out_mux_tri_25_inst : TBUF_X1 port map( A => n127, EN => n144, Z => 
                           out_mux(25));
   out_mux_tri_26_inst : TBUF_X1 port map( A => n126, EN => n144, Z => 
                           out_mux(26));
   out_mux_tri_27_inst : TBUF_X1 port map( A => n125, EN => n144, Z => 
                           out_mux(27));
   out_mux_tri_28_inst : TBUF_X1 port map( A => n124, EN => n144, Z => 
                           out_mux(28));
   out_mux_tri_29_inst : TBUF_X1 port map( A => n123, EN => n144, Z => 
                           out_mux(29));
   out_mux_tri_30_inst : TBUF_X1 port map( A => n122, EN => n144, Z => 
                           out_mux(30));
   out_mux_tri_31_inst : TBUF_X1 port map( A => n121, EN => n144, Z => 
                           out_mux(31));
   U2 : BUF_X1 port map( A => n38, Z => n104);
   U3 : BUF_X1 port map( A => n38, Z => n105);
   U4 : BUF_X1 port map( A => n38, Z => n106);
   U5 : NOR3_X1 port map( A1 => n30, A2 => n25, A3 => n101, ZN => n38);
   U6 : BUF_X1 port map( A => n17, Z => n113);
   U7 : BUF_X1 port map( A => n17, Z => n114);
   U8 : BUF_X1 port map( A => n37, Z => n107);
   U9 : BUF_X1 port map( A => n37, Z => n108);
   U10 : BUF_X1 port map( A => n16, Z => n116);
   U11 : BUF_X1 port map( A => n16, Z => n117);
   U12 : BUF_X1 port map( A => n36, Z => n110);
   U13 : BUF_X1 port map( A => n36, Z => n111);
   U14 : BUF_X1 port map( A => n16, Z => n118);
   U15 : BUF_X1 port map( A => n36, Z => n112);
   U16 : AOI22_X1 port map( A1 => n24, A2 => gt, B1 => n25, B2 => let, ZN => 
                           n23);
   U17 : BUF_X1 port map( A => n2, Z => n120);
   U18 : BUF_X1 port map( A => n2, Z => n119);
   U19 : INV_X1 port map( A => n102, ZN => n25);
   U20 : BUF_X1 port map( A => n2, Z => n144);
   U21 : BUF_X1 port map( A => n17, Z => n115);
   U22 : NAND2_X1 port map( A1 => n10, A2 => n12, ZN => n101);
   U23 : BUF_X1 port map( A => n37, Z => n109);
   U24 : INV_X1 port map( A => n24, ZN => n13);
   U25 : INV_X1 port map( A => n35, ZN => n29);
   U26 : AOI22_X1 port map( A1 => get, A2 => n25, B1 => n26, B2 => gt, ZN => 
                           n35);
   U27 : NAND2_X1 port map( A1 => sel(1), A2 => n28, ZN => n103);
   U28 : NOR4_X1 port map( A1 => n13, A2 => n12, A3 => n30, A4 => sel(1), ZN =>
                           n17);
   U29 : NOR4_X1 port map( A1 => n101, A2 => n25, A3 => n24, A4 => sel(2), ZN 
                           => n36);
   U30 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n127);
   U31 : AOI22_X1 port map( A1 => log(25), A2 => n104, B1 => addsub(25), B2 => 
                           n110, ZN => n87);
   U32 : AOI222_X1 port map( A1 => mul(25), A2 => n108, B1 => shift(25), B2 => 
                           n116, C1 => lhi(25), C2 => n114, ZN => n88);
   U33 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => n128);
   U34 : AOI22_X1 port map( A1 => log(24), A2 => n104, B1 => addsub(24), B2 => 
                           n110, ZN => n85);
   U35 : AOI222_X1 port map( A1 => mul(24), A2 => n108, B1 => shift(24), B2 => 
                           n116, C1 => lhi(24), C2 => n114, ZN => n86);
   U36 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => n129);
   U37 : AOI22_X1 port map( A1 => log(23), A2 => n104, B1 => addsub(23), B2 => 
                           n110, ZN => n83);
   U38 : AOI222_X1 port map( A1 => mul(23), A2 => n108, B1 => shift(23), B2 => 
                           n116, C1 => lhi(23), C2 => n114, ZN => n84);
   U39 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n130);
   U40 : AOI22_X1 port map( A1 => log(22), A2 => n104, B1 => addsub(22), B2 => 
                           n110, ZN => n81);
   U41 : AOI222_X1 port map( A1 => mul(22), A2 => n108, B1 => shift(22), B2 => 
                           n116, C1 => lhi(22), C2 => n114, ZN => n82);
   U42 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n131);
   U43 : AOI22_X1 port map( A1 => log(21), A2 => n104, B1 => addsub(21), B2 => 
                           n110, ZN => n79);
   U44 : AOI222_X1 port map( A1 => mul(21), A2 => n108, B1 => shift(21), B2 => 
                           n116, C1 => lhi(21), C2 => n114, ZN => n80);
   U45 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n132);
   U46 : AOI22_X1 port map( A1 => log(20), A2 => n104, B1 => addsub(20), B2 => 
                           n110, ZN => n77);
   U47 : AOI222_X1 port map( A1 => mul(20), A2 => n108, B1 => shift(20), B2 => 
                           n116, C1 => lhi(20), C2 => n114, ZN => n78);
   U48 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => n133);
   U49 : AOI22_X1 port map( A1 => log(19), A2 => n105, B1 => addsub(19), B2 => 
                           n111, ZN => n75);
   U50 : AOI222_X1 port map( A1 => mul(19), A2 => n108, B1 => shift(19), B2 => 
                           n117, C1 => lhi(19), C2 => n114, ZN => n76);
   U51 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => n134);
   U52 : AOI22_X1 port map( A1 => log(18), A2 => n105, B1 => addsub(18), B2 => 
                           n111, ZN => n73);
   U53 : AOI222_X1 port map( A1 => mul(18), A2 => n108, B1 => shift(18), B2 => 
                           n117, C1 => lhi(18), C2 => n114, ZN => n74);
   U54 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n135);
   U55 : AOI22_X1 port map( A1 => log(17), A2 => n105, B1 => addsub(17), B2 => 
                           n111, ZN => n71);
   U56 : AOI222_X1 port map( A1 => mul(17), A2 => n108, B1 => shift(17), B2 => 
                           n117, C1 => lhi(17), C2 => n114, ZN => n72);
   U57 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => n136);
   U58 : AOI22_X1 port map( A1 => log(16), A2 => n105, B1 => addsub(16), B2 => 
                           n111, ZN => n69);
   U59 : AOI222_X1 port map( A1 => mul(16), A2 => n108, B1 => shift(16), B2 => 
                           n117, C1 => lhi(16), C2 => n114, ZN => n70);
   U60 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => n137);
   U61 : AOI22_X1 port map( A1 => log(15), A2 => n105, B1 => addsub(15), B2 => 
                           n111, ZN => n67);
   U62 : AOI222_X1 port map( A1 => mul(15), A2 => n108, B1 => shift(15), B2 => 
                           n117, C1 => lhi(15), C2 => n114, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => n138);
   U64 : AOI22_X1 port map( A1 => log(14), A2 => n105, B1 => addsub(14), B2 => 
                           n111, ZN => n65);
   U65 : AOI222_X1 port map( A1 => mul(14), A2 => n108, B1 => shift(14), B2 => 
                           n117, C1 => lhi(14), C2 => n114, ZN => n66);
   U66 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n139);
   U67 : AOI22_X1 port map( A1 => log(13), A2 => n105, B1 => addsub(13), B2 => 
                           n111, ZN => n63);
   U68 : AOI222_X1 port map( A1 => mul(13), A2 => n108, B1 => shift(13), B2 => 
                           n117, C1 => lhi(13), C2 => n114, ZN => n64);
   U69 : NOR3_X1 port map( A1 => n102, A2 => sel(2), A3 => n101, ZN => n37);
   U70 : NOR2_X1 port map( A1 => sel(3), A2 => sel(4), ZN => n24);
   U71 : AOI21_X1 port map( B1 => n10, B2 => n11, A => n12, ZN => n2);
   U72 : NAND2_X1 port map( A1 => sel(2), A2 => n13, ZN => n11);
   U73 : NOR2_X1 port map( A1 => n28, A2 => sel(4), ZN => n26);
   U74 : INV_X1 port map( A => sel(2), ZN => n30);
   U75 : AOI21_X1 port map( B1 => n26, B2 => lt, A => n27, ZN => n22);
   U76 : AND3_X1 port map( A1 => get, A2 => n28, A3 => sel(4), ZN => n27);
   U77 : AOI21_X1 port map( B1 => n32, B2 => n33, A => n30, ZN => n31);
   U78 : AOI21_X1 port map( B1 => eq, B2 => n26, A => n34, ZN => n33);
   U79 : AOI22_X1 port map( A1 => neq, A2 => n25, B1 => n24, B2 => lt, ZN => 
                           n32);
   U80 : AND3_X1 port map( A1 => let, A2 => n28, A3 => sel(4), ZN => n34);
   U81 : INV_X1 port map( A => sel(0), ZN => n12);
   U82 : OAI21_X1 port map( B1 => n19, B2 => n10, A => n20, ZN => n18);
   U83 : INV_X1 port map( A => n21, ZN => n20);
   U84 : AOI21_X1 port map( B1 => n29, B2 => n30, A => n31, ZN => n19);
   U85 : AOI211_X1 port map( C1 => n22, C2 => n23, A => sel(2), B => n12, ZN =>
                           n21);
   U86 : NAND2_X1 port map( A1 => sel(3), A2 => sel(4), ZN => n102);
   U87 : INV_X1 port map( A => sel(3), ZN => n28);
   U88 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n153);
   U89 : AOI222_X1 port map( A1 => addsub(0), A2 => n112, B1 => mul(0), B2 => 
                           n107, C1 => log(0), C2 => n106, ZN => n14);
   U90 : AOI221_X1 port map( B1 => shift(0), B2 => n118, C1 => lhi(0), C2 => 
                           n113, A => n18, ZN => n15);
   U91 : INV_X1 port map( A => sel(1), ZN => n10);
   U92 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => n146);
   U93 : AOI22_X1 port map( A1 => log(7), A2 => n106, B1 => addsub(7), B2 => 
                           n112, ZN => n51);
   U94 : AOI222_X1 port map( A1 => mul(7), A2 => n107, B1 => shift(7), B2 => 
                           n118, C1 => lhi(7), C2 => n113, ZN => n52);
   U95 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n147);
   U96 : AOI22_X1 port map( A1 => log(6), A2 => n106, B1 => addsub(6), B2 => 
                           n112, ZN => n49);
   U97 : AOI222_X1 port map( A1 => mul(6), A2 => n107, B1 => shift(6), B2 => 
                           n118, C1 => lhi(6), C2 => n113, ZN => n50);
   U98 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => n148);
   U99 : AOI22_X1 port map( A1 => log(5), A2 => n106, B1 => addsub(5), B2 => 
                           n112, ZN => n47);
   U100 : AOI222_X1 port map( A1 => mul(5), A2 => n107, B1 => shift(5), B2 => 
                           n118, C1 => lhi(5), C2 => n113, ZN => n48);
   U101 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n149);
   U102 : AOI22_X1 port map( A1 => log(4), A2 => n106, B1 => addsub(4), B2 => 
                           n112, ZN => n45);
   U103 : AOI222_X1 port map( A1 => mul(4), A2 => n107, B1 => shift(4), B2 => 
                           n118, C1 => lhi(4), C2 => n113, ZN => n46);
   U104 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n150);
   U105 : AOI22_X1 port map( A1 => log(3), A2 => n106, B1 => addsub(3), B2 => 
                           n112, ZN => n43);
   U106 : AOI222_X1 port map( A1 => mul(3), A2 => n107, B1 => shift(3), B2 => 
                           n118, C1 => lhi(3), C2 => n113, ZN => n44);
   U107 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n151);
   U108 : AOI22_X1 port map( A1 => log(2), A2 => n106, B1 => addsub(2), B2 => 
                           n112, ZN => n41);
   U109 : AOI222_X1 port map( A1 => mul(2), A2 => n107, B1 => shift(2), B2 => 
                           n118, C1 => lhi(2), C2 => n113, ZN => n42);
   U110 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n152);
   U111 : AOI22_X1 port map( A1 => log(1), A2 => n106, B1 => addsub(1), B2 => 
                           n112, ZN => n39);
   U112 : AOI222_X1 port map( A1 => mul(1), A2 => n107, B1 => shift(1), B2 => 
                           n118, C1 => lhi(1), C2 => n113, ZN => n40);
   U113 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n121);
   U114 : AOI22_X1 port map( A1 => log(31), A2 => n104, B1 => addsub(31), B2 =>
                           n110, ZN => n99);
   U115 : AOI222_X1 port map( A1 => mul(31), A2 => n109, B1 => shift(31), B2 =>
                           n116, C1 => lhi(31), C2 => n115, ZN => n100);
   U116 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n122);
   U117 : AOI22_X1 port map( A1 => log(30), A2 => n104, B1 => addsub(30), B2 =>
                           n110, ZN => n97);
   U118 : AOI222_X1 port map( A1 => mul(30), A2 => n109, B1 => shift(30), B2 =>
                           n116, C1 => lhi(30), C2 => n115, ZN => n98);
   U119 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n123);
   U120 : AOI22_X1 port map( A1 => log(29), A2 => n104, B1 => addsub(29), B2 =>
                           n110, ZN => n95);
   U121 : AOI222_X1 port map( A1 => mul(29), A2 => n109, B1 => shift(29), B2 =>
                           n116, C1 => lhi(29), C2 => n115, ZN => n96);
   U122 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => n124);
   U123 : AOI22_X1 port map( A1 => log(28), A2 => n104, B1 => addsub(28), B2 =>
                           n110, ZN => n93);
   U124 : AOI222_X1 port map( A1 => mul(28), A2 => n109, B1 => shift(28), B2 =>
                           n116, C1 => lhi(28), C2 => n115, ZN => n94);
   U125 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => n125);
   U126 : AOI22_X1 port map( A1 => log(27), A2 => n104, B1 => addsub(27), B2 =>
                           n110, ZN => n91);
   U127 : AOI222_X1 port map( A1 => mul(27), A2 => n109, B1 => shift(27), B2 =>
                           n116, C1 => lhi(27), C2 => n115, ZN => n92);
   U129 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n126);
   U130 : AOI22_X1 port map( A1 => log(26), A2 => n104, B1 => addsub(26), B2 =>
                           n110, ZN => n89);
   U131 : AOI222_X1 port map( A1 => mul(26), A2 => n109, B1 => shift(26), B2 =>
                           n116, C1 => lhi(26), C2 => n115, ZN => n90);
   U132 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n140);
   U133 : AOI22_X1 port map( A1 => log(12), A2 => n105, B1 => addsub(12), B2 =>
                           n111, ZN => n61);
   U134 : AOI222_X1 port map( A1 => mul(12), A2 => n107, B1 => shift(12), B2 =>
                           n117, C1 => lhi(12), C2 => n113, ZN => n62);
   U135 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => n141);
   U136 : AOI22_X1 port map( A1 => log(11), A2 => n105, B1 => addsub(11), B2 =>
                           n111, ZN => n59);
   U137 : AOI222_X1 port map( A1 => mul(11), A2 => n107, B1 => shift(11), B2 =>
                           n117, C1 => lhi(11), C2 => n113, ZN => n60);
   U138 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n142);
   U139 : AOI22_X1 port map( A1 => log(10), A2 => n105, B1 => addsub(10), B2 =>
                           n111, ZN => n57);
   U140 : AOI222_X1 port map( A1 => mul(10), A2 => n107, B1 => shift(10), B2 =>
                           n117, C1 => lhi(10), C2 => n113, ZN => n58);
   U141 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n143);
   U142 : AOI22_X1 port map( A1 => log(9), A2 => n105, B1 => addsub(9), B2 => 
                           n111, ZN => n55);
   U143 : AOI222_X1 port map( A1 => mul(9), A2 => n107, B1 => shift(9), B2 => 
                           n117, C1 => lhi(9), C2 => n113, ZN => n56);
   U144 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n145);
   U145 : AOI22_X1 port map( A1 => log(8), A2 => n105, B1 => addsub(8), B2 => 
                           n111, ZN => n53);
   U146 : AOI222_X1 port map( A1 => mul(8), A2 => n107, B1 => shift(8), B2 => 
                           n117, C1 => lhi(8), C2 => n113, ZN => n54);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity comparator is

   port( C : in std_logic;  Sum : in std_logic_vector (31 downto 0);  sign : in
         std_logic;  gt, get, lt, let, eq, neq : out std_logic);

end comparator;

architecture SYN_behav of comparator is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal gt_port, get_port, lt_port, eq_port, n4, n5, n6, n7, n8, n9, n10, n11
      , n12, n13 : std_logic;

begin
   gt <= gt_port;
   get <= get_port;
   lt <= lt_port;
   eq <= eq_port;
   
   U16 : XOR2_X1 port map( A => sign, B => C, Z => get_port);
   U1 : INV_X1 port map( A => gt_port, ZN => let);
   U2 : INV_X1 port map( A => eq_port, ZN => neq);
   U3 : NOR4_X1 port map( A1 => Sum(23), A2 => Sum(22), A3 => Sum(21), A4 => 
                           Sum(20), ZN => n9);
   U4 : NOR4_X1 port map( A1 => Sum(9), A2 => Sum(8), A3 => Sum(7), A4 => 
                           Sum(6), ZN => n13);
   U5 : NOR4_X1 port map( A1 => Sum(16), A2 => Sum(15), A3 => Sum(14), A4 => 
                           Sum(13), ZN => n7);
   U6 : NOR2_X1 port map( A1 => lt_port, A2 => eq_port, ZN => gt_port);
   U7 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => eq_port);
   U8 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => n4
                           );
   U9 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U10 : NOR4_X1 port map( A1 => Sum(27), A2 => Sum(26), A3 => Sum(25), A4 => 
                           Sum(24), ZN => n10);
   U11 : NOR4_X1 port map( A1 => Sum(1), A2 => Sum(19), A3 => Sum(18), A4 => 
                           Sum(17), ZN => n8);
   U12 : NOR4_X1 port map( A1 => Sum(5), A2 => Sum(4), A3 => Sum(3), A4 => 
                           Sum(31), ZN => n12);
   U13 : NOR4_X1 port map( A1 => Sum(30), A2 => Sum(2), A3 => Sum(29), A4 => 
                           Sum(28), ZN => n11);
   U14 : NOR4_X1 port map( A1 => Sum(12), A2 => Sum(11), A3 => Sum(10), A4 => 
                           Sum(0), ZN => n6);
   U15 : INV_X1 port map( A => get_port, ZN => lt_port);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity shifter is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (1 downto 0);  C : out std_logic_vector (31 downto 0));

end shifter;

architecture SYN_struct of shifter is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_thirdLevel
      port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector 
            (38 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_secondLevel
      port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : 
            in std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 
            downto 0));
   end component;
   
   component shift_firstLevel
      port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
            (1 downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 
            downto 0));
   end component;
   
   signal s3_2_port, s3_1_port, s3_0_port, m0_38_port, m0_37_port, m0_36_port, 
      m0_35_port, m0_34_port, m0_33_port, m0_32_port, m0_31_port, m0_30_port, 
      m0_29_port, m0_28_port, m0_27_port, m0_26_port, m0_25_port, m0_24_port, 
      m0_23_port, m0_22_port, m0_21_port, m0_20_port, m0_19_port, m0_18_port, 
      m0_17_port, m0_16_port, m0_15_port, m0_14_port, m0_13_port, m0_12_port, 
      m0_11_port, m0_10_port, m0_9_port, m0_8_port, m0_7_port, m0_6_port, 
      m0_5_port, m0_4_port, m0_3_port, m0_2_port, m0_1_port, m0_0_port, 
      m8_38_port, m8_37_port, m8_36_port, m8_35_port, m8_34_port, m8_33_port, 
      m8_32_port, m8_31_port, m8_30_port, m8_29_port, m8_28_port, m8_27_port, 
      m8_26_port, m8_25_port, m8_24_port, m8_23_port, m8_22_port, m8_21_port, 
      m8_20_port, m8_19_port, m8_18_port, m8_17_port, m8_16_port, m8_15_port, 
      m8_14_port, m8_13_port, m8_12_port, m8_11_port, m8_10_port, m8_9_port, 
      m8_8_port, m8_7_port, m8_6_port, m8_5_port, m8_4_port, m8_3_port, 
      m8_2_port, m8_1_port, m8_0_port, m16_38_port, m16_37_port, m16_36_port, 
      m16_35_port, m16_34_port, m16_33_port, m16_32_port, m16_31_port, 
      m16_30_port, m16_29_port, m16_28_port, m16_27_port, m16_26_port, 
      m16_25_port, m16_24_port, m16_23_port, m16_22_port, m16_21_port, 
      m16_20_port, m16_19_port, m16_18_port, m16_17_port, m16_16_port, 
      m16_15_port, m16_14_port, m16_13_port, m16_12_port, m16_11_port, 
      m16_10_port, m16_9_port, m16_8_port, m16_7_port, m16_6_port, m16_5_port, 
      m16_4_port, m16_3_port, m16_2_port, m16_1_port, m16_0_port, y_38_port, 
      y_37_port, y_36_port, y_35_port, y_34_port, y_33_port, y_32_port, 
      y_31_port, y_30_port, y_29_port, y_28_port, y_27_port, y_26_port, 
      y_25_port, y_24_port, y_23_port, y_22_port, y_21_port, y_20_port, 
      y_19_port, y_18_port, y_17_port, y_16_port, y_15_port, y_14_port, 
      y_13_port, y_12_port, y_11_port, y_10_port, y_9_port, y_8_port, y_7_port,
      y_6_port, y_5_port, y_4_port, y_3_port, y_2_port, y_1_port, y_0_port, n6,
      n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   IL : shift_firstLevel port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), sel(1) => sel(1), sel(0) => sel(0), 
                           mask00(38) => m0_38_port, mask00(37) => m0_37_port, 
                           mask00(36) => m0_36_port, mask00(35) => m0_35_port, 
                           mask00(34) => m0_34_port, mask00(33) => m0_33_port, 
                           mask00(32) => m0_32_port, mask00(31) => m0_31_port, 
                           mask00(30) => m0_30_port, mask00(29) => m0_29_port, 
                           mask00(28) => m0_28_port, mask00(27) => m0_27_port, 
                           mask00(26) => m0_26_port, mask00(25) => m0_25_port, 
                           mask00(24) => m0_24_port, mask00(23) => m0_23_port, 
                           mask00(22) => m0_22_port, mask00(21) => m0_21_port, 
                           mask00(20) => m0_20_port, mask00(19) => m0_19_port, 
                           mask00(18) => m0_18_port, mask00(17) => m0_17_port, 
                           mask00(16) => m0_16_port, mask00(15) => m0_15_port, 
                           mask00(14) => m0_14_port, mask00(13) => m0_13_port, 
                           mask00(12) => m0_12_port, mask00(11) => m0_11_port, 
                           mask00(10) => m0_10_port, mask00(9) => m0_9_port, 
                           mask00(8) => m0_8_port, mask00(7) => m0_7_port, 
                           mask00(6) => m0_6_port, mask00(5) => m0_5_port, 
                           mask00(4) => m0_4_port, mask00(3) => m0_3_port, 
                           mask00(2) => m0_2_port, mask00(1) => m0_1_port, 
                           mask00(0) => m0_0_port, mask08(38) => m8_38_port, 
                           mask08(37) => m8_37_port, mask08(36) => m8_36_port, 
                           mask08(35) => m8_35_port, mask08(34) => m8_34_port, 
                           mask08(33) => m8_33_port, mask08(32) => m8_32_port, 
                           mask08(31) => m8_31_port, mask08(30) => m8_30_port, 
                           mask08(29) => m8_29_port, mask08(28) => m8_28_port, 
                           mask08(27) => m8_27_port, mask08(26) => m8_26_port, 
                           mask08(25) => m8_25_port, mask08(24) => m8_24_port, 
                           mask08(23) => m8_23_port, mask08(22) => m8_22_port, 
                           mask08(21) => m8_21_port, mask08(20) => m8_20_port, 
                           mask08(19) => m8_19_port, mask08(18) => m8_18_port, 
                           mask08(17) => m8_17_port, mask08(16) => m8_16_port, 
                           mask08(15) => m8_15_port, mask08(14) => m8_14_port, 
                           mask08(13) => m8_13_port, mask08(12) => m8_12_port, 
                           mask08(11) => m8_11_port, mask08(10) => m8_10_port, 
                           mask08(9) => m8_9_port, mask08(8) => m8_8_port, 
                           mask08(7) => m8_7_port, mask08(6) => m8_6_port, 
                           mask08(5) => m8_5_port, mask08(4) => m8_4_port, 
                           mask08(3) => m8_3_port, mask08(2) => m8_2_port, 
                           mask08(1) => m8_1_port, mask08(0) => m8_0_port, 
                           mask16(38) => m16_38_port, mask16(37) => m16_37_port
                           , mask16(36) => m16_36_port, mask16(35) => 
                           m16_35_port, mask16(34) => m16_34_port, mask16(33) 
                           => m16_33_port, mask16(32) => m16_32_port, 
                           mask16(31) => m16_31_port, mask16(30) => m16_30_port
                           , mask16(29) => m16_29_port, mask16(28) => 
                           m16_28_port, mask16(27) => m16_27_port, mask16(26) 
                           => m16_26_port, mask16(25) => m16_25_port, 
                           mask16(24) => m16_24_port, mask16(23) => m16_23_port
                           , mask16(22) => m16_22_port, mask16(21) => 
                           m16_21_port, mask16(20) => m16_20_port, mask16(19) 
                           => m16_19_port, mask16(18) => m16_18_port, 
                           mask16(17) => m16_17_port, mask16(16) => m16_16_port
                           , mask16(15) => m16_15_port, mask16(14) => 
                           m16_14_port, mask16(13) => m16_13_port, mask16(12) 
                           => m16_12_port, mask16(11) => m16_11_port, 
                           mask16(10) => m16_10_port, mask16(9) => m16_9_port, 
                           mask16(8) => m16_8_port, mask16(7) => m16_7_port, 
                           mask16(6) => m16_6_port, mask16(5) => m16_5_port, 
                           mask16(4) => m16_4_port, mask16(3) => m16_3_port, 
                           mask16(2) => m16_2_port, mask16(1) => m16_1_port, 
                           mask16(0) => m16_0_port);
   IIL : shift_secondLevel port map( sel(1) => B(4), sel(0) => B(3), mask00(38)
                           => m0_38_port, mask00(37) => m0_37_port, mask00(36) 
                           => m0_36_port, mask00(35) => m0_35_port, mask00(34) 
                           => m0_34_port, mask00(33) => m0_33_port, mask00(32) 
                           => m0_32_port, mask00(31) => m0_31_port, mask00(30) 
                           => m0_30_port, mask00(29) => m0_29_port, mask00(28) 
                           => m0_28_port, mask00(27) => m0_27_port, mask00(26) 
                           => m0_26_port, mask00(25) => m0_25_port, mask00(24) 
                           => m0_24_port, mask00(23) => m0_23_port, mask00(22) 
                           => m0_22_port, mask00(21) => m0_21_port, mask00(20) 
                           => m0_20_port, mask00(19) => m0_19_port, mask00(18) 
                           => m0_18_port, mask00(17) => m0_17_port, mask00(16) 
                           => m0_16_port, mask00(15) => m0_15_port, mask00(14) 
                           => m0_14_port, mask00(13) => m0_13_port, mask00(12) 
                           => m0_12_port, mask00(11) => m0_11_port, mask00(10) 
                           => m0_10_port, mask00(9) => m0_9_port, mask00(8) => 
                           m0_8_port, mask00(7) => m0_7_port, mask00(6) => 
                           m0_6_port, mask00(5) => m0_5_port, mask00(4) => 
                           m0_4_port, mask00(3) => m0_3_port, mask00(2) => 
                           m0_2_port, mask00(1) => m0_1_port, mask00(0) => 
                           m0_0_port, mask08(38) => m8_38_port, mask08(37) => 
                           m8_37_port, mask08(36) => m8_36_port, mask08(35) => 
                           m8_35_port, mask08(34) => m8_34_port, mask08(33) => 
                           m8_33_port, mask08(32) => m8_32_port, mask08(31) => 
                           m8_31_port, mask08(30) => m8_30_port, mask08(29) => 
                           m8_29_port, mask08(28) => m8_28_port, mask08(27) => 
                           m8_27_port, mask08(26) => m8_26_port, mask08(25) => 
                           m8_25_port, mask08(24) => m8_24_port, mask08(23) => 
                           m8_23_port, mask08(22) => m8_22_port, mask08(21) => 
                           m8_21_port, mask08(20) => m8_20_port, mask08(19) => 
                           m8_19_port, mask08(18) => m8_18_port, mask08(17) => 
                           m8_17_port, mask08(16) => m8_16_port, mask08(15) => 
                           m8_15_port, mask08(14) => m8_14_port, mask08(13) => 
                           m8_13_port, mask08(12) => m8_12_port, mask08(11) => 
                           m8_11_port, mask08(10) => m8_10_port, mask08(9) => 
                           m8_9_port, mask08(8) => m8_8_port, mask08(7) => 
                           m8_7_port, mask08(6) => m8_6_port, mask08(5) => 
                           m8_5_port, mask08(4) => m8_4_port, mask08(3) => 
                           m8_3_port, mask08(2) => m8_2_port, mask08(1) => 
                           m8_1_port, mask08(0) => m8_0_port, mask16(38) => 
                           m16_38_port, mask16(37) => m16_37_port, mask16(36) 
                           => m16_36_port, mask16(35) => m16_35_port, 
                           mask16(34) => m16_34_port, mask16(33) => m16_33_port
                           , mask16(32) => m16_32_port, mask16(31) => 
                           m16_31_port, mask16(30) => m16_30_port, mask16(29) 
                           => m16_29_port, mask16(28) => m16_28_port, 
                           mask16(27) => m16_27_port, mask16(26) => m16_26_port
                           , mask16(25) => m16_25_port, mask16(24) => 
                           m16_24_port, mask16(23) => m16_23_port, mask16(22) 
                           => m16_22_port, mask16(21) => m16_21_port, 
                           mask16(20) => m16_20_port, mask16(19) => m16_19_port
                           , mask16(18) => m16_18_port, mask16(17) => 
                           m16_17_port, mask16(16) => m16_16_port, mask16(15) 
                           => m16_15_port, mask16(14) => m16_14_port, 
                           mask16(13) => m16_13_port, mask16(12) => m16_12_port
                           , mask16(11) => m16_11_port, mask16(10) => 
                           m16_10_port, mask16(9) => m16_9_port, mask16(8) => 
                           m16_8_port, mask16(7) => m16_7_port, mask16(6) => 
                           m16_6_port, mask16(5) => m16_5_port, mask16(4) => 
                           m16_4_port, mask16(3) => m16_3_port, mask16(2) => 
                           m16_2_port, mask16(1) => m16_1_port, mask16(0) => 
                           m16_0_port, Y(38) => y_38_port, Y(37) => y_37_port, 
                           Y(36) => y_36_port, Y(35) => y_35_port, Y(34) => 
                           y_34_port, Y(33) => y_33_port, Y(32) => y_32_port, 
                           Y(31) => y_31_port, Y(30) => y_30_port, Y(29) => 
                           y_29_port, Y(28) => y_28_port, Y(27) => y_27_port, 
                           Y(26) => y_26_port, Y(25) => y_25_port, Y(24) => 
                           y_24_port, Y(23) => y_23_port, Y(22) => y_22_port, 
                           Y(21) => y_21_port, Y(20) => y_20_port, Y(19) => 
                           y_19_port, Y(18) => y_18_port, Y(17) => y_17_port, 
                           Y(16) => y_16_port, Y(15) => y_15_port, Y(14) => 
                           y_14_port, Y(13) => y_13_port, Y(12) => y_12_port, 
                           Y(11) => y_11_port, Y(10) => y_10_port, Y(9) => 
                           y_9_port, Y(8) => y_8_port, Y(7) => y_7_port, Y(6) 
                           => y_6_port, Y(5) => y_5_port, Y(4) => y_4_port, 
                           Y(3) => y_3_port, Y(2) => y_2_port, Y(1) => y_1_port
                           , Y(0) => y_0_port);
   IIIL : shift_thirdLevel port map( sel(2) => s3_2_port, sel(1) => s3_1_port, 
                           sel(0) => s3_0_port, A(38) => y_38_port, A(37) => 
                           y_37_port, A(36) => y_36_port, A(35) => y_35_port, 
                           A(34) => y_34_port, A(33) => y_33_port, A(32) => 
                           y_32_port, A(31) => y_31_port, A(30) => y_30_port, 
                           A(29) => y_29_port, A(28) => y_28_port, A(27) => 
                           y_27_port, A(26) => y_26_port, A(25) => y_25_port, 
                           A(24) => y_24_port, A(23) => y_23_port, A(22) => 
                           y_22_port, A(21) => y_21_port, A(20) => y_20_port, 
                           A(19) => y_19_port, A(18) => y_18_port, A(17) => 
                           y_17_port, A(16) => y_16_port, A(15) => y_15_port, 
                           A(14) => y_14_port, A(13) => y_13_port, A(12) => 
                           y_12_port, A(11) => y_11_port, A(10) => y_10_port, 
                           A(9) => y_9_port, A(8) => y_8_port, A(7) => y_7_port
                           , A(6) => y_6_port, A(5) => y_5_port, A(4) => 
                           y_4_port, A(3) => y_3_port, A(2) => y_2_port, A(1) 
                           => y_1_port, A(0) => y_0_port, Y(31) => C(31), Y(30)
                           => C(30), Y(29) => C(29), Y(28) => C(28), Y(27) => 
                           C(27), Y(26) => C(26), Y(25) => C(25), Y(24) => 
                           C(24), Y(23) => C(23), Y(22) => C(22), Y(21) => 
                           C(21), Y(20) => C(20), Y(19) => C(19), Y(18) => 
                           C(18), Y(17) => C(17), Y(16) => C(16), Y(15) => 
                           C(15), Y(14) => C(14), Y(13) => C(13), Y(12) => 
                           C(12), Y(11) => C(11), Y(10) => C(10), Y(9) => C(9),
                           Y(8) => C(8), Y(7) => C(7), Y(6) => C(6), Y(5) => 
                           C(5), Y(4) => C(4), Y(3) => C(3), Y(2) => C(2), Y(1)
                           => C(1), Y(0) => C(0));
   U1 : AOI221_X1 port map( B1 => n6, B2 => n7, C1 => sel(0), C2 => B(2), A => 
                           n8, ZN => s3_2_port);
   U2 : INV_X1 port map( A => n6, ZN => n11);
   U3 : INV_X1 port map( A => B(2), ZN => n7);
   U4 : INV_X1 port map( A => n9, ZN => n8);
   U5 : OAI21_X1 port map( B1 => B(2), B2 => sel(0), A => sel(1), ZN => n9);
   U6 : OAI22_X1 port map( A1 => B(0), A2 => n10, B1 => n11, B2 => n13, ZN => 
                           s3_0_port);
   U7 : INV_X1 port map( A => B(0), ZN => n13);
   U8 : OAI22_X1 port map( A1 => B(1), A2 => n10, B1 => n11, B2 => n12, ZN => 
                           s3_1_port);
   U9 : INV_X1 port map( A => B(1), ZN => n12);
   U10 : XNOR2_X1 port map( A => sel(1), B => sel(0), ZN => n10);
   U11 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n6);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity logical is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (3 downto 0);  Y : out std_logic_vector (31 downto 0));

end logical;

architecture SYN_behav of logical is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201 : 
      std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n121, A2 => n122, B1 => B(25), B2 => n123, ZN 
                           => Y(25));
   U2 : OAI22_X1 port map( A1 => n125, A2 => n126, B1 => B(24), B2 => n127, ZN 
                           => Y(24));
   U3 : OAI22_X1 port map( A1 => n129, A2 => n130, B1 => B(23), B2 => n131, ZN 
                           => Y(23));
   U4 : OAI22_X1 port map( A1 => n133, A2 => n134, B1 => B(22), B2 => n135, ZN 
                           => Y(22));
   U5 : OAI22_X1 port map( A1 => n137, A2 => n138, B1 => B(21), B2 => n139, ZN 
                           => Y(21));
   U6 : OAI22_X1 port map( A1 => n141, A2 => n142, B1 => B(20), B2 => n143, ZN 
                           => Y(20));
   U7 : OAI22_X1 port map( A1 => n149, A2 => n150, B1 => B(19), B2 => n151, ZN 
                           => Y(19));
   U8 : OAI22_X1 port map( A1 => n153, A2 => n154, B1 => B(18), B2 => n155, ZN 
                           => Y(18));
   U9 : OAI22_X1 port map( A1 => n157, A2 => n158, B1 => B(17), B2 => n159, ZN 
                           => Y(17));
   U10 : OAI22_X1 port map( A1 => n161, A2 => n162, B1 => B(16), B2 => n163, ZN
                           => Y(16));
   U11 : OAI22_X1 port map( A1 => n165, A2 => n166, B1 => B(15), B2 => n167, ZN
                           => Y(15));
   U12 : OAI22_X1 port map( A1 => n169, A2 => n170, B1 => B(14), B2 => n171, ZN
                           => Y(14));
   U13 : OAI22_X1 port map( A1 => n173, A2 => n174, B1 => B(13), B2 => n175, ZN
                           => Y(13));
   U14 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => B(7), B2 => n75, ZN => 
                           Y(7));
   U15 : OAI22_X1 port map( A1 => n77, A2 => n78, B1 => B(6), B2 => n79, ZN => 
                           Y(6));
   U16 : OAI22_X1 port map( A1 => n81, A2 => n82, B1 => B(5), B2 => n83, ZN => 
                           Y(5));
   U17 : OAI22_X1 port map( A1 => n85, A2 => n86, B1 => B(4), B2 => n87, ZN => 
                           Y(4));
   U18 : OAI22_X1 port map( A1 => n89, A2 => n90, B1 => B(3), B2 => n91, ZN => 
                           Y(3));
   U19 : OAI22_X1 port map( A1 => n101, A2 => n102, B1 => B(2), B2 => n103, ZN 
                           => Y(2));
   U20 : OAI22_X1 port map( A1 => n145, A2 => n146, B1 => B(1), B2 => n147, ZN 
                           => Y(1));
   U21 : OAI22_X1 port map( A1 => n93, A2 => n94, B1 => B(31), B2 => n95, ZN =>
                           Y(31));
   U22 : OAI22_X1 port map( A1 => n97, A2 => n98, B1 => B(30), B2 => n99, ZN =>
                           Y(30));
   U23 : OAI22_X1 port map( A1 => n105, A2 => n106, B1 => B(29), B2 => n107, ZN
                           => Y(29));
   U24 : OAI22_X1 port map( A1 => n109, A2 => n110, B1 => B(28), B2 => n111, ZN
                           => Y(28));
   U25 : OAI22_X1 port map( A1 => n113, A2 => n114, B1 => B(27), B2 => n115, ZN
                           => Y(27));
   U26 : OAI22_X1 port map( A1 => n117, A2 => n118, B1 => B(26), B2 => n119, ZN
                           => Y(26));
   U27 : OAI22_X1 port map( A1 => n177, A2 => n178, B1 => B(12), B2 => n179, ZN
                           => Y(12));
   U28 : OAI22_X1 port map( A1 => n181, A2 => n182, B1 => B(11), B2 => n183, ZN
                           => Y(11));
   U29 : OAI22_X1 port map( A1 => n185, A2 => n186, B1 => B(10), B2 => n187, ZN
                           => Y(10));
   U30 : OAI22_X1 port map( A1 => n65, A2 => n66, B1 => B(9), B2 => n67, ZN => 
                           Y(9));
   U31 : OAI22_X1 port map( A1 => n69, A2 => n70, B1 => B(8), B2 => n71, ZN => 
                           Y(8));
   U32 : BUF_X1 port map( A => sel(1), Z => n197);
   U33 : BUF_X1 port map( A => sel(0), Z => n194);
   U34 : BUF_X1 port map( A => sel(1), Z => n196);
   U35 : BUF_X1 port map( A => sel(0), Z => n193);
   U36 : OAI22_X1 port map( A1 => n189, A2 => n190, B1 => B(0), B2 => n191, ZN 
                           => Y(0));
   U37 : INV_X1 port map( A => B(0), ZN => n190);
   U38 : AOI22_X1 port map( A1 => n199, A2 => n192, B1 => A(0), B2 => n193, ZN 
                           => n189);
   U39 : AOI22_X1 port map( A1 => sel(3), A2 => n192, B1 => A(0), B2 => n196, 
                           ZN => n191);
   U40 : BUF_X1 port map( A => sel(2), Z => n200);
   U41 : BUF_X1 port map( A => sel(2), Z => n199);
   U42 : BUF_X1 port map( A => sel(1), Z => n198);
   U43 : BUF_X1 port map( A => sel(0), Z => n195);
   U44 : BUF_X1 port map( A => sel(2), Z => n201);
   U45 : AOI22_X1 port map( A1 => sel(3), A2 => n96, B1 => A(31), B2 => n198, 
                           ZN => n95);
   U46 : AOI22_X1 port map( A1 => sel(3), A2 => n72, B1 => A(8), B2 => n198, ZN
                           => n71);
   U47 : AOI22_X1 port map( A1 => sel(3), A2 => n76, B1 => A(7), B2 => n198, ZN
                           => n75);
   U48 : AOI22_X1 port map( A1 => sel(3), A2 => n80, B1 => A(6), B2 => n198, ZN
                           => n79);
   U49 : AOI22_X1 port map( A1 => sel(3), A2 => n84, B1 => A(5), B2 => n198, ZN
                           => n83);
   U50 : AOI22_X1 port map( A1 => sel(3), A2 => n88, B1 => A(4), B2 => n198, ZN
                           => n87);
   U51 : AOI22_X1 port map( A1 => sel(3), A2 => n92, B1 => A(3), B2 => n198, ZN
                           => n91);
   U52 : AOI22_X1 port map( A1 => sel(3), A2 => n68, B1 => n198, B2 => A(9), ZN
                           => n67);
   U53 : AOI22_X1 port map( A1 => sel(3), A2 => n100, B1 => A(30), B2 => n197, 
                           ZN => n99);
   U54 : AOI22_X1 port map( A1 => sel(3), A2 => n108, B1 => A(29), B2 => n197, 
                           ZN => n107);
   U55 : AOI22_X1 port map( A1 => sel(3), A2 => n112, B1 => A(28), B2 => n197, 
                           ZN => n111);
   U56 : AOI22_X1 port map( A1 => sel(3), A2 => n116, B1 => A(27), B2 => n197, 
                           ZN => n115);
   U57 : AOI22_X1 port map( A1 => sel(3), A2 => n120, B1 => A(26), B2 => n197, 
                           ZN => n119);
   U58 : AOI22_X1 port map( A1 => sel(3), A2 => n124, B1 => A(25), B2 => n197, 
                           ZN => n123);
   U59 : AOI22_X1 port map( A1 => sel(3), A2 => n128, B1 => A(24), B2 => n197, 
                           ZN => n127);
   U60 : AOI22_X1 port map( A1 => sel(3), A2 => n132, B1 => A(23), B2 => n197, 
                           ZN => n131);
   U61 : AOI22_X1 port map( A1 => sel(3), A2 => n136, B1 => A(22), B2 => n197, 
                           ZN => n135);
   U62 : AOI22_X1 port map( A1 => sel(3), A2 => n140, B1 => A(21), B2 => n197, 
                           ZN => n139);
   U63 : AOI22_X1 port map( A1 => sel(3), A2 => n144, B1 => A(20), B2 => n197, 
                           ZN => n143);
   U64 : AOI22_X1 port map( A1 => sel(3), A2 => n152, B1 => A(19), B2 => n196, 
                           ZN => n151);
   U65 : AOI22_X1 port map( A1 => sel(3), A2 => n156, B1 => A(18), B2 => n196, 
                           ZN => n155);
   U66 : AOI22_X1 port map( A1 => sel(3), A2 => n160, B1 => A(17), B2 => n196, 
                           ZN => n159);
   U67 : AOI22_X1 port map( A1 => sel(3), A2 => n164, B1 => A(16), B2 => n196, 
                           ZN => n163);
   U68 : AOI22_X1 port map( A1 => sel(3), A2 => n168, B1 => A(15), B2 => n196, 
                           ZN => n167);
   U69 : AOI22_X1 port map( A1 => sel(3), A2 => n172, B1 => A(14), B2 => n196, 
                           ZN => n171);
   U70 : AOI22_X1 port map( A1 => sel(3), A2 => n176, B1 => A(13), B2 => n196, 
                           ZN => n175);
   U71 : AOI22_X1 port map( A1 => sel(3), A2 => n180, B1 => A(12), B2 => n196, 
                           ZN => n179);
   U72 : AOI22_X1 port map( A1 => sel(3), A2 => n184, B1 => A(11), B2 => n196, 
                           ZN => n183);
   U73 : AOI22_X1 port map( A1 => sel(3), A2 => n188, B1 => A(10), B2 => n196, 
                           ZN => n187);
   U74 : AOI22_X1 port map( A1 => sel(3), A2 => n104, B1 => A(2), B2 => n197, 
                           ZN => n103);
   U75 : AOI22_X1 port map( A1 => sel(3), A2 => n148, B1 => A(1), B2 => n196, 
                           ZN => n147);
   U76 : AOI22_X1 port map( A1 => n201, A2 => n96, B1 => A(31), B2 => n195, ZN 
                           => n93);
   U77 : AOI22_X1 port map( A1 => n201, A2 => n72, B1 => A(8), B2 => n195, ZN 
                           => n69);
   U78 : AOI22_X1 port map( A1 => n201, A2 => n76, B1 => A(7), B2 => n195, ZN 
                           => n73);
   U79 : AOI22_X1 port map( A1 => n201, A2 => n80, B1 => A(6), B2 => n195, ZN 
                           => n77);
   U80 : AOI22_X1 port map( A1 => n201, A2 => n84, B1 => A(5), B2 => n195, ZN 
                           => n81);
   U81 : AOI22_X1 port map( A1 => n201, A2 => n88, B1 => A(4), B2 => n195, ZN 
                           => n85);
   U82 : AOI22_X1 port map( A1 => n201, A2 => n92, B1 => A(3), B2 => n195, ZN 
                           => n89);
   U83 : AOI22_X1 port map( A1 => n201, A2 => n68, B1 => n195, B2 => A(9), ZN 
                           => n65);
   U84 : AOI22_X1 port map( A1 => n200, A2 => n100, B1 => A(30), B2 => n194, ZN
                           => n97);
   U85 : AOI22_X1 port map( A1 => n200, A2 => n108, B1 => A(29), B2 => n194, ZN
                           => n105);
   U86 : AOI22_X1 port map( A1 => n200, A2 => n112, B1 => A(28), B2 => n194, ZN
                           => n109);
   U87 : AOI22_X1 port map( A1 => n200, A2 => n116, B1 => A(27), B2 => n194, ZN
                           => n113);
   U88 : AOI22_X1 port map( A1 => n200, A2 => n120, B1 => A(26), B2 => n194, ZN
                           => n117);
   U89 : AOI22_X1 port map( A1 => n200, A2 => n124, B1 => A(25), B2 => n194, ZN
                           => n121);
   U90 : AOI22_X1 port map( A1 => n200, A2 => n128, B1 => A(24), B2 => n194, ZN
                           => n125);
   U91 : AOI22_X1 port map( A1 => n200, A2 => n132, B1 => A(23), B2 => n194, ZN
                           => n129);
   U92 : AOI22_X1 port map( A1 => n200, A2 => n136, B1 => A(22), B2 => n194, ZN
                           => n133);
   U93 : AOI22_X1 port map( A1 => n200, A2 => n140, B1 => A(21), B2 => n194, ZN
                           => n137);
   U94 : AOI22_X1 port map( A1 => n200, A2 => n144, B1 => A(20), B2 => n194, ZN
                           => n141);
   U95 : AOI22_X1 port map( A1 => n199, A2 => n152, B1 => A(19), B2 => n193, ZN
                           => n149);
   U96 : AOI22_X1 port map( A1 => n199, A2 => n156, B1 => A(18), B2 => n193, ZN
                           => n153);
   U97 : AOI22_X1 port map( A1 => n199, A2 => n160, B1 => A(17), B2 => n193, ZN
                           => n157);
   U98 : AOI22_X1 port map( A1 => n199, A2 => n164, B1 => A(16), B2 => n193, ZN
                           => n161);
   U99 : AOI22_X1 port map( A1 => n199, A2 => n168, B1 => A(15), B2 => n193, ZN
                           => n165);
   U100 : AOI22_X1 port map( A1 => n199, A2 => n172, B1 => A(14), B2 => n193, 
                           ZN => n169);
   U101 : AOI22_X1 port map( A1 => n199, A2 => n176, B1 => A(13), B2 => n193, 
                           ZN => n173);
   U102 : AOI22_X1 port map( A1 => n199, A2 => n180, B1 => A(12), B2 => n193, 
                           ZN => n177);
   U103 : AOI22_X1 port map( A1 => n199, A2 => n184, B1 => A(11), B2 => n193, 
                           ZN => n181);
   U104 : AOI22_X1 port map( A1 => n199, A2 => n188, B1 => A(10), B2 => n193, 
                           ZN => n185);
   U105 : AOI22_X1 port map( A1 => n200, A2 => n104, B1 => A(2), B2 => n194, ZN
                           => n101);
   U106 : AOI22_X1 port map( A1 => n199, A2 => n148, B1 => A(1), B2 => n193, ZN
                           => n145);
   U107 : INV_X1 port map( A => A(9), ZN => n68);
   U108 : INV_X1 port map( A => A(31), ZN => n96);
   U109 : INV_X1 port map( A => A(30), ZN => n100);
   U110 : INV_X1 port map( A => A(29), ZN => n108);
   U111 : INV_X1 port map( A => A(28), ZN => n112);
   U112 : INV_X1 port map( A => A(27), ZN => n116);
   U113 : INV_X1 port map( A => A(26), ZN => n120);
   U114 : INV_X1 port map( A => A(25), ZN => n124);
   U115 : INV_X1 port map( A => A(24), ZN => n128);
   U116 : INV_X1 port map( A => A(23), ZN => n132);
   U117 : INV_X1 port map( A => A(22), ZN => n136);
   U118 : INV_X1 port map( A => A(21), ZN => n140);
   U119 : INV_X1 port map( A => A(20), ZN => n144);
   U120 : INV_X1 port map( A => A(19), ZN => n152);
   U121 : INV_X1 port map( A => A(18), ZN => n156);
   U122 : INV_X1 port map( A => A(17), ZN => n160);
   U123 : INV_X1 port map( A => A(16), ZN => n164);
   U124 : INV_X1 port map( A => A(15), ZN => n168);
   U125 : INV_X1 port map( A => A(14), ZN => n172);
   U126 : INV_X1 port map( A => A(13), ZN => n176);
   U127 : INV_X1 port map( A => A(12), ZN => n180);
   U128 : INV_X1 port map( A => A(11), ZN => n184);
   U129 : INV_X1 port map( A => A(10), ZN => n188);
   U130 : INV_X1 port map( A => A(8), ZN => n72);
   U131 : INV_X1 port map( A => A(7), ZN => n76);
   U132 : INV_X1 port map( A => A(6), ZN => n80);
   U133 : INV_X1 port map( A => A(5), ZN => n84);
   U134 : INV_X1 port map( A => A(4), ZN => n88);
   U135 : INV_X1 port map( A => A(3), ZN => n92);
   U136 : INV_X1 port map( A => A(2), ZN => n104);
   U137 : INV_X1 port map( A => A(1), ZN => n148);
   U138 : INV_X1 port map( A => A(0), ZN => n192);
   U139 : INV_X1 port map( A => B(31), ZN => n94);
   U140 : INV_X1 port map( A => B(30), ZN => n98);
   U141 : INV_X1 port map( A => B(29), ZN => n106);
   U142 : INV_X1 port map( A => B(28), ZN => n110);
   U143 : INV_X1 port map( A => B(27), ZN => n114);
   U144 : INV_X1 port map( A => B(26), ZN => n118);
   U145 : INV_X1 port map( A => B(25), ZN => n122);
   U146 : INV_X1 port map( A => B(24), ZN => n126);
   U147 : INV_X1 port map( A => B(23), ZN => n130);
   U148 : INV_X1 port map( A => B(22), ZN => n134);
   U149 : INV_X1 port map( A => B(21), ZN => n138);
   U150 : INV_X1 port map( A => B(20), ZN => n142);
   U151 : INV_X1 port map( A => B(19), ZN => n150);
   U152 : INV_X1 port map( A => B(18), ZN => n154);
   U153 : INV_X1 port map( A => B(17), ZN => n158);
   U154 : INV_X1 port map( A => B(16), ZN => n162);
   U155 : INV_X1 port map( A => B(15), ZN => n166);
   U156 : INV_X1 port map( A => B(14), ZN => n170);
   U157 : INV_X1 port map( A => B(13), ZN => n174);
   U158 : INV_X1 port map( A => B(12), ZN => n178);
   U159 : INV_X1 port map( A => B(11), ZN => n182);
   U160 : INV_X1 port map( A => B(10), ZN => n186);
   U161 : INV_X1 port map( A => B(9), ZN => n66);
   U162 : INV_X1 port map( A => B(8), ZN => n70);
   U163 : INV_X1 port map( A => B(7), ZN => n74);
   U164 : INV_X1 port map( A => B(6), ZN => n78);
   U165 : INV_X1 port map( A => B(5), ZN => n82);
   U166 : INV_X1 port map( A => B(4), ZN => n86);
   U167 : INV_X1 port map( A => B(3), ZN => n90);
   U168 : INV_X1 port map( A => B(2), ZN => n102);
   U169 : INV_X1 port map( A => B(1), ZN => n146);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity booth_mul_N16 is

   port( A, B : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end booth_mul_N16;

architecture SYN_struct of booth_mul_N16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component cla_adder_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_4
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_5
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CSA_Nbits32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  S, Cout : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux_N32_1
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_2
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_3
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_4
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_5
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_6
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_7
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_N32_0
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component shift_mul_N16_S14
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S12
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S10
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S8
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S6
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S4
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S2
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component shift_mul_N16_S0
      port( A : in std_logic_vector (15 downto 0);  B, C, D, E : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, muxInE_7_31_port, muxInE_7_30_port, muxInE_7_29_port, 
      muxInE_7_28_port, muxInE_7_27_port, muxInE_7_26_port, muxInE_7_25_port, 
      muxInE_7_24_port, muxInE_7_23_port, muxInE_7_22_port, muxInE_7_21_port, 
      muxInE_7_20_port, muxInE_7_19_port, muxInE_7_18_port, muxInE_7_17_port, 
      muxInE_7_16_port, muxInE_7_15_port, muxInE_7_14_port, muxInE_7_13_port, 
      muxInE_7_12_port, muxInE_7_11_port, muxInE_7_10_port, muxInE_7_9_port, 
      muxInE_7_8_port, muxInE_7_7_port, muxInE_7_6_port, muxInE_7_5_port, 
      muxInE_7_4_port, muxInE_7_3_port, muxInE_7_2_port, muxInE_7_1_port, 
      muxInE_7_0_port, muxInE_6_31_port, muxInE_6_30_port, muxInE_6_29_port, 
      muxInE_6_28_port, muxInE_6_27_port, muxInE_6_26_port, muxInE_6_25_port, 
      muxInE_6_24_port, muxInE_6_23_port, muxInE_6_22_port, muxInE_6_21_port, 
      muxInE_6_20_port, muxInE_6_19_port, muxInE_6_18_port, muxInE_6_17_port, 
      muxInE_6_16_port, muxInE_6_15_port, muxInE_6_14_port, muxInE_6_13_port, 
      muxInE_6_12_port, muxInE_6_11_port, muxInE_6_10_port, muxInE_6_9_port, 
      muxInE_6_8_port, muxInE_6_7_port, muxInE_6_6_port, muxInE_6_5_port, 
      muxInE_6_4_port, muxInE_6_3_port, muxInE_6_2_port, muxInE_6_1_port, 
      muxInE_6_0_port, muxInE_5_31_port, muxInE_5_30_port, muxInE_5_29_port, 
      muxInE_5_28_port, muxInE_5_27_port, muxInE_5_26_port, muxInE_5_25_port, 
      muxInE_5_24_port, muxInE_5_23_port, muxInE_5_22_port, muxInE_5_21_port, 
      muxInE_5_20_port, muxInE_5_19_port, muxInE_5_18_port, muxInE_5_17_port, 
      muxInE_5_16_port, muxInE_5_15_port, muxInE_5_14_port, muxInE_5_13_port, 
      muxInE_5_12_port, muxInE_5_11_port, muxInE_5_10_port, muxInE_5_9_port, 
      muxInE_5_8_port, muxInE_5_7_port, muxInE_5_6_port, muxInE_5_5_port, 
      muxInE_5_4_port, muxInE_5_3_port, muxInE_5_2_port, muxInE_5_1_port, 
      muxInE_5_0_port, muxInE_4_31_port, muxInE_4_30_port, muxInE_4_29_port, 
      muxInE_4_28_port, muxInE_4_27_port, muxInE_4_26_port, muxInE_4_25_port, 
      muxInE_4_24_port, muxInE_4_23_port, muxInE_4_22_port, muxInE_4_21_port, 
      muxInE_4_20_port, muxInE_4_19_port, muxInE_4_18_port, muxInE_4_17_port, 
      muxInE_4_16_port, muxInE_4_15_port, muxInE_4_14_port, muxInE_4_13_port, 
      muxInE_4_12_port, muxInE_4_11_port, muxInE_4_10_port, muxInE_4_9_port, 
      muxInE_4_8_port, muxInE_4_7_port, muxInE_4_6_port, muxInE_4_5_port, 
      muxInE_4_4_port, muxInE_4_3_port, muxInE_4_2_port, muxInE_4_1_port, 
      muxInE_4_0_port, muxInE_3_31_port, muxInE_3_30_port, muxInE_3_29_port, 
      muxInE_3_28_port, muxInE_3_27_port, muxInE_3_26_port, muxInE_3_25_port, 
      muxInE_3_24_port, muxInE_3_23_port, muxInE_3_22_port, muxInE_3_21_port, 
      muxInE_3_20_port, muxInE_3_19_port, muxInE_3_18_port, muxInE_3_17_port, 
      muxInE_3_16_port, muxInE_3_15_port, muxInE_3_14_port, muxInE_3_13_port, 
      muxInE_3_12_port, muxInE_3_11_port, muxInE_3_10_port, muxInE_3_9_port, 
      muxInE_3_8_port, muxInE_3_7_port, muxInE_3_6_port, muxInE_3_5_port, 
      muxInE_3_4_port, muxInE_3_3_port, muxInE_3_2_port, muxInE_3_1_port, 
      muxInE_3_0_port, muxInE_2_31_port, muxInE_2_30_port, muxInE_2_29_port, 
      muxInE_2_28_port, muxInE_2_27_port, muxInE_2_26_port, muxInE_2_25_port, 
      muxInE_2_24_port, muxInE_2_23_port, muxInE_2_22_port, muxInE_2_21_port, 
      muxInE_2_19_port, muxInE_2_18_port, muxInE_2_17_port, muxInE_2_16_port, 
      muxInE_2_15_port, muxInE_2_14_port, muxInE_2_13_port, muxInE_2_12_port, 
      muxInE_2_11_port, muxInE_2_10_port, muxInE_2_9_port, muxInE_2_8_port, 
      muxInE_2_7_port, muxInE_2_6_port, muxInE_2_5_port, muxInE_2_4_port, 
      muxInE_2_3_port, muxInE_2_2_port, muxInE_2_1_port, muxInE_2_0_port, 
      muxInE_1_31_port, muxInE_1_30_port, muxInE_1_29_port, muxInE_1_28_port, 
      muxInE_1_27_port, muxInE_1_26_port, muxInE_1_25_port, muxInE_1_24_port, 
      muxInE_1_23_port, muxInE_1_22_port, muxInE_1_21_port, muxInE_1_20_port, 
      muxInE_1_19_port, muxInE_1_18_port, muxInE_1_17_port, muxInE_1_16_port, 
      muxInE_1_15_port, muxInE_1_14_port, muxInE_1_13_port, muxInE_1_12_port, 
      muxInE_1_11_port, muxInE_1_10_port, muxInE_1_9_port, muxInE_1_8_port, 
      muxInE_1_7_port, muxInE_1_6_port, muxInE_1_5_port, muxInE_1_4_port, 
      muxInE_1_3_port, muxInE_1_2_port, muxInE_1_1_port, muxInE_1_0_port, 
      muxInE_0_31_port, muxInE_0_30_port, muxInE_0_29_port, muxInE_0_28_port, 
      muxInE_0_27_port, muxInE_0_26_port, muxInE_0_24_port, muxInE_0_23_port, 
      muxInE_0_21_port, muxInE_0_20_port, muxInE_0_19_port, muxInE_0_18_port, 
      muxInE_0_16_port, muxInE_0_15_port, muxInE_0_14_port, muxInE_0_13_port, 
      muxInE_0_12_port, muxInE_0_11_port, muxInE_0_10_port, muxInE_0_9_port, 
      muxInE_0_8_port, muxInE_0_7_port, muxInE_0_6_port, muxInE_0_5_port, 
      muxInE_0_4_port, muxInE_0_3_port, muxInE_0_2_port, muxInE_0_1_port, 
      muxInE_0_0_port, muxInD_7_31_port, muxInD_7_30_port, muxInD_7_29_port, 
      muxInD_7_28_port, muxInD_7_27_port, muxInD_7_26_port, muxInD_7_25_port, 
      muxInD_7_24_port, muxInD_7_23_port, muxInD_7_22_port, muxInD_7_21_port, 
      muxInD_7_20_port, muxInD_7_19_port, muxInD_7_18_port, muxInD_7_17_port, 
      muxInD_7_16_port, muxInD_7_15_port, muxInD_7_14_port, muxInD_7_13_port, 
      muxInD_7_12_port, muxInD_7_11_port, muxInD_7_10_port, muxInD_7_9_port, 
      muxInD_7_8_port, muxInD_7_7_port, muxInD_7_6_port, muxInD_7_5_port, 
      muxInD_7_4_port, muxInD_7_3_port, muxInD_7_2_port, muxInD_7_1_port, 
      muxInD_7_0_port, muxInD_6_31_port, muxInD_6_30_port, muxInD_6_29_port, 
      muxInD_6_28_port, muxInD_6_27_port, muxInD_6_26_port, muxInD_6_25_port, 
      muxInD_6_24_port, muxInD_6_23_port, muxInD_6_22_port, muxInD_6_21_port, 
      muxInD_6_20_port, muxInD_6_19_port, muxInD_6_18_port, muxInD_6_17_port, 
      muxInD_6_16_port, muxInD_6_15_port, muxInD_6_14_port, muxInD_6_13_port, 
      muxInD_6_12_port, muxInD_6_11_port, muxInD_6_10_port, muxInD_6_9_port, 
      muxInD_6_8_port, muxInD_6_7_port, muxInD_6_6_port, muxInD_6_5_port, 
      muxInD_6_4_port, muxInD_6_3_port, muxInD_6_2_port, muxInD_6_1_port, 
      muxInD_6_0_port, muxInD_5_31_port, muxInD_5_30_port, muxInD_5_29_port, 
      muxInD_5_28_port, muxInD_5_27_port, muxInD_5_26_port, muxInD_5_25_port, 
      muxInD_5_24_port, muxInD_5_23_port, muxInD_5_22_port, muxInD_5_21_port, 
      muxInD_5_20_port, muxInD_5_19_port, muxInD_5_18_port, muxInD_5_17_port, 
      muxInD_5_16_port, muxInD_5_15_port, muxInD_5_14_port, muxInD_5_13_port, 
      muxInD_5_12_port, muxInD_5_11_port, muxInD_5_10_port, muxInD_5_9_port, 
      muxInD_5_8_port, muxInD_5_7_port, muxInD_5_6_port, muxInD_5_5_port, 
      muxInD_5_4_port, muxInD_5_3_port, muxInD_5_2_port, muxInD_5_1_port, 
      muxInD_5_0_port, muxInD_4_31_port, muxInD_4_30_port, muxInD_4_29_port, 
      muxInD_4_28_port, muxInD_4_27_port, muxInD_4_26_port, muxInD_4_25_port, 
      muxInD_4_24_port, muxInD_4_23_port, muxInD_4_22_port, muxInD_4_21_port, 
      muxInD_4_20_port, muxInD_4_19_port, muxInD_4_18_port, muxInD_4_17_port, 
      muxInD_4_16_port, muxInD_4_15_port, muxInD_4_14_port, muxInD_4_13_port, 
      muxInD_4_12_port, muxInD_4_11_port, muxInD_4_10_port, muxInD_4_9_port, 
      muxInD_4_8_port, muxInD_4_7_port, muxInD_4_6_port, muxInD_4_5_port, 
      muxInD_4_4_port, muxInD_4_3_port, muxInD_4_2_port, muxInD_4_1_port, 
      muxInD_4_0_port, muxInD_3_31_port, muxInD_3_30_port, muxInD_3_29_port, 
      muxInD_3_28_port, muxInD_3_27_port, muxInD_3_26_port, muxInD_3_25_port, 
      muxInD_3_24_port, muxInD_3_23_port, muxInD_3_22_port, muxInD_3_21_port, 
      muxInD_3_20_port, muxInD_3_19_port, muxInD_3_18_port, muxInD_3_17_port, 
      muxInD_3_16_port, muxInD_3_15_port, muxInD_3_14_port, muxInD_3_13_port, 
      muxInD_3_12_port, muxInD_3_11_port, muxInD_3_10_port, muxInD_3_9_port, 
      muxInD_3_8_port, muxInD_3_7_port, muxInD_3_6_port, muxInD_3_5_port, 
      muxInD_3_4_port, muxInD_3_3_port, muxInD_3_2_port, muxInD_3_1_port, 
      muxInD_3_0_port, muxInD_2_31_port, muxInD_2_30_port, muxInD_2_29_port, 
      muxInD_2_28_port, muxInD_2_27_port, muxInD_2_26_port, muxInD_2_25_port, 
      muxInD_2_24_port, muxInD_2_23_port, muxInD_2_22_port, muxInD_2_21_port, 
      muxInD_2_20_port, muxInD_2_19_port, muxInD_2_18_port, muxInD_2_17_port, 
      muxInD_2_16_port, muxInD_2_15_port, muxInD_2_14_port, muxInD_2_13_port, 
      muxInD_2_12_port, muxInD_2_11_port, muxInD_2_10_port, muxInD_2_9_port, 
      muxInD_2_8_port, muxInD_2_7_port, muxInD_2_6_port, muxInD_2_5_port, 
      muxInD_2_4_port, muxInD_2_3_port, muxInD_2_2_port, muxInD_2_1_port, 
      muxInD_2_0_port, muxInD_1_31_port, muxInD_1_30_port, muxInD_1_29_port, 
      muxInD_1_28_port, muxInD_1_27_port, muxInD_1_26_port, muxInD_1_25_port, 
      muxInD_1_24_port, muxInD_1_23_port, muxInD_1_22_port, muxInD_1_21_port, 
      muxInD_1_20_port, muxInD_1_19_port, muxInD_1_18_port, muxInD_1_17_port, 
      muxInD_1_16_port, muxInD_1_15_port, muxInD_1_14_port, muxInD_1_13_port, 
      muxInD_1_12_port, muxInD_1_11_port, muxInD_1_10_port, muxInD_1_9_port, 
      muxInD_1_8_port, muxInD_1_7_port, muxInD_1_6_port, muxInD_1_5_port, 
      muxInD_1_4_port, muxInD_1_3_port, muxInD_1_2_port, muxInD_1_1_port, 
      muxInD_1_0_port, muxInD_0_31_port, muxInD_0_30_port, muxInD_0_29_port, 
      muxInD_0_28_port, muxInD_0_27_port, muxInD_0_26_port, muxInD_0_25_port, 
      muxInD_0_24_port, muxInD_0_23_port, muxInD_0_22_port, muxInD_0_21_port, 
      muxInD_0_20_port, muxInD_0_19_port, muxInD_0_18_port, muxInD_0_17_port, 
      muxInD_0_16_port, muxInD_0_15_port, muxInD_0_14_port, muxInD_0_13_port, 
      muxInD_0_12_port, muxInD_0_11_port, muxInD_0_10_port, muxInD_0_9_port, 
      muxInD_0_8_port, muxInD_0_7_port, muxInD_0_6_port, muxInD_0_5_port, 
      muxInD_0_4_port, muxInD_0_3_port, muxInD_0_2_port, muxInD_0_1_port, 
      muxInD_0_0_port, muxInC_7_31_port, muxInC_7_30_port, muxInC_7_29_port, 
      muxInC_7_28_port, muxInC_7_27_port, muxInC_7_26_port, muxInC_7_25_port, 
      muxInC_7_24_port, muxInC_7_23_port, muxInC_7_22_port, muxInC_7_21_port, 
      muxInC_7_20_port, muxInC_7_19_port, muxInC_7_18_port, muxInC_7_17_port, 
      muxInC_7_16_port, muxInC_7_15_port, muxInC_7_14_port, muxInC_7_13_port, 
      muxInC_7_12_port, muxInC_7_11_port, muxInC_7_10_port, muxInC_7_9_port, 
      muxInC_7_8_port, muxInC_7_7_port, muxInC_7_6_port, muxInC_7_5_port, 
      muxInC_7_4_port, muxInC_7_3_port, muxInC_7_2_port, muxInC_7_1_port, 
      muxInC_7_0_port, muxInC_6_31_port, muxInC_6_30_port, muxInC_6_29_port, 
      muxInC_6_28_port, muxInC_6_27_port, muxInC_6_26_port, muxInC_6_25_port, 
      muxInC_6_24_port, muxInC_6_23_port, muxInC_6_22_port, muxInC_6_21_port, 
      muxInC_6_20_port, muxInC_6_19_port, muxInC_6_18_port, muxInC_6_17_port, 
      muxInC_6_16_port, muxInC_6_15_port, muxInC_6_14_port, muxInC_6_13_port, 
      muxInC_6_12_port, muxInC_6_11_port, muxInC_6_10_port, muxInC_6_9_port, 
      muxInC_6_8_port, muxInC_6_7_port, muxInC_6_6_port, muxInC_6_5_port, 
      muxInC_6_4_port, muxInC_6_3_port, muxInC_6_2_port, muxInC_6_1_port, 
      muxInC_6_0_port, muxInC_5_31_port, muxInC_5_30_port, muxInC_5_29_port, 
      muxInC_5_28_port, muxInC_5_27_port, muxInC_5_26_port, muxInC_5_25_port, 
      muxInC_5_24_port, muxInC_5_23_port, muxInC_5_22_port, muxInC_5_21_port, 
      muxInC_5_20_port, muxInC_5_19_port, muxInC_5_18_port, muxInC_5_17_port, 
      muxInC_5_16_port, muxInC_5_15_port, muxInC_5_14_port, muxInC_5_13_port, 
      muxInC_5_12_port, muxInC_5_11_port, muxInC_5_10_port, muxInC_5_9_port, 
      muxInC_5_8_port, muxInC_5_7_port, muxInC_5_6_port, muxInC_5_5_port, 
      muxInC_5_4_port, muxInC_5_3_port, muxInC_5_2_port, muxInC_5_1_port, 
      muxInC_5_0_port, muxInC_4_31_port, muxInC_4_30_port, muxInC_4_29_port, 
      muxInC_4_28_port, muxInC_4_27_port, muxInC_4_26_port, muxInC_4_25_port, 
      muxInC_4_24_port, muxInC_4_23_port, muxInC_4_22_port, muxInC_4_21_port, 
      muxInC_4_20_port, muxInC_4_19_port, muxInC_4_18_port, muxInC_4_17_port, 
      muxInC_4_16_port, muxInC_4_15_port, muxInC_4_14_port, muxInC_4_13_port, 
      muxInC_4_12_port, muxInC_4_11_port, muxInC_4_10_port, muxInC_4_9_port, 
      muxInC_4_8_port, muxInC_4_7_port, muxInC_4_6_port, muxInC_4_5_port, 
      muxInC_4_4_port, muxInC_4_3_port, muxInC_4_2_port, muxInC_4_1_port, 
      muxInC_4_0_port, muxInC_3_31_port, muxInC_3_30_port, muxInC_3_29_port, 
      muxInC_3_28_port, muxInC_3_27_port, muxInC_3_26_port, muxInC_3_25_port, 
      muxInC_3_24_port, muxInC_3_23_port, muxInC_3_22_port, muxInC_3_21_port, 
      muxInC_3_20_port, muxInC_3_19_port, muxInC_3_18_port, muxInC_3_17_port, 
      muxInC_3_16_port, muxInC_3_15_port, muxInC_3_14_port, muxInC_3_13_port, 
      muxInC_3_12_port, muxInC_3_11_port, muxInC_3_10_port, muxInC_3_9_port, 
      muxInC_3_8_port, muxInC_3_7_port, muxInC_3_6_port, muxInC_3_5_port, 
      muxInC_3_4_port, muxInC_3_3_port, muxInC_3_2_port, muxInC_3_1_port, 
      muxInC_3_0_port, muxInC_2_31_port, muxInC_2_30_port, muxInC_2_29_port, 
      muxInC_2_28_port, muxInC_2_27_port, muxInC_2_26_port, muxInC_2_25_port, 
      muxInC_2_24_port, muxInC_2_23_port, muxInC_2_22_port, muxInC_2_21_port, 
      muxInC_2_20_port, muxInC_2_19_port, muxInC_2_18_port, muxInC_2_17_port, 
      muxInC_2_16_port, muxInC_2_15_port, muxInC_2_14_port, muxInC_2_13_port, 
      muxInC_2_12_port, muxInC_2_11_port, muxInC_2_10_port, muxInC_2_9_port, 
      muxInC_2_8_port, muxInC_2_7_port, muxInC_2_6_port, muxInC_2_5_port, 
      muxInC_2_4_port, muxInC_2_3_port, muxInC_2_2_port, muxInC_2_1_port, 
      muxInC_2_0_port, muxInC_1_31_port, muxInC_1_30_port, muxInC_1_29_port, 
      muxInC_1_28_port, muxInC_1_27_port, muxInC_1_26_port, muxInC_1_25_port, 
      muxInC_1_24_port, muxInC_1_23_port, muxInC_1_22_port, muxInC_1_21_port, 
      muxInC_1_20_port, muxInC_1_18_port, muxInC_1_17_port, muxInC_1_16_port, 
      muxInC_1_15_port, muxInC_1_14_port, muxInC_1_13_port, muxInC_1_12_port, 
      muxInC_1_11_port, muxInC_1_10_port, muxInC_1_9_port, muxInC_1_8_port, 
      muxInC_1_7_port, muxInC_1_6_port, muxInC_1_5_port, muxInC_1_4_port, 
      muxInC_1_3_port, muxInC_1_2_port, muxInC_1_1_port, muxInC_1_0_port, 
      muxInC_0_31_port, muxInC_0_30_port, muxInC_0_29_port, muxInC_0_28_port, 
      muxInC_0_27_port, muxInC_0_26_port, muxInC_0_25_port, muxInC_0_24_port, 
      muxInC_0_23_port, muxInC_0_22_port, muxInC_0_21_port, muxInC_0_20_port, 
      muxInC_0_19_port, muxInC_0_18_port, muxInC_0_17_port, muxInC_0_16_port, 
      muxInC_0_15_port, muxInC_0_14_port, muxInC_0_13_port, muxInC_0_12_port, 
      muxInC_0_11_port, muxInC_0_10_port, muxInC_0_9_port, muxInC_0_8_port, 
      muxInC_0_7_port, muxInC_0_6_port, muxInC_0_5_port, muxInC_0_4_port, 
      muxInC_0_3_port, muxInC_0_2_port, muxInC_0_1_port, muxInC_0_0_port, 
      muxInB_7_31_port, muxInB_7_30_port, muxInB_7_29_port, muxInB_7_28_port, 
      muxInB_7_27_port, muxInB_7_26_port, muxInB_7_25_port, muxInB_7_24_port, 
      muxInB_7_23_port, muxInB_7_22_port, muxInB_7_21_port, muxInB_7_20_port, 
      muxInB_7_19_port, muxInB_7_18_port, muxInB_7_17_port, muxInB_7_16_port, 
      muxInB_7_15_port, muxInB_7_14_port, muxInB_7_13_port, muxInB_7_12_port, 
      muxInB_7_11_port, muxInB_7_10_port, muxInB_7_9_port, muxInB_7_8_port, 
      muxInB_7_7_port, muxInB_7_6_port, muxInB_7_5_port, muxInB_7_4_port, 
      muxInB_7_3_port, muxInB_7_2_port, muxInB_7_1_port, muxInB_7_0_port, 
      muxInB_6_31_port, muxInB_6_30_port, muxInB_6_29_port, muxInB_6_28_port, 
      muxInB_6_27_port, muxInB_6_26_port, muxInB_6_25_port, muxInB_6_24_port, 
      muxInB_6_23_port, muxInB_6_22_port, muxInB_6_21_port, muxInB_6_20_port, 
      muxInB_6_19_port, muxInB_6_18_port, muxInB_6_17_port, muxInB_6_16_port, 
      muxInB_6_15_port, muxInB_6_14_port, muxInB_6_13_port, muxInB_6_12_port, 
      muxInB_6_11_port, muxInB_6_10_port, muxInB_6_9_port, muxInB_6_8_port, 
      muxInB_6_7_port, muxInB_6_6_port, muxInB_6_5_port, muxInB_6_4_port, 
      muxInB_6_3_port, muxInB_6_2_port, muxInB_6_1_port, muxInB_6_0_port, 
      muxInB_5_31_port, muxInB_5_30_port, muxInB_5_29_port, muxInB_5_28_port, 
      muxInB_5_27_port, muxInB_5_26_port, muxInB_5_25_port, muxInB_5_24_port, 
      muxInB_5_23_port, muxInB_5_22_port, muxInB_5_21_port, muxInB_5_20_port, 
      muxInB_5_19_port, muxInB_5_18_port, muxInB_5_17_port, muxInB_5_16_port, 
      muxInB_5_15_port, muxInB_5_14_port, muxInB_5_13_port, muxInB_5_12_port, 
      muxInB_5_11_port, muxInB_5_10_port, muxInB_5_9_port, muxInB_5_8_port, 
      muxInB_5_7_port, muxInB_5_6_port, muxInB_5_5_port, muxInB_5_4_port, 
      muxInB_5_3_port, muxInB_5_2_port, muxInB_5_1_port, muxInB_5_0_port, 
      muxInB_4_31_port, muxInB_4_30_port, muxInB_4_29_port, muxInB_4_28_port, 
      muxInB_4_27_port, muxInB_4_26_port, muxInB_4_25_port, muxInB_4_24_port, 
      muxInB_4_23_port, muxInB_4_22_port, muxInB_4_21_port, muxInB_4_20_port, 
      muxInB_4_19_port, muxInB_4_18_port, muxInB_4_17_port, muxInB_4_16_port, 
      muxInB_4_15_port, muxInB_4_14_port, muxInB_4_13_port, muxInB_4_12_port, 
      muxInB_4_11_port, muxInB_4_10_port, muxInB_4_9_port, muxInB_4_8_port, 
      muxInB_4_7_port, muxInB_4_6_port, muxInB_4_5_port, muxInB_4_4_port, 
      muxInB_4_3_port, muxInB_4_2_port, muxInB_4_1_port, muxInB_4_0_port, 
      muxInB_3_31_port, muxInB_3_30_port, muxInB_3_29_port, muxInB_3_28_port, 
      muxInB_3_27_port, muxInB_3_26_port, muxInB_3_25_port, muxInB_3_24_port, 
      muxInB_3_23_port, muxInB_3_22_port, muxInB_3_21_port, muxInB_3_20_port, 
      muxInB_3_19_port, muxInB_3_18_port, muxInB_3_17_port, muxInB_3_16_port, 
      muxInB_3_15_port, muxInB_3_14_port, muxInB_3_13_port, muxInB_3_12_port, 
      muxInB_3_11_port, muxInB_3_10_port, muxInB_3_9_port, muxInB_3_8_port, 
      muxInB_3_7_port, muxInB_3_6_port, muxInB_3_5_port, muxInB_3_4_port, 
      muxInB_3_3_port, muxInB_3_2_port, muxInB_3_1_port, muxInB_3_0_port, 
      muxInB_2_31_port, muxInB_2_30_port, muxInB_2_29_port, muxInB_2_28_port, 
      muxInB_2_27_port, muxInB_2_26_port, muxInB_2_25_port, muxInB_2_24_port, 
      muxInB_2_23_port, muxInB_2_22_port, muxInB_2_21_port, muxInB_2_20_port, 
      muxInB_2_19_port, muxInB_2_18_port, muxInB_2_17_port, muxInB_2_16_port, 
      muxInB_2_15_port, muxInB_2_14_port, muxInB_2_13_port, muxInB_2_12_port, 
      muxInB_2_11_port, muxInB_2_10_port, muxInB_2_9_port, muxInB_2_8_port, 
      muxInB_2_7_port, muxInB_2_6_port, muxInB_2_5_port, muxInB_2_4_port, 
      muxInB_2_3_port, muxInB_2_2_port, muxInB_2_1_port, muxInB_2_0_port, 
      muxInB_1_31_port, muxInB_1_30_port, muxInB_1_29_port, muxInB_1_28_port, 
      muxInB_1_27_port, muxInB_1_26_port, muxInB_1_25_port, muxInB_1_24_port, 
      muxInB_1_23_port, muxInB_1_22_port, muxInB_1_21_port, muxInB_1_20_port, 
      muxInB_1_19_port, muxInB_1_18_port, muxInB_1_17_port, muxInB_1_16_port, 
      muxInB_1_15_port, muxInB_1_14_port, muxInB_1_13_port, muxInB_1_12_port, 
      muxInB_1_11_port, muxInB_1_10_port, muxInB_1_9_port, muxInB_1_8_port, 
      muxInB_1_7_port, muxInB_1_6_port, muxInB_1_5_port, muxInB_1_4_port, 
      muxInB_1_3_port, muxInB_1_2_port, muxInB_1_1_port, muxInB_1_0_port, 
      muxInB_0_31_port, muxInB_0_30_port, muxInB_0_29_port, muxInB_0_28_port, 
      muxInB_0_27_port, muxInB_0_26_port, muxInB_0_25_port, muxInB_0_24_port, 
      muxInB_0_23_port, muxInB_0_22_port, muxInB_0_21_port, muxInB_0_20_port, 
      muxInB_0_19_port, muxInB_0_18_port, muxInB_0_17_port, muxInB_0_16_port, 
      muxInB_0_15_port, muxInB_0_14_port, muxInB_0_13_port, muxInB_0_12_port, 
      muxInB_0_11_port, muxInB_0_10_port, muxInB_0_9_port, muxInB_0_8_port, 
      muxInB_0_7_port, muxInB_0_6_port, muxInB_0_5_port, muxInB_0_4_port, 
      muxInB_0_3_port, muxInB_0_2_port, muxInB_0_1_port, muxInB_0_0_port, 
      outmux_7_31_port, outmux_7_30_port, outmux_7_29_port, outmux_7_28_port, 
      outmux_7_27_port, outmux_7_26_port, outmux_7_25_port, outmux_7_24_port, 
      outmux_7_23_port, outmux_7_22_port, outmux_7_21_port, outmux_7_20_port, 
      outmux_7_19_port, outmux_7_18_port, outmux_7_17_port, outmux_7_16_port, 
      outmux_7_15_port, outmux_7_14_port, outmux_7_13_port, outmux_7_12_port, 
      outmux_7_11_port, outmux_7_10_port, outmux_7_9_port, outmux_7_8_port, 
      outmux_7_7_port, outmux_7_6_port, outmux_7_5_port, outmux_7_4_port, 
      outmux_7_3_port, outmux_7_2_port, outmux_7_1_port, outmux_7_0_port, 
      outmux_6_31_port, outmux_6_30_port, outmux_6_29_port, outmux_6_28_port, 
      outmux_6_27_port, outmux_6_26_port, outmux_6_25_port, outmux_6_24_port, 
      outmux_6_23_port, outmux_6_22_port, outmux_6_21_port, outmux_6_20_port, 
      outmux_6_19_port, outmux_6_18_port, outmux_6_17_port, outmux_6_16_port, 
      outmux_6_15_port, outmux_6_14_port, outmux_6_13_port, outmux_6_12_port, 
      outmux_6_11_port, outmux_6_10_port, outmux_6_9_port, outmux_6_8_port, 
      outmux_6_7_port, outmux_6_6_port, outmux_6_5_port, outmux_6_4_port, 
      outmux_6_3_port, outmux_6_2_port, outmux_6_1_port, outmux_6_0_port, 
      outmux_5_31_port, outmux_5_30_port, outmux_5_29_port, outmux_5_28_port, 
      outmux_5_27_port, outmux_5_26_port, outmux_5_25_port, outmux_5_24_port, 
      outmux_5_23_port, outmux_5_22_port, outmux_5_21_port, outmux_5_20_port, 
      outmux_5_19_port, outmux_5_18_port, outmux_5_17_port, outmux_5_16_port, 
      outmux_5_15_port, outmux_5_14_port, outmux_5_13_port, outmux_5_12_port, 
      outmux_5_11_port, outmux_5_10_port, outmux_5_9_port, outmux_5_8_port, 
      outmux_5_7_port, outmux_5_6_port, outmux_5_5_port, outmux_5_4_port, 
      outmux_5_3_port, outmux_5_2_port, outmux_5_1_port, outmux_5_0_port, 
      outmux_4_31_port, outmux_4_30_port, outmux_4_29_port, outmux_4_28_port, 
      outmux_4_27_port, outmux_4_26_port, outmux_4_25_port, outmux_4_24_port, 
      outmux_4_23_port, outmux_4_22_port, outmux_4_21_port, outmux_4_20_port, 
      outmux_4_19_port, outmux_4_18_port, outmux_4_17_port, outmux_4_16_port, 
      outmux_4_15_port, outmux_4_14_port, outmux_4_13_port, outmux_4_12_port, 
      outmux_4_11_port, outmux_4_10_port, outmux_4_9_port, outmux_4_8_port, 
      outmux_4_7_port, outmux_4_6_port, outmux_4_5_port, outmux_4_4_port, 
      outmux_4_3_port, outmux_4_2_port, outmux_4_1_port, outmux_4_0_port, 
      outmux_3_31_port, outmux_3_30_port, outmux_3_29_port, outmux_3_28_port, 
      outmux_3_27_port, outmux_3_26_port, outmux_3_25_port, outmux_3_24_port, 
      outmux_3_23_port, outmux_3_22_port, outmux_3_21_port, outmux_3_20_port, 
      outmux_3_19_port, outmux_3_18_port, outmux_3_17_port, outmux_3_16_port, 
      outmux_3_15_port, outmux_3_14_port, outmux_3_13_port, outmux_3_12_port, 
      outmux_3_11_port, outmux_3_10_port, outmux_3_9_port, outmux_3_8_port, 
      outmux_3_7_port, outmux_3_6_port, outmux_3_5_port, outmux_3_4_port, 
      outmux_3_3_port, outmux_3_2_port, outmux_3_1_port, outmux_3_0_port, 
      outmux_2_31_port, outmux_2_30_port, outmux_2_29_port, outmux_2_28_port, 
      outmux_2_27_port, outmux_2_26_port, outmux_2_25_port, outmux_2_24_port, 
      outmux_2_23_port, outmux_2_22_port, outmux_2_21_port, outmux_2_20_port, 
      outmux_2_19_port, outmux_2_18_port, outmux_2_17_port, outmux_2_16_port, 
      outmux_2_15_port, outmux_2_14_port, outmux_2_13_port, outmux_2_12_port, 
      outmux_2_11_port, outmux_2_10_port, outmux_2_9_port, outmux_2_8_port, 
      outmux_2_7_port, outmux_2_6_port, outmux_2_5_port, outmux_2_4_port, 
      outmux_2_3_port, outmux_2_2_port, outmux_2_1_port, outmux_2_0_port, 
      outmux_1_31_port, outmux_1_30_port, outmux_1_29_port, outmux_1_28_port, 
      outmux_1_27_port, outmux_1_26_port, outmux_1_25_port, outmux_1_24_port, 
      outmux_1_23_port, outmux_1_22_port, outmux_1_21_port, outmux_1_20_port, 
      outmux_1_19_port, outmux_1_18_port, outmux_1_17_port, outmux_1_16_port, 
      outmux_1_15_port, outmux_1_14_port, outmux_1_13_port, outmux_1_12_port, 
      outmux_1_11_port, outmux_1_10_port, outmux_1_9_port, outmux_1_8_port, 
      outmux_1_7_port, outmux_1_6_port, outmux_1_5_port, outmux_1_4_port, 
      outmux_1_3_port, outmux_1_2_port, outmux_1_1_port, outmux_1_0_port, 
      outmux_0_31_port, outmux_0_30_port, outmux_0_29_port, outmux_0_28_port, 
      outmux_0_27_port, outmux_0_26_port, outmux_0_25_port, outmux_0_24_port, 
      outmux_0_23_port, outmux_0_22_port, outmux_0_21_port, outmux_0_20_port, 
      outmux_0_19_port, outmux_0_18_port, outmux_0_17_port, outmux_0_16_port, 
      outmux_0_15_port, outmux_0_14_port, outmux_0_13_port, outmux_0_12_port, 
      outmux_0_11_port, outmux_0_10_port, outmux_0_9_port, outmux_0_8_port, 
      outmux_0_7_port, outmux_0_6_port, outmux_0_5_port, outmux_0_4_port, 
      outmux_0_3_port, outmux_0_2_port, outmux_0_1_port, outmux_0_0_port, 
      cout_array_5_31_port, cout_array_5_30_port, cout_array_5_29_port, 
      cout_array_5_28_port, cout_array_5_27_port, cout_array_5_26_port, 
      cout_array_5_25_port, cout_array_5_24_port, cout_array_5_23_port, 
      cout_array_5_22_port, cout_array_5_21_port, cout_array_5_20_port, 
      cout_array_5_19_port, cout_array_5_18_port, cout_array_5_17_port, 
      cout_array_5_16_port, cout_array_5_15_port, cout_array_5_14_port, 
      cout_array_5_13_port, cout_array_5_12_port, cout_array_5_11_port, 
      cout_array_5_10_port, cout_array_5_9_port, cout_array_5_8_port, 
      cout_array_5_7_port, cout_array_5_6_port, cout_array_5_5_port, 
      cout_array_5_4_port, cout_array_5_3_port, cout_array_5_2_port, 
      cout_array_5_1_port, cout_array_5_0_port, cout_array_4_31_port, 
      cout_array_4_30_port, cout_array_4_29_port, cout_array_4_28_port, 
      cout_array_4_27_port, cout_array_4_26_port, cout_array_4_25_port, 
      cout_array_4_24_port, cout_array_4_23_port, cout_array_4_22_port, 
      cout_array_4_21_port, cout_array_4_20_port, cout_array_4_19_port, 
      cout_array_4_18_port, cout_array_4_17_port, cout_array_4_16_port, 
      cout_array_4_15_port, cout_array_4_14_port, cout_array_4_13_port, 
      cout_array_4_12_port, cout_array_4_11_port, cout_array_4_10_port, 
      cout_array_4_9_port, cout_array_4_8_port, cout_array_4_7_port, 
      cout_array_4_6_port, cout_array_4_5_port, cout_array_4_4_port, 
      cout_array_4_3_port, cout_array_4_2_port, cout_array_4_1_port, 
      cout_array_4_0_port, cout_array_3_31_port, cout_array_3_30_port, 
      cout_array_3_29_port, cout_array_3_28_port, cout_array_3_27_port, 
      cout_array_3_26_port, cout_array_3_25_port, cout_array_3_24_port, 
      cout_array_3_23_port, cout_array_3_22_port, cout_array_3_21_port, 
      cout_array_3_20_port, cout_array_3_19_port, cout_array_3_18_port, 
      cout_array_3_17_port, cout_array_3_16_port, cout_array_3_15_port, 
      cout_array_3_14_port, cout_array_3_13_port, cout_array_3_12_port, 
      cout_array_3_11_port, cout_array_3_10_port, cout_array_3_9_port, 
      cout_array_3_8_port, cout_array_3_7_port, cout_array_3_6_port, 
      cout_array_3_5_port, cout_array_3_4_port, cout_array_3_3_port, 
      cout_array_3_2_port, cout_array_3_1_port, cout_array_3_0_port, 
      cout_array_2_31_port, cout_array_2_30_port, cout_array_2_29_port, 
      cout_array_2_28_port, cout_array_2_27_port, cout_array_2_26_port, 
      cout_array_2_25_port, cout_array_2_24_port, cout_array_2_23_port, 
      cout_array_2_22_port, cout_array_2_21_port, cout_array_2_20_port, 
      cout_array_2_19_port, cout_array_2_18_port, cout_array_2_17_port, 
      cout_array_2_16_port, cout_array_2_15_port, cout_array_2_14_port, 
      cout_array_2_13_port, cout_array_2_12_port, cout_array_2_11_port, 
      cout_array_2_10_port, cout_array_2_9_port, cout_array_2_8_port, 
      cout_array_2_7_port, cout_array_2_6_port, cout_array_2_5_port, 
      cout_array_2_4_port, cout_array_2_3_port, cout_array_2_2_port, 
      cout_array_2_1_port, cout_array_2_0_port, cout_array_1_31_port, 
      cout_array_1_30_port, cout_array_1_29_port, cout_array_1_28_port, 
      cout_array_1_27_port, cout_array_1_26_port, cout_array_1_25_port, 
      cout_array_1_24_port, cout_array_1_23_port, cout_array_1_22_port, 
      cout_array_1_21_port, cout_array_1_20_port, cout_array_1_19_port, 
      cout_array_1_18_port, cout_array_1_17_port, cout_array_1_16_port, 
      cout_array_1_15_port, cout_array_1_14_port, cout_array_1_13_port, 
      cout_array_1_12_port, cout_array_1_11_port, cout_array_1_10_port, 
      cout_array_1_9_port, cout_array_1_8_port, cout_array_1_7_port, 
      cout_array_1_6_port, cout_array_1_5_port, cout_array_1_4_port, 
      cout_array_1_3_port, cout_array_1_2_port, cout_array_1_1_port, 
      cout_array_1_0_port, cout_array_0_31_port, cout_array_0_30_port, 
      cout_array_0_29_port, cout_array_0_28_port, cout_array_0_27_port, 
      cout_array_0_26_port, cout_array_0_25_port, cout_array_0_24_port, 
      cout_array_0_23_port, cout_array_0_22_port, cout_array_0_21_port, 
      cout_array_0_20_port, cout_array_0_19_port, cout_array_0_18_port, 
      cout_array_0_17_port, cout_array_0_16_port, cout_array_0_15_port, 
      cout_array_0_14_port, cout_array_0_13_port, cout_array_0_12_port, 
      cout_array_0_11_port, cout_array_0_10_port, cout_array_0_9_port, 
      cout_array_0_8_port, cout_array_0_7_port, cout_array_0_6_port, 
      cout_array_0_5_port, cout_array_0_4_port, cout_array_0_3_port, 
      cout_array_0_2_port, cout_array_0_1_port, cout_array_0_0_port, 
      sum_array_5_31_port, sum_array_5_30_port, sum_array_5_29_port, 
      sum_array_5_28_port, sum_array_5_27_port, sum_array_5_26_port, 
      sum_array_5_25_port, sum_array_5_24_port, sum_array_5_23_port, 
      sum_array_5_22_port, sum_array_5_21_port, sum_array_5_20_port, 
      sum_array_5_19_port, sum_array_5_18_port, sum_array_5_17_port, 
      sum_array_5_16_port, sum_array_5_15_port, sum_array_5_14_port, 
      sum_array_5_13_port, sum_array_5_12_port, sum_array_5_11_port, 
      sum_array_5_10_port, sum_array_5_9_port, sum_array_5_8_port, 
      sum_array_5_7_port, sum_array_5_6_port, sum_array_5_5_port, 
      sum_array_5_4_port, sum_array_5_3_port, sum_array_5_2_port, 
      sum_array_5_1_port, sum_array_5_0_port, sum_array_4_31_port, 
      sum_array_4_30_port, sum_array_4_29_port, sum_array_4_28_port, 
      sum_array_4_27_port, sum_array_4_26_port, sum_array_4_25_port, 
      sum_array_4_24_port, sum_array_4_23_port, sum_array_4_22_port, 
      sum_array_4_21_port, sum_array_4_20_port, sum_array_4_19_port, 
      sum_array_4_18_port, sum_array_4_17_port, sum_array_4_16_port, 
      sum_array_4_15_port, sum_array_4_14_port, sum_array_4_13_port, 
      sum_array_4_12_port, sum_array_4_11_port, sum_array_4_10_port, 
      sum_array_4_9_port, sum_array_4_8_port, sum_array_4_7_port, 
      sum_array_4_6_port, sum_array_4_5_port, sum_array_4_4_port, 
      sum_array_4_3_port, sum_array_4_2_port, sum_array_4_1_port, 
      sum_array_4_0_port, sum_array_3_31_port, sum_array_3_30_port, 
      sum_array_3_29_port, sum_array_3_28_port, sum_array_3_27_port, 
      sum_array_3_26_port, sum_array_3_25_port, sum_array_3_24_port, 
      sum_array_3_23_port, sum_array_3_22_port, sum_array_3_21_port, 
      sum_array_3_20_port, sum_array_3_19_port, sum_array_3_18_port, 
      sum_array_3_17_port, sum_array_3_16_port, sum_array_3_15_port, 
      sum_array_3_14_port, sum_array_3_13_port, sum_array_3_12_port, 
      sum_array_3_11_port, sum_array_3_10_port, sum_array_3_9_port, 
      sum_array_3_8_port, sum_array_3_7_port, sum_array_3_6_port, 
      sum_array_3_5_port, sum_array_3_4_port, sum_array_3_3_port, 
      sum_array_3_2_port, sum_array_3_1_port, sum_array_3_0_port, 
      sum_array_2_31_port, sum_array_2_30_port, sum_array_2_29_port, 
      sum_array_2_28_port, sum_array_2_27_port, sum_array_2_26_port, 
      sum_array_2_25_port, sum_array_2_24_port, sum_array_2_23_port, 
      sum_array_2_22_port, sum_array_2_21_port, sum_array_2_20_port, 
      sum_array_2_19_port, sum_array_2_18_port, sum_array_2_17_port, 
      sum_array_2_16_port, sum_array_2_15_port, sum_array_2_14_port, 
      sum_array_2_13_port, sum_array_2_12_port, sum_array_2_11_port, 
      sum_array_2_10_port, sum_array_2_9_port, sum_array_2_8_port, 
      sum_array_2_7_port, sum_array_2_6_port, sum_array_2_5_port, 
      sum_array_2_4_port, sum_array_2_3_port, sum_array_2_2_port, 
      sum_array_2_1_port, sum_array_2_0_port, sum_array_1_31_port, 
      sum_array_1_30_port, sum_array_1_29_port, sum_array_1_28_port, 
      sum_array_1_27_port, sum_array_1_26_port, sum_array_1_25_port, 
      sum_array_1_24_port, sum_array_1_23_port, sum_array_1_22_port, 
      sum_array_1_21_port, sum_array_1_20_port, sum_array_1_19_port, 
      sum_array_1_18_port, sum_array_1_17_port, sum_array_1_16_port, 
      sum_array_1_15_port, sum_array_1_14_port, sum_array_1_13_port, 
      sum_array_1_12_port, sum_array_1_11_port, sum_array_1_10_port, 
      sum_array_1_9_port, sum_array_1_8_port, sum_array_1_7_port, 
      sum_array_1_6_port, sum_array_1_5_port, sum_array_1_4_port, 
      sum_array_1_3_port, sum_array_1_2_port, sum_array_1_1_port, 
      sum_array_1_0_port, sum_array_0_31_port, sum_array_0_30_port, 
      sum_array_0_29_port, sum_array_0_28_port, sum_array_0_27_port, 
      sum_array_0_26_port, sum_array_0_25_port, sum_array_0_24_port, 
      sum_array_0_23_port, sum_array_0_22_port, sum_array_0_21_port, 
      sum_array_0_20_port, sum_array_0_19_port, sum_array_0_18_port, 
      sum_array_0_17_port, sum_array_0_16_port, sum_array_0_15_port, 
      sum_array_0_14_port, sum_array_0_13_port, sum_array_0_12_port, 
      sum_array_0_11_port, sum_array_0_10_port, sum_array_0_9_port, 
      sum_array_0_8_port, sum_array_0_7_port, sum_array_0_6_port, 
      sum_array_0_5_port, sum_array_0_4_port, sum_array_0_3_port, 
      sum_array_0_2_port, sum_array_0_1_port, sum_array_0_0_port, net6197, n20,
      net51440, net51450, net51451, net51452, n2, n3, n10, n11, n13, n14, n15, 
      n17, n18, n19, n21, n22, n25, n26, n27, n28, net59829, net59830, net59831
      , net59832, net59833, net59834, net59835, net59836, net59837, net59838, 
      net59839, net59840, net59841, net59842, net59843, net59844, net59845, 
      net59846, net59847, net59848, net59849, net59850, net59851, net59852, 
      net59853, net59854, net59855, net59856, net59857, net59858, net59859, 
      net59860, net59861, net59862, net59863, net59864, net59865, net59866, 
      net59867, net59868, net59869, net59870, net59871, net59872, net59873, 
      net59874, net59875, net59876, net59877, net59878, net59879, net59880, 
      net59881, net59882, net59883, net59884, net59885, net59886, net59887, 
      net59888, net59889, net59890, net59891, net59892, net59893, net59894, 
      net59895, net59896, net59897, net59898, net59899, net59900, net59901, 
      net59902, net59903, net59904, net59905, net59906, net59907, net59908, 
      net59909, net59910, net59911, net59912, net59913, net59914, net59915, 
      net59916, net59917, net59918, net59919, net59920, net59921, net59922, 
      net59923, net59924, net59925, net59926, net59927, net59928, net59929, 
      net59930, net59931, net59932, net59933, net59934, net59935, net59936, 
      net59937, net59938, net59939, net59940, net59941, net59942, net59943, 
      net59944, net59945, net59946, net59947, net59948, net59949, net59950, 
      net59951, net59952, net59953, net59954, net59955, net59956, net59957, 
      net59958, net59959, net59960, net59961, net59962, net59963, net59964, 
      net59965, net59966, net59967, net59968, net59969, net59970, net59971, 
      net59972, net59973, net59974, net59975, net59976, net59977, net59978, 
      net59979, net59980, net59981, net59982, net59983, net59984, net59985, 
      net59986, net59987, net59988, net59989, net59990, net59991, net59992, 
      net59993, net59994, net59995, net59996, net59997, net59998, net59999, 
      net60000, net60001, net60002, net60003, net60004, net60005, net60006, 
      net60007, net60008, net60009, net60010, net60011, net60012, net60013, 
      net60014, net60015, net60016, net60017, net60018, net60019, net60020, 
      net60021, net60022, net60023, net60024, net60025, net60026, net60027, 
      net60028, net60029, net60030, net60031, net60032, net60033, net60034, 
      net60035, net60036, net60037, net60038, net60039, net60040, net60041, 
      net60042, net60043, net60044, net60045, net60046, net60047, net60048, 
      net60049, net60050, net60051, net60052, net60053, net60054, net60055, 
      net60056, net60057, net60058, net60059, net60060, net60061, net60062, 
      net60063, net60064, net60065, net60066, net60067, net60068, net60069, 
      net60070, net60071, net60072, net60073, net60074 : std_logic;

begin
   
   X_Logic0_port <= '0';
   SHIFTERS_0 : shift_mul_N16_S0 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_0_31_port, B(30)
                           => muxInB_0_30_port, B(29) => muxInB_0_29_port, 
                           B(28) => muxInB_0_28_port, B(27) => muxInB_0_27_port
                           , B(26) => muxInB_0_26_port, B(25) => 
                           muxInB_0_25_port, B(24) => muxInB_0_24_port, B(23) 
                           => muxInB_0_23_port, B(22) => muxInB_0_22_port, 
                           B(21) => muxInB_0_21_port, B(20) => muxInB_0_20_port
                           , B(19) => muxInB_0_19_port, B(18) => 
                           muxInB_0_18_port, B(17) => muxInB_0_17_port, B(16) 
                           => muxInB_0_16_port, B(15) => muxInB_0_15_port, 
                           B(14) => muxInB_0_14_port, B(13) => muxInB_0_13_port
                           , B(12) => muxInB_0_12_port, B(11) => 
                           muxInB_0_11_port, B(10) => muxInB_0_10_port, B(9) =>
                           muxInB_0_9_port, B(8) => muxInB_0_8_port, B(7) => 
                           muxInB_0_7_port, B(6) => muxInB_0_6_port, B(5) => 
                           muxInB_0_5_port, B(4) => muxInB_0_4_port, B(3) => 
                           muxInB_0_3_port, B(2) => muxInB_0_2_port, B(1) => 
                           muxInB_0_1_port, B(0) => muxInB_0_0_port, C(31) => 
                           muxInC_0_31_port, C(30) => muxInC_0_30_port, C(29) 
                           => muxInC_0_29_port, C(28) => muxInC_0_28_port, 
                           C(27) => muxInC_0_27_port, C(26) => muxInC_0_26_port
                           , C(25) => muxInC_0_25_port, C(24) => 
                           muxInC_0_24_port, C(23) => muxInC_0_23_port, C(22) 
                           => muxInC_0_22_port, C(21) => muxInC_0_21_port, 
                           C(20) => muxInC_0_20_port, C(19) => muxInC_0_19_port
                           , C(18) => muxInC_0_18_port, C(17) => 
                           muxInC_0_17_port, C(16) => muxInC_0_16_port, C(15) 
                           => muxInC_0_15_port, C(14) => muxInC_0_14_port, 
                           C(13) => muxInC_0_13_port, C(12) => muxInC_0_12_port
                           , C(11) => muxInC_0_11_port, C(10) => 
                           muxInC_0_10_port, C(9) => muxInC_0_9_port, C(8) => 
                           muxInC_0_8_port, C(7) => muxInC_0_7_port, C(6) => 
                           muxInC_0_6_port, C(5) => muxInC_0_5_port, C(4) => 
                           muxInC_0_4_port, C(3) => muxInC_0_3_port, C(2) => 
                           muxInC_0_2_port, C(1) => muxInC_0_1_port, C(0) => 
                           muxInC_0_0_port, D(31) => muxInD_0_31_port, D(30) =>
                           muxInD_0_30_port, D(29) => muxInD_0_29_port, D(28) 
                           => muxInD_0_28_port, D(27) => muxInD_0_27_port, 
                           D(26) => muxInD_0_26_port, D(25) => muxInD_0_25_port
                           , D(24) => muxInD_0_24_port, D(23) => 
                           muxInD_0_23_port, D(22) => muxInD_0_22_port, D(21) 
                           => muxInD_0_21_port, D(20) => muxInD_0_20_port, 
                           D(19) => muxInD_0_19_port, D(18) => muxInD_0_18_port
                           , D(17) => muxInD_0_17_port, D(16) => 
                           muxInD_0_16_port, D(15) => muxInD_0_15_port, D(14) 
                           => muxInD_0_14_port, D(13) => muxInD_0_13_port, 
                           D(12) => muxInD_0_12_port, D(11) => muxInD_0_11_port
                           , D(10) => muxInD_0_10_port, D(9) => muxInD_0_9_port
                           , D(8) => muxInD_0_8_port, D(7) => muxInD_0_7_port, 
                           D(6) => muxInD_0_6_port, D(5) => muxInD_0_5_port, 
                           D(4) => muxInD_0_4_port, D(3) => muxInD_0_3_port, 
                           D(2) => muxInD_0_2_port, D(1) => muxInD_0_1_port, 
                           D(0) => net60073, E(31) => muxInE_0_31_port, E(30) 
                           => muxInE_0_30_port, E(29) => muxInE_0_29_port, 
                           E(28) => muxInE_0_28_port, E(27) => muxInE_0_27_port
                           , E(26) => muxInE_0_26_port, E(25) => net51450, 
                           E(24) => muxInE_0_24_port, E(23) => muxInE_0_23_port
                           , E(22) => net51451, E(21) => muxInE_0_21_port, 
                           E(20) => muxInE_0_20_port, E(19) => muxInE_0_19_port
                           , E(18) => muxInE_0_18_port, E(17) => net51452, 
                           E(16) => muxInE_0_16_port, E(15) => muxInE_0_15_port
                           , E(14) => muxInE_0_14_port, E(13) => 
                           muxInE_0_13_port, E(12) => muxInE_0_12_port, E(11) 
                           => muxInE_0_11_port, E(10) => muxInE_0_10_port, E(9)
                           => muxInE_0_9_port, E(8) => muxInE_0_8_port, E(7) =>
                           muxInE_0_7_port, E(6) => muxInE_0_6_port, E(5) => 
                           muxInE_0_5_port, E(4) => muxInE_0_4_port, E(3) => 
                           muxInE_0_3_port, E(2) => muxInE_0_2_port, E(1) => 
                           muxInE_0_1_port, E(0) => net60074);
   SHIFTERS_1 : shift_mul_N16_S2 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_1_31_port, B(30)
                           => muxInB_1_30_port, B(29) => muxInB_1_29_port, 
                           B(28) => muxInB_1_28_port, B(27) => muxInB_1_27_port
                           , B(26) => muxInB_1_26_port, B(25) => 
                           muxInB_1_25_port, B(24) => muxInB_1_24_port, B(23) 
                           => muxInB_1_23_port, B(22) => muxInB_1_22_port, 
                           B(21) => muxInB_1_21_port, B(20) => muxInB_1_20_port
                           , B(19) => muxInB_1_19_port, B(18) => 
                           muxInB_1_18_port, B(17) => muxInB_1_17_port, B(16) 
                           => muxInB_1_16_port, B(15) => muxInB_1_15_port, 
                           B(14) => muxInB_1_14_port, B(13) => muxInB_1_13_port
                           , B(12) => muxInB_1_12_port, B(11) => 
                           muxInB_1_11_port, B(10) => muxInB_1_10_port, B(9) =>
                           muxInB_1_9_port, B(8) => muxInB_1_8_port, B(7) => 
                           muxInB_1_7_port, B(6) => muxInB_1_6_port, B(5) => 
                           muxInB_1_5_port, B(4) => muxInB_1_4_port, B(3) => 
                           muxInB_1_3_port, B(2) => muxInB_1_2_port, B(1) => 
                           net60063, B(0) => net60064, C(31) => 
                           muxInC_1_31_port, C(30) => muxInC_1_30_port, C(29) 
                           => muxInC_1_29_port, C(28) => muxInC_1_28_port, 
                           C(27) => muxInC_1_27_port, C(26) => muxInC_1_26_port
                           , C(25) => muxInC_1_25_port, C(24) => 
                           muxInC_1_24_port, C(23) => muxInC_1_23_port, C(22) 
                           => muxInC_1_22_port, C(21) => muxInC_1_21_port, 
                           C(20) => muxInC_1_20_port, C(19) => net51440, C(18) 
                           => muxInC_1_18_port, C(17) => muxInC_1_17_port, 
                           C(16) => muxInC_1_16_port, C(15) => muxInC_1_15_port
                           , C(14) => muxInC_1_14_port, C(13) => 
                           muxInC_1_13_port, C(12) => muxInC_1_12_port, C(11) 
                           => muxInC_1_11_port, C(10) => muxInC_1_10_port, C(9)
                           => muxInC_1_9_port, C(8) => muxInC_1_8_port, C(7) =>
                           muxInC_1_7_port, C(6) => muxInC_1_6_port, C(5) => 
                           muxInC_1_5_port, C(4) => muxInC_1_4_port, C(3) => 
                           muxInC_1_3_port, C(2) => muxInC_1_2_port, C(1) => 
                           net60065, C(0) => net60066, D(31) => 
                           muxInD_1_31_port, D(30) => muxInD_1_30_port, D(29) 
                           => muxInD_1_29_port, D(28) => muxInD_1_28_port, 
                           D(27) => muxInD_1_27_port, D(26) => muxInD_1_26_port
                           , D(25) => muxInD_1_25_port, D(24) => 
                           muxInD_1_24_port, D(23) => muxInD_1_23_port, D(22) 
                           => muxInD_1_22_port, D(21) => muxInD_1_21_port, 
                           D(20) => muxInD_1_20_port, D(19) => muxInD_1_19_port
                           , D(18) => muxInD_1_18_port, D(17) => 
                           muxInD_1_17_port, D(16) => muxInD_1_16_port, D(15) 
                           => muxInD_1_15_port, D(14) => muxInD_1_14_port, 
                           D(13) => muxInD_1_13_port, D(12) => muxInD_1_12_port
                           , D(11) => muxInD_1_11_port, D(10) => 
                           muxInD_1_10_port, D(9) => muxInD_1_9_port, D(8) => 
                           muxInD_1_8_port, D(7) => muxInD_1_7_port, D(6) => 
                           muxInD_1_6_port, D(5) => muxInD_1_5_port, D(4) => 
                           muxInD_1_4_port, D(3) => muxInD_1_3_port, D(2) => 
                           net60067, D(1) => net60068, D(0) => net60069, E(31) 
                           => muxInE_1_31_port, E(30) => muxInE_1_30_port, 
                           E(29) => muxInE_1_29_port, E(28) => muxInE_1_28_port
                           , E(27) => muxInE_1_27_port, E(26) => 
                           muxInE_1_26_port, E(25) => muxInE_1_25_port, E(24) 
                           => muxInE_1_24_port, E(23) => muxInE_1_23_port, 
                           E(22) => muxInE_1_22_port, E(21) => muxInE_1_21_port
                           , E(20) => muxInE_1_20_port, E(19) => 
                           muxInE_1_19_port, E(18) => muxInE_1_18_port, E(17) 
                           => muxInE_1_17_port, E(16) => muxInE_1_16_port, 
                           E(15) => muxInE_1_15_port, E(14) => muxInE_1_14_port
                           , E(13) => muxInE_1_13_port, E(12) => 
                           muxInE_1_12_port, E(11) => muxInE_1_11_port, E(10) 
                           => muxInE_1_10_port, E(9) => muxInE_1_9_port, E(8) 
                           => muxInE_1_8_port, E(7) => muxInE_1_7_port, E(6) =>
                           muxInE_1_6_port, E(5) => muxInE_1_5_port, E(4) => 
                           muxInE_1_4_port, E(3) => muxInE_1_3_port, E(2) => 
                           net60070, E(1) => net60071, E(0) => net60072);
   SHIFTERS_2 : shift_mul_N16_S4 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_2_31_port, B(30)
                           => muxInB_2_30_port, B(29) => muxInB_2_29_port, 
                           B(28) => muxInB_2_28_port, B(27) => muxInB_2_27_port
                           , B(26) => muxInB_2_26_port, B(25) => 
                           muxInB_2_25_port, B(24) => muxInB_2_24_port, B(23) 
                           => muxInB_2_23_port, B(22) => muxInB_2_22_port, 
                           B(21) => muxInB_2_21_port, B(20) => muxInB_2_20_port
                           , B(19) => muxInB_2_19_port, B(18) => 
                           muxInB_2_18_port, B(17) => muxInB_2_17_port, B(16) 
                           => muxInB_2_16_port, B(15) => muxInB_2_15_port, 
                           B(14) => muxInB_2_14_port, B(13) => muxInB_2_13_port
                           , B(12) => muxInB_2_12_port, B(11) => 
                           muxInB_2_11_port, B(10) => muxInB_2_10_port, B(9) =>
                           muxInB_2_9_port, B(8) => muxInB_2_8_port, B(7) => 
                           muxInB_2_7_port, B(6) => muxInB_2_6_port, B(5) => 
                           muxInB_2_5_port, B(4) => muxInB_2_4_port, B(3) => 
                           net60045, B(2) => net60046, B(1) => net60047, B(0) 
                           => net60048, C(31) => muxInC_2_31_port, C(30) => 
                           muxInC_2_30_port, C(29) => muxInC_2_29_port, C(28) 
                           => muxInC_2_28_port, C(27) => muxInC_2_27_port, 
                           C(26) => muxInC_2_26_port, C(25) => muxInC_2_25_port
                           , C(24) => muxInC_2_24_port, C(23) => 
                           muxInC_2_23_port, C(22) => muxInC_2_22_port, C(21) 
                           => muxInC_2_21_port, C(20) => muxInC_2_20_port, 
                           C(19) => muxInC_2_19_port, C(18) => muxInC_2_18_port
                           , C(17) => muxInC_2_17_port, C(16) => 
                           muxInC_2_16_port, C(15) => muxInC_2_15_port, C(14) 
                           => muxInC_2_14_port, C(13) => muxInC_2_13_port, 
                           C(12) => muxInC_2_12_port, C(11) => muxInC_2_11_port
                           , C(10) => muxInC_2_10_port, C(9) => muxInC_2_9_port
                           , C(8) => muxInC_2_8_port, C(7) => muxInC_2_7_port, 
                           C(6) => muxInC_2_6_port, C(5) => muxInC_2_5_port, 
                           C(4) => muxInC_2_4_port, C(3) => net60049, C(2) => 
                           net60050, C(1) => net60051, C(0) => net60052, D(31) 
                           => muxInD_2_31_port, D(30) => muxInD_2_30_port, 
                           D(29) => muxInD_2_29_port, D(28) => muxInD_2_28_port
                           , D(27) => muxInD_2_27_port, D(26) => 
                           muxInD_2_26_port, D(25) => muxInD_2_25_port, D(24) 
                           => muxInD_2_24_port, D(23) => muxInD_2_23_port, 
                           D(22) => muxInD_2_22_port, D(21) => muxInD_2_21_port
                           , D(20) => muxInD_2_20_port, D(19) => 
                           muxInD_2_19_port, D(18) => muxInD_2_18_port, D(17) 
                           => muxInD_2_17_port, D(16) => muxInD_2_16_port, 
                           D(15) => muxInD_2_15_port, D(14) => muxInD_2_14_port
                           , D(13) => muxInD_2_13_port, D(12) => 
                           muxInD_2_12_port, D(11) => muxInD_2_11_port, D(10) 
                           => muxInD_2_10_port, D(9) => muxInD_2_9_port, D(8) 
                           => muxInD_2_8_port, D(7) => muxInD_2_7_port, D(6) =>
                           muxInD_2_6_port, D(5) => muxInD_2_5_port, D(4) => 
                           net60053, D(3) => net60054, D(2) => net60055, D(1) 
                           => net60056, D(0) => net60057, E(31) => 
                           muxInE_2_31_port, E(30) => muxInE_2_30_port, E(29) 
                           => muxInE_2_29_port, E(28) => muxInE_2_28_port, 
                           E(27) => muxInE_2_27_port, E(26) => muxInE_2_26_port
                           , E(25) => muxInE_2_25_port, E(24) => 
                           muxInE_2_24_port, E(23) => muxInE_2_23_port, E(22) 
                           => muxInE_2_22_port, E(21) => muxInE_2_21_port, 
                           E(20) => n20, E(19) => muxInE_2_19_port, E(18) => 
                           muxInE_2_18_port, E(17) => muxInE_2_17_port, E(16) 
                           => muxInE_2_16_port, E(15) => muxInE_2_15_port, 
                           E(14) => muxInE_2_14_port, E(13) => muxInE_2_13_port
                           , E(12) => muxInE_2_12_port, E(11) => 
                           muxInE_2_11_port, E(10) => muxInE_2_10_port, E(9) =>
                           muxInE_2_9_port, E(8) => muxInE_2_8_port, E(7) => 
                           muxInE_2_7_port, E(6) => muxInE_2_6_port, E(5) => 
                           muxInE_2_5_port, E(4) => net60058, E(3) => net60059,
                           E(2) => net60060, E(1) => net60061, E(0) => net60062
                           );
   SHIFTERS_3 : shift_mul_N16_S6 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n3, B(31) => muxInB_3_31_port, B(30)
                           => muxInB_3_30_port, B(29) => muxInB_3_29_port, 
                           B(28) => muxInB_3_28_port, B(27) => muxInB_3_27_port
                           , B(26) => muxInB_3_26_port, B(25) => 
                           muxInB_3_25_port, B(24) => muxInB_3_24_port, B(23) 
                           => muxInB_3_23_port, B(22) => muxInB_3_22_port, 
                           B(21) => muxInB_3_21_port, B(20) => muxInB_3_20_port
                           , B(19) => muxInB_3_19_port, B(18) => 
                           muxInB_3_18_port, B(17) => muxInB_3_17_port, B(16) 
                           => muxInB_3_16_port, B(15) => muxInB_3_15_port, 
                           B(14) => muxInB_3_14_port, B(13) => muxInB_3_13_port
                           , B(12) => muxInB_3_12_port, B(11) => 
                           muxInB_3_11_port, B(10) => muxInB_3_10_port, B(9) =>
                           muxInB_3_9_port, B(8) => muxInB_3_8_port, B(7) => 
                           muxInB_3_7_port, B(6) => muxInB_3_6_port, B(5) => 
                           net60019, B(4) => net60020, B(3) => net60021, B(2) 
                           => net60022, B(1) => net60023, B(0) => net60024, 
                           C(31) => muxInC_3_31_port, C(30) => muxInC_3_30_port
                           , C(29) => muxInC_3_29_port, C(28) => 
                           muxInC_3_28_port, C(27) => muxInC_3_27_port, C(26) 
                           => muxInC_3_26_port, C(25) => muxInC_3_25_port, 
                           C(24) => muxInC_3_24_port, C(23) => muxInC_3_23_port
                           , C(22) => muxInC_3_22_port, C(21) => 
                           muxInC_3_21_port, C(20) => muxInC_3_20_port, C(19) 
                           => muxInC_3_19_port, C(18) => muxInC_3_18_port, 
                           C(17) => muxInC_3_17_port, C(16) => muxInC_3_16_port
                           , C(15) => muxInC_3_15_port, C(14) => 
                           muxInC_3_14_port, C(13) => muxInC_3_13_port, C(12) 
                           => muxInC_3_12_port, C(11) => muxInC_3_11_port, 
                           C(10) => muxInC_3_10_port, C(9) => muxInC_3_9_port, 
                           C(8) => muxInC_3_8_port, C(7) => muxInC_3_7_port, 
                           C(6) => muxInC_3_6_port, C(5) => net60025, C(4) => 
                           net60026, C(3) => net60027, C(2) => net60028, C(1) 
                           => net60029, C(0) => net60030, D(31) => 
                           muxInD_3_31_port, D(30) => muxInD_3_30_port, D(29) 
                           => muxInD_3_29_port, D(28) => muxInD_3_28_port, 
                           D(27) => muxInD_3_27_port, D(26) => muxInD_3_26_port
                           , D(25) => muxInD_3_25_port, D(24) => 
                           muxInD_3_24_port, D(23) => muxInD_3_23_port, D(22) 
                           => muxInD_3_22_port, D(21) => muxInD_3_21_port, 
                           D(20) => muxInD_3_20_port, D(19) => muxInD_3_19_port
                           , D(18) => muxInD_3_18_port, D(17) => 
                           muxInD_3_17_port, D(16) => muxInD_3_16_port, D(15) 
                           => muxInD_3_15_port, D(14) => muxInD_3_14_port, 
                           D(13) => muxInD_3_13_port, D(12) => muxInD_3_12_port
                           , D(11) => muxInD_3_11_port, D(10) => 
                           muxInD_3_10_port, D(9) => muxInD_3_9_port, D(8) => 
                           muxInD_3_8_port, D(7) => muxInD_3_7_port, D(6) => 
                           net60031, D(5) => net60032, D(4) => net60033, D(3) 
                           => net60034, D(2) => net60035, D(1) => net60036, 
                           D(0) => net60037, E(31) => muxInE_3_31_port, E(30) 
                           => muxInE_3_30_port, E(29) => muxInE_3_29_port, 
                           E(28) => muxInE_3_28_port, E(27) => muxInE_3_27_port
                           , E(26) => muxInE_3_26_port, E(25) => 
                           muxInE_3_25_port, E(24) => muxInE_3_24_port, E(23) 
                           => muxInE_3_23_port, E(22) => muxInE_3_22_port, 
                           E(21) => muxInE_3_21_port, E(20) => muxInE_3_20_port
                           , E(19) => muxInE_3_19_port, E(18) => 
                           muxInE_3_18_port, E(17) => muxInE_3_17_port, E(16) 
                           => muxInE_3_16_port, E(15) => muxInE_3_15_port, 
                           E(14) => muxInE_3_14_port, E(13) => muxInE_3_13_port
                           , E(12) => muxInE_3_12_port, E(11) => 
                           muxInE_3_11_port, E(10) => muxInE_3_10_port, E(9) =>
                           muxInE_3_9_port, E(8) => muxInE_3_8_port, E(7) => 
                           muxInE_3_7_port, E(6) => net60038, E(5) => net60039,
                           E(4) => net60040, E(3) => net60041, E(2) => net60042
                           , E(1) => net60043, E(0) => net60044);
   SHIFTERS_4 : shift_mul_N16_S8 port map( A(15) => n28, A(14) => n27, A(13) =>
                           n26, A(12) => n25, A(11) => n22, A(10) => n21, A(9) 
                           => n19, A(8) => n18, A(7) => n17, A(6) => n15, A(5) 
                           => n14, A(4) => n13, A(3) => n11, A(2) => A(2), A(1)
                           => n10, A(0) => n2, B(31) => muxInB_4_31_port, B(30)
                           => muxInB_4_30_port, B(29) => muxInB_4_29_port, 
                           B(28) => muxInB_4_28_port, B(27) => muxInB_4_27_port
                           , B(26) => muxInB_4_26_port, B(25) => 
                           muxInB_4_25_port, B(24) => muxInB_4_24_port, B(23) 
                           => muxInB_4_23_port, B(22) => muxInB_4_22_port, 
                           B(21) => muxInB_4_21_port, B(20) => muxInB_4_20_port
                           , B(19) => muxInB_4_19_port, B(18) => 
                           muxInB_4_18_port, B(17) => muxInB_4_17_port, B(16) 
                           => muxInB_4_16_port, B(15) => muxInB_4_15_port, 
                           B(14) => muxInB_4_14_port, B(13) => muxInB_4_13_port
                           , B(12) => muxInB_4_12_port, B(11) => 
                           muxInB_4_11_port, B(10) => muxInB_4_10_port, B(9) =>
                           muxInB_4_9_port, B(8) => muxInB_4_8_port, B(7) => 
                           net59985, B(6) => net59986, B(5) => net59987, B(4) 
                           => net59988, B(3) => net59989, B(2) => net59990, 
                           B(1) => net59991, B(0) => net59992, C(31) => 
                           muxInC_4_31_port, C(30) => muxInC_4_30_port, C(29) 
                           => muxInC_4_29_port, C(28) => muxInC_4_28_port, 
                           C(27) => muxInC_4_27_port, C(26) => muxInC_4_26_port
                           , C(25) => muxInC_4_25_port, C(24) => 
                           muxInC_4_24_port, C(23) => muxInC_4_23_port, C(22) 
                           => muxInC_4_22_port, C(21) => muxInC_4_21_port, 
                           C(20) => muxInC_4_20_port, C(19) => muxInC_4_19_port
                           , C(18) => muxInC_4_18_port, C(17) => 
                           muxInC_4_17_port, C(16) => muxInC_4_16_port, C(15) 
                           => muxInC_4_15_port, C(14) => muxInC_4_14_port, 
                           C(13) => muxInC_4_13_port, C(12) => muxInC_4_12_port
                           , C(11) => muxInC_4_11_port, C(10) => 
                           muxInC_4_10_port, C(9) => muxInC_4_9_port, C(8) => 
                           muxInC_4_8_port, C(7) => net59993, C(6) => net59994,
                           C(5) => net59995, C(4) => net59996, C(3) => net59997
                           , C(2) => net59998, C(1) => net59999, C(0) => 
                           net60000, D(31) => muxInD_4_31_port, D(30) => 
                           muxInD_4_30_port, D(29) => muxInD_4_29_port, D(28) 
                           => muxInD_4_28_port, D(27) => muxInD_4_27_port, 
                           D(26) => muxInD_4_26_port, D(25) => muxInD_4_25_port
                           , D(24) => muxInD_4_24_port, D(23) => 
                           muxInD_4_23_port, D(22) => muxInD_4_22_port, D(21) 
                           => muxInD_4_21_port, D(20) => muxInD_4_20_port, 
                           D(19) => muxInD_4_19_port, D(18) => muxInD_4_18_port
                           , D(17) => muxInD_4_17_port, D(16) => 
                           muxInD_4_16_port, D(15) => muxInD_4_15_port, D(14) 
                           => muxInD_4_14_port, D(13) => muxInD_4_13_port, 
                           D(12) => muxInD_4_12_port, D(11) => muxInD_4_11_port
                           , D(10) => muxInD_4_10_port, D(9) => muxInD_4_9_port
                           , D(8) => net60001, D(7) => net60002, D(6) => 
                           net60003, D(5) => net60004, D(4) => net60005, D(3) 
                           => net60006, D(2) => net60007, D(1) => net60008, 
                           D(0) => net60009, E(31) => muxInE_4_31_port, E(30) 
                           => muxInE_4_30_port, E(29) => muxInE_4_29_port, 
                           E(28) => muxInE_4_28_port, E(27) => muxInE_4_27_port
                           , E(26) => muxInE_4_26_port, E(25) => 
                           muxInE_4_25_port, E(24) => muxInE_4_24_port, E(23) 
                           => muxInE_4_23_port, E(22) => muxInE_4_22_port, 
                           E(21) => muxInE_4_21_port, E(20) => muxInE_4_20_port
                           , E(19) => muxInE_4_19_port, E(18) => 
                           muxInE_4_18_port, E(17) => muxInE_4_17_port, E(16) 
                           => muxInE_4_16_port, E(15) => muxInE_4_15_port, 
                           E(14) => muxInE_4_14_port, E(13) => muxInE_4_13_port
                           , E(12) => muxInE_4_12_port, E(11) => 
                           muxInE_4_11_port, E(10) => muxInE_4_10_port, E(9) =>
                           muxInE_4_9_port, E(8) => net60010, E(7) => net60011,
                           E(6) => net60012, E(5) => net60013, E(4) => net60014
                           , E(3) => net60015, E(2) => net60016, E(1) => 
                           net60017, E(0) => net60018);
   SHIFTERS_5 : shift_mul_N16_S10 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n3, B(31) => muxInB_5_31_port, 
                           B(30) => muxInB_5_30_port, B(29) => muxInB_5_29_port
                           , B(28) => muxInB_5_28_port, B(27) => 
                           muxInB_5_27_port, B(26) => muxInB_5_26_port, B(25) 
                           => muxInB_5_25_port, B(24) => muxInB_5_24_port, 
                           B(23) => muxInB_5_23_port, B(22) => muxInB_5_22_port
                           , B(21) => muxInB_5_21_port, B(20) => 
                           muxInB_5_20_port, B(19) => muxInB_5_19_port, B(18) 
                           => muxInB_5_18_port, B(17) => muxInB_5_17_port, 
                           B(16) => muxInB_5_16_port, B(15) => muxInB_5_15_port
                           , B(14) => muxInB_5_14_port, B(13) => 
                           muxInB_5_13_port, B(12) => muxInB_5_12_port, B(11) 
                           => muxInB_5_11_port, B(10) => muxInB_5_10_port, B(9)
                           => net59943, B(8) => net59944, B(7) => net59945, 
                           B(6) => net59946, B(5) => net59947, B(4) => net59948
                           , B(3) => net59949, B(2) => net59950, B(1) => 
                           net59951, B(0) => net59952, C(31) => 
                           muxInC_5_31_port, C(30) => muxInC_5_30_port, C(29) 
                           => muxInC_5_29_port, C(28) => muxInC_5_28_port, 
                           C(27) => muxInC_5_27_port, C(26) => muxInC_5_26_port
                           , C(25) => muxInC_5_25_port, C(24) => 
                           muxInC_5_24_port, C(23) => muxInC_5_23_port, C(22) 
                           => muxInC_5_22_port, C(21) => muxInC_5_21_port, 
                           C(20) => muxInC_5_20_port, C(19) => muxInC_5_19_port
                           , C(18) => muxInC_5_18_port, C(17) => 
                           muxInC_5_17_port, C(16) => muxInC_5_16_port, C(15) 
                           => muxInC_5_15_port, C(14) => muxInC_5_14_port, 
                           C(13) => muxInC_5_13_port, C(12) => muxInC_5_12_port
                           , C(11) => muxInC_5_11_port, C(10) => 
                           muxInC_5_10_port, C(9) => net59953, C(8) => net59954
                           , C(7) => net59955, C(6) => net59956, C(5) => 
                           net59957, C(4) => net59958, C(3) => net59959, C(2) 
                           => net59960, C(1) => net59961, C(0) => net59962, 
                           D(31) => muxInD_5_31_port, D(30) => muxInD_5_30_port
                           , D(29) => muxInD_5_29_port, D(28) => 
                           muxInD_5_28_port, D(27) => muxInD_5_27_port, D(26) 
                           => muxInD_5_26_port, D(25) => muxInD_5_25_port, 
                           D(24) => muxInD_5_24_port, D(23) => muxInD_5_23_port
                           , D(22) => muxInD_5_22_port, D(21) => 
                           muxInD_5_21_port, D(20) => muxInD_5_20_port, D(19) 
                           => muxInD_5_19_port, D(18) => muxInD_5_18_port, 
                           D(17) => muxInD_5_17_port, D(16) => muxInD_5_16_port
                           , D(15) => muxInD_5_15_port, D(14) => 
                           muxInD_5_14_port, D(13) => muxInD_5_13_port, D(12) 
                           => muxInD_5_12_port, D(11) => muxInD_5_11_port, 
                           D(10) => net59963, D(9) => net59964, D(8) => 
                           net59965, D(7) => net59966, D(6) => net59967, D(5) 
                           => net59968, D(4) => net59969, D(3) => net59970, 
                           D(2) => net59971, D(1) => net59972, D(0) => net59973
                           , E(31) => muxInE_5_31_port, E(30) => 
                           muxInE_5_30_port, E(29) => muxInE_5_29_port, E(28) 
                           => muxInE_5_28_port, E(27) => muxInE_5_27_port, 
                           E(26) => muxInE_5_26_port, E(25) => muxInE_5_25_port
                           , E(24) => muxInE_5_24_port, E(23) => 
                           muxInE_5_23_port, E(22) => muxInE_5_22_port, E(21) 
                           => muxInE_5_21_port, E(20) => muxInE_5_20_port, 
                           E(19) => muxInE_5_19_port, E(18) => muxInE_5_18_port
                           , E(17) => muxInE_5_17_port, E(16) => 
                           muxInE_5_16_port, E(15) => muxInE_5_15_port, E(14) 
                           => muxInE_5_14_port, E(13) => muxInE_5_13_port, 
                           E(12) => muxInE_5_12_port, E(11) => muxInE_5_11_port
                           , E(10) => net59974, E(9) => net59975, E(8) => 
                           net59976, E(7) => net59977, E(6) => net59978, E(5) 
                           => net59979, E(4) => net59980, E(3) => net59981, 
                           E(2) => net59982, E(1) => net59983, E(0) => net59984
                           );
   SHIFTERS_6 : shift_mul_N16_S12 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n3, B(31) => muxInB_6_31_port, 
                           B(30) => muxInB_6_30_port, B(29) => muxInB_6_29_port
                           , B(28) => muxInB_6_28_port, B(27) => 
                           muxInB_6_27_port, B(26) => muxInB_6_26_port, B(25) 
                           => muxInB_6_25_port, B(24) => muxInB_6_24_port, 
                           B(23) => muxInB_6_23_port, B(22) => muxInB_6_22_port
                           , B(21) => muxInB_6_21_port, B(20) => 
                           muxInB_6_20_port, B(19) => muxInB_6_19_port, B(18) 
                           => muxInB_6_18_port, B(17) => muxInB_6_17_port, 
                           B(16) => muxInB_6_16_port, B(15) => muxInB_6_15_port
                           , B(14) => muxInB_6_14_port, B(13) => 
                           muxInB_6_13_port, B(12) => muxInB_6_12_port, B(11) 
                           => net59893, B(10) => net59894, B(9) => net59895, 
                           B(8) => net59896, B(7) => net59897, B(6) => net59898
                           , B(5) => net59899, B(4) => net59900, B(3) => 
                           net59901, B(2) => net59902, B(1) => net59903, B(0) 
                           => net59904, C(31) => muxInC_6_31_port, C(30) => 
                           muxInC_6_30_port, C(29) => muxInC_6_29_port, C(28) 
                           => muxInC_6_28_port, C(27) => muxInC_6_27_port, 
                           C(26) => muxInC_6_26_port, C(25) => muxInC_6_25_port
                           , C(24) => muxInC_6_24_port, C(23) => 
                           muxInC_6_23_port, C(22) => muxInC_6_22_port, C(21) 
                           => muxInC_6_21_port, C(20) => muxInC_6_20_port, 
                           C(19) => muxInC_6_19_port, C(18) => muxInC_6_18_port
                           , C(17) => muxInC_6_17_port, C(16) => 
                           muxInC_6_16_port, C(15) => muxInC_6_15_port, C(14) 
                           => muxInC_6_14_port, C(13) => muxInC_6_13_port, 
                           C(12) => muxInC_6_12_port, C(11) => net59905, C(10) 
                           => net59906, C(9) => net59907, C(8) => net59908, 
                           C(7) => net59909, C(6) => net59910, C(5) => net59911
                           , C(4) => net59912, C(3) => net59913, C(2) => 
                           net59914, C(1) => net59915, C(0) => net59916, D(31) 
                           => muxInD_6_31_port, D(30) => muxInD_6_30_port, 
                           D(29) => muxInD_6_29_port, D(28) => muxInD_6_28_port
                           , D(27) => muxInD_6_27_port, D(26) => 
                           muxInD_6_26_port, D(25) => muxInD_6_25_port, D(24) 
                           => muxInD_6_24_port, D(23) => muxInD_6_23_port, 
                           D(22) => muxInD_6_22_port, D(21) => muxInD_6_21_port
                           , D(20) => muxInD_6_20_port, D(19) => 
                           muxInD_6_19_port, D(18) => muxInD_6_18_port, D(17) 
                           => muxInD_6_17_port, D(16) => muxInD_6_16_port, 
                           D(15) => muxInD_6_15_port, D(14) => muxInD_6_14_port
                           , D(13) => muxInD_6_13_port, D(12) => net59917, 
                           D(11) => net59918, D(10) => net59919, D(9) => 
                           net59920, D(8) => net59921, D(7) => net59922, D(6) 
                           => net59923, D(5) => net59924, D(4) => net59925, 
                           D(3) => net59926, D(2) => net59927, D(1) => net59928
                           , D(0) => net59929, E(31) => muxInE_6_31_port, E(30)
                           => muxInE_6_30_port, E(29) => muxInE_6_29_port, 
                           E(28) => muxInE_6_28_port, E(27) => muxInE_6_27_port
                           , E(26) => muxInE_6_26_port, E(25) => 
                           muxInE_6_25_port, E(24) => muxInE_6_24_port, E(23) 
                           => muxInE_6_23_port, E(22) => muxInE_6_22_port, 
                           E(21) => muxInE_6_21_port, E(20) => muxInE_6_20_port
                           , E(19) => muxInE_6_19_port, E(18) => 
                           muxInE_6_18_port, E(17) => muxInE_6_17_port, E(16) 
                           => muxInE_6_16_port, E(15) => muxInE_6_15_port, 
                           E(14) => muxInE_6_14_port, E(13) => muxInE_6_13_port
                           , E(12) => net59930, E(11) => net59931, E(10) => 
                           net59932, E(9) => net59933, E(8) => net59934, E(7) 
                           => net59935, E(6) => net59936, E(5) => net59937, 
                           E(4) => net59938, E(3) => net59939, E(2) => net59940
                           , E(1) => net59941, E(0) => net59942);
   SHIFTERS_7 : shift_mul_N16_S14 port map( A(15) => n28, A(14) => n27, A(13) 
                           => n26, A(12) => n25, A(11) => n22, A(10) => n21, 
                           A(9) => n19, A(8) => n18, A(7) => n17, A(6) => n15, 
                           A(5) => n14, A(4) => n13, A(3) => n11, A(2) => A(2),
                           A(1) => n10, A(0) => n2, B(31) => muxInB_7_31_port, 
                           B(30) => muxInB_7_30_port, B(29) => muxInB_7_29_port
                           , B(28) => muxInB_7_28_port, B(27) => 
                           muxInB_7_27_port, B(26) => muxInB_7_26_port, B(25) 
                           => muxInB_7_25_port, B(24) => muxInB_7_24_port, 
                           B(23) => muxInB_7_23_port, B(22) => muxInB_7_22_port
                           , B(21) => muxInB_7_21_port, B(20) => 
                           muxInB_7_20_port, B(19) => muxInB_7_19_port, B(18) 
                           => muxInB_7_18_port, B(17) => muxInB_7_17_port, 
                           B(16) => muxInB_7_16_port, B(15) => muxInB_7_15_port
                           , B(14) => muxInB_7_14_port, B(13) => net59835, 
                           B(12) => net59836, B(11) => net59837, B(10) => 
                           net59838, B(9) => net59839, B(8) => net59840, B(7) 
                           => net59841, B(6) => net59842, B(5) => net59843, 
                           B(4) => net59844, B(3) => net59845, B(2) => net59846
                           , B(1) => net59847, B(0) => net59848, C(31) => 
                           muxInC_7_31_port, C(30) => muxInC_7_30_port, C(29) 
                           => muxInC_7_29_port, C(28) => muxInC_7_28_port, 
                           C(27) => muxInC_7_27_port, C(26) => muxInC_7_26_port
                           , C(25) => muxInC_7_25_port, C(24) => 
                           muxInC_7_24_port, C(23) => muxInC_7_23_port, C(22) 
                           => muxInC_7_22_port, C(21) => muxInC_7_21_port, 
                           C(20) => muxInC_7_20_port, C(19) => muxInC_7_19_port
                           , C(18) => muxInC_7_18_port, C(17) => 
                           muxInC_7_17_port, C(16) => muxInC_7_16_port, C(15) 
                           => muxInC_7_15_port, C(14) => muxInC_7_14_port, 
                           C(13) => net59849, C(12) => net59850, C(11) => 
                           net59851, C(10) => net59852, C(9) => net59853, C(8) 
                           => net59854, C(7) => net59855, C(6) => net59856, 
                           C(5) => net59857, C(4) => net59858, C(3) => net59859
                           , C(2) => net59860, C(1) => net59861, C(0) => 
                           net59862, D(31) => muxInD_7_31_port, D(30) => 
                           muxInD_7_30_port, D(29) => muxInD_7_29_port, D(28) 
                           => muxInD_7_28_port, D(27) => muxInD_7_27_port, 
                           D(26) => muxInD_7_26_port, D(25) => muxInD_7_25_port
                           , D(24) => muxInD_7_24_port, D(23) => 
                           muxInD_7_23_port, D(22) => muxInD_7_22_port, D(21) 
                           => muxInD_7_21_port, D(20) => muxInD_7_20_port, 
                           D(19) => muxInD_7_19_port, D(18) => muxInD_7_18_port
                           , D(17) => muxInD_7_17_port, D(16) => 
                           muxInD_7_16_port, D(15) => muxInD_7_15_port, D(14) 
                           => net59863, D(13) => net59864, D(12) => net59865, 
                           D(11) => net59866, D(10) => net59867, D(9) => 
                           net59868, D(8) => net59869, D(7) => net59870, D(6) 
                           => net59871, D(5) => net59872, D(4) => net59873, 
                           D(3) => net59874, D(2) => net59875, D(1) => net59876
                           , D(0) => net59877, E(31) => muxInE_7_31_port, E(30)
                           => muxInE_7_30_port, E(29) => muxInE_7_29_port, 
                           E(28) => muxInE_7_28_port, E(27) => muxInE_7_27_port
                           , E(26) => muxInE_7_26_port, E(25) => 
                           muxInE_7_25_port, E(24) => muxInE_7_24_port, E(23) 
                           => muxInE_7_23_port, E(22) => muxInE_7_22_port, 
                           E(21) => muxInE_7_21_port, E(20) => muxInE_7_20_port
                           , E(19) => muxInE_7_19_port, E(18) => 
                           muxInE_7_18_port, E(17) => muxInE_7_17_port, E(16) 
                           => muxInE_7_16_port, E(15) => muxInE_7_15_port, 
                           E(14) => net59878, E(13) => net59879, E(12) => 
                           net59880, E(11) => net59881, E(10) => net59882, E(9)
                           => net59883, E(8) => net59884, E(7) => net59885, 
                           E(6) => net59886, E(5) => net59887, E(4) => net59888
                           , E(3) => net59889, E(2) => net59890, E(1) => 
                           net59891, E(0) => net59892);
   MUXGEN_0 : mux_N32_0 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_0_31_port, B(30) => 
                           muxInB_0_30_port, B(29) => muxInB_0_29_port, B(28) 
                           => muxInB_0_28_port, B(27) => muxInB_0_27_port, 
                           B(26) => muxInB_0_26_port, B(25) => muxInB_0_25_port
                           , B(24) => muxInB_0_24_port, B(23) => 
                           muxInB_0_23_port, B(22) => muxInB_0_22_port, B(21) 
                           => muxInB_0_21_port, B(20) => muxInB_0_20_port, 
                           B(19) => muxInB_0_19_port, B(18) => muxInB_0_18_port
                           , B(17) => muxInB_0_17_port, B(16) => 
                           muxInB_0_16_port, B(15) => muxInB_0_15_port, B(14) 
                           => muxInB_0_14_port, B(13) => muxInB_0_13_port, 
                           B(12) => muxInB_0_12_port, B(11) => muxInB_0_11_port
                           , B(10) => muxInB_0_10_port, B(9) => muxInB_0_9_port
                           , B(8) => muxInB_0_8_port, B(7) => muxInB_0_7_port, 
                           B(6) => muxInB_0_6_port, B(5) => muxInB_0_5_port, 
                           B(4) => muxInB_0_4_port, B(3) => muxInB_0_3_port, 
                           B(2) => muxInB_0_2_port, B(1) => muxInB_0_1_port, 
                           B(0) => muxInB_0_0_port, C(31) => muxInC_0_31_port, 
                           C(30) => muxInC_0_30_port, C(29) => muxInC_0_29_port
                           , C(28) => muxInC_0_28_port, C(27) => 
                           muxInC_0_20_port, C(26) => muxInC_0_26_port, C(25) 
                           => muxInC_0_25_port, C(24) => muxInC_0_24_port, 
                           C(23) => muxInC_0_23_port, C(22) => muxInC_0_22_port
                           , C(21) => muxInC_0_21_port, C(20) => 
                           muxInC_0_20_port, C(19) => muxInC_0_19_port, C(18) 
                           => muxInC_0_18_port, C(17) => muxInC_0_17_port, 
                           C(16) => muxInC_0_16_port, C(15) => muxInC_0_15_port
                           , C(14) => muxInC_0_14_port, C(13) => 
                           muxInC_0_13_port, C(12) => muxInC_0_12_port, C(11) 
                           => muxInC_0_11_port, C(10) => muxInC_0_10_port, C(9)
                           => muxInC_0_9_port, C(8) => muxInC_0_8_port, C(7) =>
                           muxInC_0_7_port, C(6) => muxInC_0_6_port, C(5) => 
                           muxInC_0_5_port, C(4) => muxInC_0_4_port, C(3) => 
                           muxInC_0_3_port, C(2) => muxInC_0_2_port, C(1) => 
                           muxInC_0_1_port, C(0) => muxInC_0_0_port, D(31) => 
                           muxInD_0_31_port, D(30) => muxInD_0_30_port, D(29) 
                           => muxInD_0_29_port, D(28) => muxInD_0_28_port, 
                           D(27) => muxInD_0_27_port, D(26) => muxInD_0_26_port
                           , D(25) => muxInD_0_25_port, D(24) => 
                           muxInD_0_24_port, D(23) => muxInD_0_23_port, D(22) 
                           => muxInD_0_22_port, D(21) => muxInD_0_21_port, 
                           D(20) => muxInD_0_20_port, D(19) => muxInD_0_19_port
                           , D(18) => muxInD_0_18_port, D(17) => 
                           muxInD_0_17_port, D(16) => muxInD_0_16_port, D(15) 
                           => muxInD_0_15_port, D(14) => muxInD_0_14_port, 
                           D(13) => muxInD_0_13_port, D(12) => muxInD_0_12_port
                           , D(11) => muxInD_0_11_port, D(10) => 
                           muxInD_0_10_port, D(9) => muxInD_0_9_port, D(8) => 
                           muxInD_0_8_port, D(7) => muxInD_0_7_port, D(6) => 
                           muxInD_0_6_port, D(5) => muxInD_0_5_port, D(4) => 
                           muxInD_0_4_port, D(3) => muxInD_0_3_port, D(2) => 
                           muxInD_0_2_port, D(1) => muxInD_0_1_port, D(0) => 
                           muxInD_0_0_port, E(31) => muxInE_0_31_port, E(30) =>
                           muxInE_0_30_port, E(29) => muxInE_0_29_port, E(28) 
                           => muxInE_0_28_port, E(27) => muxInE_0_27_port, 
                           E(26) => muxInE_0_26_port, E(25) => muxInC_0_20_port
                           , E(24) => muxInE_0_24_port, E(23) => 
                           muxInE_0_23_port, E(22) => muxInC_0_27_port, E(21) 
                           => muxInE_0_21_port, E(20) => muxInE_0_20_port, 
                           E(19) => muxInE_0_19_port, E(18) => muxInE_0_18_port
                           , E(17) => muxInC_0_29_port, E(16) => 
                           muxInE_0_16_port, E(15) => muxInE_0_15_port, E(14) 
                           => muxInE_0_14_port, E(13) => muxInE_0_13_port, 
                           E(12) => muxInE_0_12_port, E(11) => muxInE_0_11_port
                           , E(10) => muxInE_0_10_port, E(9) => muxInE_0_9_port
                           , E(8) => muxInE_0_8_port, E(7) => muxInE_0_7_port, 
                           E(6) => muxInE_0_6_port, E(5) => muxInE_0_5_port, 
                           E(4) => muxInE_0_4_port, E(3) => muxInE_0_3_port, 
                           E(2) => muxInE_0_2_port, E(1) => muxInE_0_1_port, 
                           E(0) => muxInE_0_0_port, Sel(2) => B(1), Sel(1) => 
                           B(0), Sel(0) => X_Logic0_port, O(31) => 
                           outmux_0_31_port, O(30) => outmux_0_30_port, O(29) 
                           => outmux_0_29_port, O(28) => outmux_0_28_port, 
                           O(27) => outmux_0_27_port, O(26) => outmux_0_26_port
                           , O(25) => outmux_0_25_port, O(24) => 
                           outmux_0_24_port, O(23) => outmux_0_23_port, O(22) 
                           => outmux_0_22_port, O(21) => outmux_0_21_port, 
                           O(20) => outmux_0_20_port, O(19) => outmux_0_19_port
                           , O(18) => outmux_0_18_port, O(17) => 
                           outmux_0_17_port, O(16) => outmux_0_16_port, O(15) 
                           => outmux_0_15_port, O(14) => outmux_0_14_port, 
                           O(13) => outmux_0_13_port, O(12) => outmux_0_12_port
                           , O(11) => outmux_0_11_port, O(10) => 
                           outmux_0_10_port, O(9) => outmux_0_9_port, O(8) => 
                           outmux_0_8_port, O(7) => outmux_0_7_port, O(6) => 
                           outmux_0_6_port, O(5) => outmux_0_5_port, O(4) => 
                           outmux_0_4_port, O(3) => outmux_0_3_port, O(2) => 
                           outmux_0_2_port, O(1) => outmux_0_1_port, O(0) => 
                           outmux_0_0_port);
   MUXGEN_1 : mux_N32_7 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_1_31_port, B(30) => 
                           muxInB_1_30_port, B(29) => muxInB_1_29_port, B(28) 
                           => muxInB_1_28_port, B(27) => muxInB_1_27_port, 
                           B(26) => muxInB_1_26_port, B(25) => muxInB_1_25_port
                           , B(24) => muxInB_1_24_port, B(23) => 
                           muxInB_1_23_port, B(22) => muxInB_1_22_port, B(21) 
                           => muxInB_1_21_port, B(20) => muxInB_1_20_port, 
                           B(19) => muxInB_1_19_port, B(18) => muxInB_1_18_port
                           , B(17) => muxInB_1_17_port, B(16) => 
                           muxInB_1_16_port, B(15) => muxInB_1_15_port, B(14) 
                           => muxInB_1_14_port, B(13) => muxInB_1_13_port, 
                           B(12) => muxInB_1_12_port, B(11) => muxInB_1_11_port
                           , B(10) => muxInB_1_10_port, B(9) => muxInB_1_9_port
                           , B(8) => muxInB_1_8_port, B(7) => muxInB_1_7_port, 
                           B(6) => muxInB_1_6_port, B(5) => muxInB_1_5_port, 
                           B(4) => muxInB_1_4_port, B(3) => muxInB_1_3_port, 
                           B(2) => muxInB_1_2_port, B(1) => muxInB_1_1_port, 
                           B(0) => muxInB_1_0_port, C(31) => muxInC_1_31_port, 
                           C(30) => muxInC_1_30_port, C(29) => muxInC_1_29_port
                           , C(28) => muxInC_1_28_port, C(27) => 
                           muxInC_1_27_port, C(26) => muxInC_1_26_port, C(25) 
                           => muxInC_1_25_port, C(24) => muxInC_1_24_port, 
                           C(23) => muxInE_1_23_port, C(22) => muxInC_1_22_port
                           , C(21) => muxInC_1_21_port, C(20) => 
                           muxInC_1_20_port, C(19) => muxInC_1_23_port, C(18) 
                           => muxInC_1_18_port, C(17) => muxInC_1_17_port, 
                           C(16) => muxInC_1_16_port, C(15) => muxInC_1_15_port
                           , C(14) => muxInC_1_14_port, C(13) => 
                           muxInC_1_13_port, C(12) => muxInC_1_12_port, C(11) 
                           => muxInC_1_11_port, C(10) => muxInC_1_10_port, C(9)
                           => muxInC_1_9_port, C(8) => muxInC_1_8_port, C(7) =>
                           muxInC_1_7_port, C(6) => muxInC_1_6_port, C(5) => 
                           muxInC_1_5_port, C(4) => muxInC_1_4_port, C(3) => 
                           muxInC_1_3_port, C(2) => muxInC_1_2_port, C(1) => 
                           muxInC_1_1_port, C(0) => muxInC_1_0_port, D(31) => 
                           muxInD_1_31_port, D(30) => muxInD_1_30_port, D(29) 
                           => muxInD_1_29_port, D(28) => muxInD_1_28_port, 
                           D(27) => muxInD_1_27_port, D(26) => muxInD_1_26_port
                           , D(25) => muxInD_1_25_port, D(24) => 
                           muxInD_1_24_port, D(23) => muxInD_1_23_port, D(22) 
                           => muxInD_1_22_port, D(21) => muxInD_1_21_port, 
                           D(20) => muxInD_1_20_port, D(19) => muxInD_1_19_port
                           , D(18) => muxInD_1_18_port, D(17) => 
                           muxInD_1_17_port, D(16) => muxInD_1_16_port, D(15) 
                           => muxInD_1_15_port, D(14) => muxInD_1_14_port, 
                           D(13) => muxInD_1_13_port, D(12) => muxInD_1_12_port
                           , D(11) => muxInD_1_11_port, D(10) => 
                           muxInD_1_10_port, D(9) => muxInD_1_9_port, D(8) => 
                           muxInD_1_8_port, D(7) => muxInD_1_7_port, D(6) => 
                           muxInD_1_6_port, D(5) => muxInD_1_5_port, D(4) => 
                           muxInD_1_4_port, D(3) => muxInD_1_3_port, D(2) => 
                           muxInD_1_2_port, D(1) => muxInD_1_1_port, D(0) => 
                           muxInD_1_0_port, E(31) => muxInE_1_31_port, E(30) =>
                           muxInE_1_30_port, E(29) => muxInE_1_29_port, E(28) 
                           => muxInE_1_28_port, E(27) => muxInE_1_27_port, 
                           E(26) => muxInE_1_26_port, E(25) => muxInE_1_25_port
                           , E(24) => muxInE_1_24_port, E(23) => 
                           muxInE_1_23_port, E(22) => muxInE_1_22_port, E(21) 
                           => muxInE_1_21_port, E(20) => muxInE_1_20_port, 
                           E(19) => muxInE_1_19_port, E(18) => muxInE_1_18_port
                           , E(17) => muxInE_1_17_port, E(16) => 
                           muxInE_1_16_port, E(15) => muxInE_1_15_port, E(14) 
                           => muxInE_1_14_port, E(13) => muxInE_1_13_port, 
                           E(12) => muxInE_1_12_port, E(11) => muxInE_1_11_port
                           , E(10) => muxInE_1_10_port, E(9) => muxInE_1_9_port
                           , E(8) => muxInE_1_8_port, E(7) => muxInE_1_7_port, 
                           E(6) => muxInE_1_6_port, E(5) => muxInE_1_5_port, 
                           E(4) => muxInE_1_4_port, E(3) => muxInE_1_3_port, 
                           E(2) => muxInE_1_2_port, E(1) => muxInE_1_1_port, 
                           E(0) => muxInE_1_0_port, Sel(2) => B(3), Sel(1) => 
                           B(2), Sel(0) => B(1), O(31) => outmux_1_31_port, 
                           O(30) => outmux_1_30_port, O(29) => outmux_1_29_port
                           , O(28) => outmux_1_28_port, O(27) => 
                           outmux_1_27_port, O(26) => outmux_1_26_port, O(25) 
                           => outmux_1_25_port, O(24) => outmux_1_24_port, 
                           O(23) => outmux_1_23_port, O(22) => outmux_1_22_port
                           , O(21) => outmux_1_21_port, O(20) => 
                           outmux_1_20_port, O(19) => outmux_1_19_port, O(18) 
                           => outmux_1_18_port, O(17) => outmux_1_17_port, 
                           O(16) => outmux_1_16_port, O(15) => outmux_1_15_port
                           , O(14) => outmux_1_14_port, O(13) => 
                           outmux_1_13_port, O(12) => outmux_1_12_port, O(11) 
                           => outmux_1_11_port, O(10) => outmux_1_10_port, O(9)
                           => outmux_1_9_port, O(8) => outmux_1_8_port, O(7) =>
                           outmux_1_7_port, O(6) => outmux_1_6_port, O(5) => 
                           outmux_1_5_port, O(4) => outmux_1_4_port, O(3) => 
                           outmux_1_3_port, O(2) => outmux_1_2_port, O(1) => 
                           outmux_1_1_port, O(0) => outmux_1_0_port);
   MUXGEN_2 : mux_N32_6 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_2_31_port, B(30) => 
                           muxInB_2_30_port, B(29) => muxInB_2_29_port, B(28) 
                           => muxInB_2_28_port, B(27) => muxInB_2_27_port, 
                           B(26) => muxInB_2_26_port, B(25) => muxInB_2_25_port
                           , B(24) => muxInB_2_24_port, B(23) => 
                           muxInB_2_23_port, B(22) => muxInB_2_22_port, B(21) 
                           => muxInB_2_21_port, B(20) => muxInB_2_20_port, 
                           B(19) => muxInB_2_19_port, B(18) => muxInB_2_18_port
                           , B(17) => muxInB_2_17_port, B(16) => 
                           muxInB_2_16_port, B(15) => muxInB_2_15_port, B(14) 
                           => muxInB_2_14_port, B(13) => muxInB_2_13_port, 
                           B(12) => muxInB_2_12_port, B(11) => muxInB_2_11_port
                           , B(10) => muxInB_2_10_port, B(9) => muxInB_2_9_port
                           , B(8) => muxInB_2_8_port, B(7) => muxInB_2_7_port, 
                           B(6) => muxInB_2_6_port, B(5) => muxInB_2_5_port, 
                           B(4) => muxInB_2_4_port, B(3) => muxInB_2_3_port, 
                           B(2) => muxInB_2_2_port, B(1) => muxInB_2_1_port, 
                           B(0) => muxInB_2_0_port, C(31) => muxInC_2_31_port, 
                           C(30) => muxInC_2_30_port, C(29) => muxInC_2_29_port
                           , C(28) => muxInC_2_28_port, C(27) => 
                           muxInC_2_27_port, C(26) => muxInC_2_26_port, C(25) 
                           => muxInC_2_25_port, C(24) => muxInC_2_24_port, 
                           C(23) => muxInC_2_23_port, C(22) => muxInC_2_22_port
                           , C(21) => muxInC_2_21_port, C(20) => 
                           muxInC_2_20_port, C(19) => n20, C(18) => 
                           muxInC_2_18_port, C(17) => muxInC_2_17_port, C(16) 
                           => muxInC_2_16_port, C(15) => muxInC_2_15_port, 
                           C(14) => muxInC_2_14_port, C(13) => muxInC_2_13_port
                           , C(12) => muxInC_2_12_port, C(11) => 
                           muxInC_2_11_port, C(10) => muxInC_2_10_port, C(9) =>
                           muxInC_2_9_port, C(8) => muxInC_2_8_port, C(7) => 
                           muxInC_2_7_port, C(6) => muxInC_2_6_port, C(5) => 
                           muxInC_2_5_port, C(4) => muxInC_2_4_port, C(3) => 
                           muxInC_2_3_port, C(2) => muxInC_2_2_port, C(1) => 
                           muxInC_2_1_port, C(0) => muxInC_2_0_port, D(31) => 
                           muxInD_2_31_port, D(30) => muxInD_2_30_port, D(29) 
                           => muxInD_2_29_port, D(28) => muxInD_2_28_port, 
                           D(27) => muxInD_2_27_port, D(26) => muxInD_2_26_port
                           , D(25) => muxInD_2_25_port, D(24) => 
                           muxInD_2_24_port, D(23) => muxInD_2_23_port, D(22) 
                           => muxInD_2_22_port, D(21) => muxInD_2_21_port, 
                           D(20) => muxInD_2_20_port, D(19) => muxInD_2_19_port
                           , D(18) => muxInD_2_18_port, D(17) => 
                           muxInD_2_17_port, D(16) => muxInD_2_16_port, D(15) 
                           => muxInD_2_15_port, D(14) => muxInD_2_14_port, 
                           D(13) => muxInD_2_13_port, D(12) => muxInD_2_12_port
                           , D(11) => muxInD_2_11_port, D(10) => 
                           muxInD_2_10_port, D(9) => muxInD_2_9_port, D(8) => 
                           muxInD_2_8_port, D(7) => muxInD_2_7_port, D(6) => 
                           muxInD_2_6_port, D(5) => muxInD_2_5_port, D(4) => 
                           muxInD_2_4_port, D(3) => muxInD_2_3_port, D(2) => 
                           muxInD_2_2_port, D(1) => muxInD_2_1_port, D(0) => 
                           muxInD_2_0_port, E(31) => muxInE_2_31_port, E(30) =>
                           muxInE_2_30_port, E(29) => muxInE_2_29_port, E(28) 
                           => muxInE_2_28_port, E(27) => muxInE_2_27_port, 
                           E(26) => muxInE_2_26_port, E(25) => muxInE_2_25_port
                           , E(24) => muxInE_2_24_port, E(23) => 
                           muxInE_2_23_port, E(22) => muxInE_2_22_port, E(21) 
                           => muxInE_2_21_port, E(20) => muxInC_2_19_port, 
                           E(19) => muxInE_2_19_port, E(18) => muxInE_2_18_port
                           , E(17) => muxInE_2_17_port, E(16) => 
                           muxInE_2_16_port, E(15) => muxInE_2_15_port, E(14) 
                           => muxInE_2_14_port, E(13) => muxInE_2_13_port, 
                           E(12) => muxInE_2_12_port, E(11) => muxInE_2_11_port
                           , E(10) => muxInE_2_10_port, E(9) => muxInE_2_9_port
                           , E(8) => muxInE_2_8_port, E(7) => muxInE_2_7_port, 
                           E(6) => muxInE_2_6_port, E(5) => muxInE_2_5_port, 
                           E(4) => muxInE_2_4_port, E(3) => muxInE_2_3_port, 
                           E(2) => muxInE_2_2_port, E(1) => muxInE_2_1_port, 
                           E(0) => muxInE_2_0_port, Sel(2) => B(5), Sel(1) => 
                           B(4), Sel(0) => B(3), O(31) => outmux_2_31_port, 
                           O(30) => outmux_2_30_port, O(29) => outmux_2_29_port
                           , O(28) => outmux_2_28_port, O(27) => 
                           outmux_2_27_port, O(26) => outmux_2_26_port, O(25) 
                           => outmux_2_25_port, O(24) => outmux_2_24_port, 
                           O(23) => outmux_2_23_port, O(22) => outmux_2_22_port
                           , O(21) => outmux_2_21_port, O(20) => 
                           outmux_2_20_port, O(19) => outmux_2_19_port, O(18) 
                           => outmux_2_18_port, O(17) => outmux_2_17_port, 
                           O(16) => outmux_2_16_port, O(15) => outmux_2_15_port
                           , O(14) => outmux_2_14_port, O(13) => 
                           outmux_2_13_port, O(12) => outmux_2_12_port, O(11) 
                           => outmux_2_11_port, O(10) => outmux_2_10_port, O(9)
                           => outmux_2_9_port, O(8) => outmux_2_8_port, O(7) =>
                           outmux_2_7_port, O(6) => outmux_2_6_port, O(5) => 
                           outmux_2_5_port, O(4) => outmux_2_4_port, O(3) => 
                           outmux_2_3_port, O(2) => outmux_2_2_port, O(1) => 
                           outmux_2_1_port, O(0) => outmux_2_0_port);
   MUXGEN_3 : mux_N32_5 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_3_31_port, B(30) => 
                           muxInB_3_30_port, B(29) => muxInB_3_29_port, B(28) 
                           => muxInB_3_28_port, B(27) => muxInB_3_27_port, 
                           B(26) => muxInB_3_26_port, B(25) => muxInB_3_25_port
                           , B(24) => muxInB_3_24_port, B(23) => 
                           muxInB_3_23_port, B(22) => muxInB_3_22_port, B(21) 
                           => muxInB_3_21_port, B(20) => muxInB_3_20_port, 
                           B(19) => muxInB_3_19_port, B(18) => muxInB_3_18_port
                           , B(17) => muxInB_3_17_port, B(16) => 
                           muxInB_3_16_port, B(15) => muxInB_3_15_port, B(14) 
                           => muxInB_3_14_port, B(13) => muxInB_3_13_port, 
                           B(12) => muxInB_3_12_port, B(11) => muxInB_3_11_port
                           , B(10) => muxInB_3_10_port, B(9) => muxInB_3_9_port
                           , B(8) => muxInB_3_8_port, B(7) => muxInB_3_7_port, 
                           B(6) => muxInB_3_6_port, B(5) => muxInB_3_5_port, 
                           B(4) => muxInB_3_4_port, B(3) => muxInB_3_3_port, 
                           B(2) => muxInB_3_2_port, B(1) => muxInB_3_1_port, 
                           B(0) => muxInB_3_0_port, C(31) => muxInC_3_31_port, 
                           C(30) => muxInC_3_30_port, C(29) => muxInC_3_29_port
                           , C(28) => muxInC_3_28_port, C(27) => 
                           muxInC_3_27_port, C(26) => muxInC_3_26_port, C(25) 
                           => muxInC_3_25_port, C(24) => muxInC_3_24_port, 
                           C(23) => muxInC_3_23_port, C(22) => muxInC_3_22_port
                           , C(21) => muxInC_3_21_port, C(20) => 
                           muxInC_3_20_port, C(19) => muxInC_3_19_port, C(18) 
                           => muxInC_3_18_port, C(17) => muxInC_3_17_port, 
                           C(16) => muxInC_3_16_port, C(15) => muxInC_3_15_port
                           , C(14) => muxInC_3_14_port, C(13) => 
                           muxInC_3_13_port, C(12) => muxInC_3_12_port, C(11) 
                           => muxInC_3_11_port, C(10) => muxInC_3_10_port, C(9)
                           => muxInC_3_9_port, C(8) => muxInC_3_8_port, C(7) =>
                           muxInC_3_7_port, C(6) => muxInC_3_6_port, C(5) => 
                           muxInC_3_5_port, C(4) => muxInC_3_4_port, C(3) => 
                           muxInC_3_3_port, C(2) => muxInC_3_2_port, C(1) => 
                           muxInC_3_1_port, C(0) => muxInC_3_0_port, D(31) => 
                           muxInD_3_31_port, D(30) => muxInD_3_30_port, D(29) 
                           => muxInD_3_29_port, D(28) => muxInD_3_28_port, 
                           D(27) => muxInD_3_27_port, D(26) => muxInD_3_26_port
                           , D(25) => muxInD_3_25_port, D(24) => 
                           muxInD_3_24_port, D(23) => muxInD_3_23_port, D(22) 
                           => muxInD_3_22_port, D(21) => muxInD_3_21_port, 
                           D(20) => muxInD_3_20_port, D(19) => muxInD_3_19_port
                           , D(18) => muxInD_3_18_port, D(17) => 
                           muxInD_3_17_port, D(16) => muxInD_3_16_port, D(15) 
                           => muxInD_3_15_port, D(14) => muxInD_3_14_port, 
                           D(13) => muxInD_3_13_port, D(12) => muxInD_3_12_port
                           , D(11) => muxInD_3_11_port, D(10) => 
                           muxInD_3_10_port, D(9) => muxInD_3_9_port, D(8) => 
                           muxInD_3_8_port, D(7) => muxInD_3_7_port, D(6) => 
                           muxInD_3_6_port, D(5) => muxInD_3_5_port, D(4) => 
                           muxInD_3_4_port, D(3) => muxInD_3_3_port, D(2) => 
                           muxInD_3_2_port, D(1) => muxInD_3_1_port, D(0) => 
                           muxInD_3_0_port, E(31) => muxInE_3_31_port, E(30) =>
                           muxInE_3_30_port, E(29) => muxInE_3_29_port, E(28) 
                           => muxInE_3_28_port, E(27) => muxInE_3_27_port, 
                           E(26) => muxInE_3_26_port, E(25) => muxInE_3_25_port
                           , E(24) => muxInE_3_24_port, E(23) => 
                           muxInE_3_23_port, E(22) => muxInE_3_22_port, E(21) 
                           => muxInE_3_21_port, E(20) => muxInE_3_20_port, 
                           E(19) => muxInE_3_19_port, E(18) => muxInE_3_18_port
                           , E(17) => muxInE_3_17_port, E(16) => 
                           muxInE_3_16_port, E(15) => muxInE_3_15_port, E(14) 
                           => muxInE_3_14_port, E(13) => muxInE_3_13_port, 
                           E(12) => muxInE_3_12_port, E(11) => muxInE_3_11_port
                           , E(10) => muxInE_3_10_port, E(9) => muxInE_3_9_port
                           , E(8) => muxInE_3_8_port, E(7) => muxInE_3_7_port, 
                           E(6) => muxInE_3_6_port, E(5) => muxInE_3_5_port, 
                           E(4) => muxInE_3_4_port, E(3) => muxInE_3_3_port, 
                           E(2) => muxInE_3_2_port, E(1) => muxInE_3_1_port, 
                           E(0) => muxInE_3_0_port, Sel(2) => B(7), Sel(1) => 
                           B(6), Sel(0) => B(5), O(31) => outmux_3_31_port, 
                           O(30) => outmux_3_30_port, O(29) => outmux_3_29_port
                           , O(28) => outmux_3_28_port, O(27) => 
                           outmux_3_27_port, O(26) => outmux_3_26_port, O(25) 
                           => outmux_3_25_port, O(24) => outmux_3_24_port, 
                           O(23) => outmux_3_23_port, O(22) => outmux_3_22_port
                           , O(21) => outmux_3_21_port, O(20) => 
                           outmux_3_20_port, O(19) => outmux_3_19_port, O(18) 
                           => outmux_3_18_port, O(17) => outmux_3_17_port, 
                           O(16) => outmux_3_16_port, O(15) => outmux_3_15_port
                           , O(14) => outmux_3_14_port, O(13) => 
                           outmux_3_13_port, O(12) => outmux_3_12_port, O(11) 
                           => outmux_3_11_port, O(10) => outmux_3_10_port, O(9)
                           => outmux_3_9_port, O(8) => outmux_3_8_port, O(7) =>
                           outmux_3_7_port, O(6) => outmux_3_6_port, O(5) => 
                           outmux_3_5_port, O(4) => outmux_3_4_port, O(3) => 
                           outmux_3_3_port, O(2) => outmux_3_2_port, O(1) => 
                           outmux_3_1_port, O(0) => outmux_3_0_port);
   MUXGEN_4 : mux_N32_4 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_4_31_port, B(30) => 
                           muxInB_4_30_port, B(29) => muxInB_4_29_port, B(28) 
                           => muxInB_4_28_port, B(27) => muxInB_4_27_port, 
                           B(26) => muxInB_4_26_port, B(25) => muxInB_4_25_port
                           , B(24) => muxInB_4_24_port, B(23) => 
                           muxInB_4_23_port, B(22) => muxInB_4_22_port, B(21) 
                           => muxInB_4_21_port, B(20) => muxInB_4_20_port, 
                           B(19) => muxInB_4_19_port, B(18) => muxInB_4_18_port
                           , B(17) => muxInB_4_17_port, B(16) => 
                           muxInB_4_16_port, B(15) => muxInB_4_15_port, B(14) 
                           => muxInB_4_14_port, B(13) => muxInB_4_13_port, 
                           B(12) => muxInB_4_12_port, B(11) => muxInB_4_11_port
                           , B(10) => muxInB_4_10_port, B(9) => muxInB_4_9_port
                           , B(8) => muxInB_4_8_port, B(7) => muxInB_4_7_port, 
                           B(6) => muxInB_4_6_port, B(5) => muxInB_4_5_port, 
                           B(4) => muxInB_4_4_port, B(3) => muxInB_4_3_port, 
                           B(2) => muxInB_4_2_port, B(1) => muxInB_4_1_port, 
                           B(0) => muxInB_4_0_port, C(31) => muxInC_4_31_port, 
                           C(30) => muxInC_4_30_port, C(29) => muxInC_4_29_port
                           , C(28) => muxInC_4_28_port, C(27) => 
                           muxInC_4_27_port, C(26) => muxInC_4_26_port, C(25) 
                           => muxInC_4_25_port, C(24) => muxInC_4_24_port, 
                           C(23) => muxInC_4_23_port, C(22) => muxInC_4_22_port
                           , C(21) => muxInC_4_21_port, C(20) => 
                           muxInC_4_20_port, C(19) => muxInC_4_19_port, C(18) 
                           => muxInC_4_18_port, C(17) => muxInC_4_17_port, 
                           C(16) => muxInC_4_16_port, C(15) => muxInC_4_15_port
                           , C(14) => muxInC_4_14_port, C(13) => 
                           muxInC_4_13_port, C(12) => muxInC_4_12_port, C(11) 
                           => muxInC_4_11_port, C(10) => muxInC_4_10_port, C(9)
                           => muxInC_4_9_port, C(8) => muxInC_4_8_port, C(7) =>
                           muxInC_4_7_port, C(6) => muxInC_4_6_port, C(5) => 
                           muxInC_4_5_port, C(4) => muxInC_4_4_port, C(3) => 
                           muxInC_4_3_port, C(2) => muxInC_4_2_port, C(1) => 
                           muxInC_4_1_port, C(0) => muxInC_4_0_port, D(31) => 
                           muxInD_4_31_port, D(30) => muxInD_4_30_port, D(29) 
                           => muxInD_4_29_port, D(28) => muxInD_4_28_port, 
                           D(27) => muxInD_4_27_port, D(26) => muxInD_4_26_port
                           , D(25) => muxInD_4_25_port, D(24) => 
                           muxInD_4_24_port, D(23) => muxInD_4_23_port, D(22) 
                           => muxInD_4_22_port, D(21) => muxInD_4_21_port, 
                           D(20) => muxInD_4_20_port, D(19) => muxInD_4_19_port
                           , D(18) => muxInD_4_18_port, D(17) => 
                           muxInD_4_17_port, D(16) => muxInD_4_16_port, D(15) 
                           => muxInD_4_15_port, D(14) => muxInD_4_14_port, 
                           D(13) => muxInD_4_13_port, D(12) => muxInD_4_12_port
                           , D(11) => muxInD_4_11_port, D(10) => 
                           muxInD_4_10_port, D(9) => muxInD_4_9_port, D(8) => 
                           muxInD_4_8_port, D(7) => muxInD_4_7_port, D(6) => 
                           muxInD_4_6_port, D(5) => muxInD_4_5_port, D(4) => 
                           muxInD_4_4_port, D(3) => muxInD_4_3_port, D(2) => 
                           muxInD_4_2_port, D(1) => muxInD_4_1_port, D(0) => 
                           muxInD_4_0_port, E(31) => muxInE_4_31_port, E(30) =>
                           muxInE_4_30_port, E(29) => muxInE_4_29_port, E(28) 
                           => muxInE_4_28_port, E(27) => muxInE_4_27_port, 
                           E(26) => muxInE_4_26_port, E(25) => muxInE_4_25_port
                           , E(24) => muxInE_4_24_port, E(23) => 
                           muxInE_4_23_port, E(22) => muxInE_4_22_port, E(21) 
                           => muxInE_4_21_port, E(20) => muxInE_4_20_port, 
                           E(19) => muxInE_4_19_port, E(18) => muxInE_4_18_port
                           , E(17) => muxInE_4_17_port, E(16) => 
                           muxInE_4_16_port, E(15) => muxInE_4_15_port, E(14) 
                           => muxInE_4_14_port, E(13) => muxInE_4_13_port, 
                           E(12) => muxInE_4_12_port, E(11) => muxInE_4_11_port
                           , E(10) => muxInE_4_10_port, E(9) => muxInE_4_9_port
                           , E(8) => muxInE_4_8_port, E(7) => muxInE_4_7_port, 
                           E(6) => muxInE_4_6_port, E(5) => muxInE_4_5_port, 
                           E(4) => muxInE_4_4_port, E(3) => muxInE_4_3_port, 
                           E(2) => muxInE_4_2_port, E(1) => muxInE_4_1_port, 
                           E(0) => muxInE_4_0_port, Sel(2) => B(9), Sel(1) => 
                           B(8), Sel(0) => B(7), O(31) => outmux_4_31_port, 
                           O(30) => outmux_4_30_port, O(29) => outmux_4_29_port
                           , O(28) => outmux_4_28_port, O(27) => 
                           outmux_4_27_port, O(26) => outmux_4_26_port, O(25) 
                           => outmux_4_25_port, O(24) => outmux_4_24_port, 
                           O(23) => outmux_4_23_port, O(22) => outmux_4_22_port
                           , O(21) => outmux_4_21_port, O(20) => 
                           outmux_4_20_port, O(19) => outmux_4_19_port, O(18) 
                           => outmux_4_18_port, O(17) => outmux_4_17_port, 
                           O(16) => outmux_4_16_port, O(15) => outmux_4_15_port
                           , O(14) => outmux_4_14_port, O(13) => 
                           outmux_4_13_port, O(12) => outmux_4_12_port, O(11) 
                           => outmux_4_11_port, O(10) => outmux_4_10_port, O(9)
                           => outmux_4_9_port, O(8) => outmux_4_8_port, O(7) =>
                           outmux_4_7_port, O(6) => outmux_4_6_port, O(5) => 
                           outmux_4_5_port, O(4) => outmux_4_4_port, O(3) => 
                           outmux_4_3_port, O(2) => outmux_4_2_port, O(1) => 
                           outmux_4_1_port, O(0) => outmux_4_0_port);
   MUXGEN_5 : mux_N32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_5_31_port, B(30) => 
                           muxInB_5_30_port, B(29) => muxInB_5_29_port, B(28) 
                           => muxInB_5_28_port, B(27) => muxInB_5_27_port, 
                           B(26) => muxInB_5_26_port, B(25) => muxInB_5_25_port
                           , B(24) => muxInB_5_24_port, B(23) => 
                           muxInB_5_23_port, B(22) => muxInB_5_22_port, B(21) 
                           => muxInB_5_21_port, B(20) => muxInB_5_20_port, 
                           B(19) => muxInB_5_19_port, B(18) => muxInB_5_18_port
                           , B(17) => muxInB_5_17_port, B(16) => 
                           muxInB_5_16_port, B(15) => muxInB_5_15_port, B(14) 
                           => muxInB_5_14_port, B(13) => muxInB_5_13_port, 
                           B(12) => muxInB_5_12_port, B(11) => muxInB_5_11_port
                           , B(10) => muxInB_5_10_port, B(9) => muxInB_5_9_port
                           , B(8) => muxInB_5_8_port, B(7) => muxInB_5_7_port, 
                           B(6) => muxInB_5_6_port, B(5) => muxInB_5_5_port, 
                           B(4) => muxInB_5_4_port, B(3) => muxInB_5_3_port, 
                           B(2) => muxInB_5_2_port, B(1) => muxInB_5_1_port, 
                           B(0) => muxInB_5_0_port, C(31) => muxInC_5_31_port, 
                           C(30) => muxInC_5_30_port, C(29) => muxInC_5_29_port
                           , C(28) => muxInC_5_28_port, C(27) => 
                           muxInC_5_27_port, C(26) => muxInC_5_26_port, C(25) 
                           => muxInC_5_25_port, C(24) => muxInC_5_24_port, 
                           C(23) => muxInC_5_23_port, C(22) => muxInC_5_22_port
                           , C(21) => muxInC_5_21_port, C(20) => 
                           muxInC_5_20_port, C(19) => muxInC_5_19_port, C(18) 
                           => muxInC_5_18_port, C(17) => muxInC_5_17_port, 
                           C(16) => muxInC_5_16_port, C(15) => muxInC_5_15_port
                           , C(14) => muxInC_5_14_port, C(13) => 
                           muxInC_5_13_port, C(12) => muxInC_5_12_port, C(11) 
                           => muxInC_5_11_port, C(10) => muxInC_5_10_port, C(9)
                           => muxInC_5_9_port, C(8) => muxInC_5_8_port, C(7) =>
                           muxInC_5_7_port, C(6) => muxInC_5_6_port, C(5) => 
                           muxInC_5_5_port, C(4) => muxInC_5_4_port, C(3) => 
                           muxInC_5_3_port, C(2) => muxInC_5_2_port, C(1) => 
                           muxInC_5_1_port, C(0) => muxInC_5_0_port, D(31) => 
                           muxInD_5_31_port, D(30) => muxInD_5_30_port, D(29) 
                           => muxInD_5_29_port, D(28) => muxInD_5_28_port, 
                           D(27) => muxInD_5_27_port, D(26) => muxInD_5_26_port
                           , D(25) => muxInD_5_25_port, D(24) => 
                           muxInD_5_24_port, D(23) => muxInD_5_23_port, D(22) 
                           => muxInD_5_22_port, D(21) => muxInD_5_21_port, 
                           D(20) => muxInD_5_20_port, D(19) => muxInD_5_19_port
                           , D(18) => muxInD_5_18_port, D(17) => 
                           muxInD_5_17_port, D(16) => muxInD_5_16_port, D(15) 
                           => muxInD_5_15_port, D(14) => muxInD_5_14_port, 
                           D(13) => muxInD_5_13_port, D(12) => muxInD_5_12_port
                           , D(11) => muxInD_5_11_port, D(10) => 
                           muxInD_5_10_port, D(9) => muxInD_5_9_port, D(8) => 
                           muxInD_5_8_port, D(7) => muxInD_5_7_port, D(6) => 
                           muxInD_5_6_port, D(5) => muxInD_5_5_port, D(4) => 
                           muxInD_5_4_port, D(3) => muxInD_5_3_port, D(2) => 
                           muxInD_5_2_port, D(1) => muxInD_5_1_port, D(0) => 
                           muxInD_5_0_port, E(31) => muxInE_5_31_port, E(30) =>
                           muxInE_5_30_port, E(29) => muxInE_5_29_port, E(28) 
                           => muxInE_5_28_port, E(27) => muxInE_5_27_port, 
                           E(26) => muxInE_5_26_port, E(25) => muxInE_5_25_port
                           , E(24) => muxInE_5_24_port, E(23) => 
                           muxInE_5_23_port, E(22) => muxInE_5_22_port, E(21) 
                           => muxInE_5_21_port, E(20) => muxInE_5_20_port, 
                           E(19) => muxInE_5_19_port, E(18) => muxInE_5_18_port
                           , E(17) => muxInE_5_17_port, E(16) => 
                           muxInE_5_16_port, E(15) => muxInE_5_15_port, E(14) 
                           => muxInE_5_14_port, E(13) => muxInE_5_13_port, 
                           E(12) => muxInE_5_12_port, E(11) => muxInE_5_11_port
                           , E(10) => muxInE_5_10_port, E(9) => muxInE_5_9_port
                           , E(8) => muxInE_5_8_port, E(7) => muxInE_5_7_port, 
                           E(6) => muxInE_5_6_port, E(5) => muxInE_5_5_port, 
                           E(4) => muxInE_5_4_port, E(3) => muxInE_5_3_port, 
                           E(2) => muxInE_5_2_port, E(1) => muxInE_5_1_port, 
                           E(0) => muxInE_5_0_port, Sel(2) => B(11), Sel(1) => 
                           B(10), Sel(0) => B(9), O(31) => outmux_5_31_port, 
                           O(30) => outmux_5_30_port, O(29) => outmux_5_29_port
                           , O(28) => outmux_5_28_port, O(27) => 
                           outmux_5_27_port, O(26) => outmux_5_26_port, O(25) 
                           => outmux_5_25_port, O(24) => outmux_5_24_port, 
                           O(23) => outmux_5_23_port, O(22) => outmux_5_22_port
                           , O(21) => outmux_5_21_port, O(20) => 
                           outmux_5_20_port, O(19) => outmux_5_19_port, O(18) 
                           => outmux_5_18_port, O(17) => outmux_5_17_port, 
                           O(16) => outmux_5_16_port, O(15) => outmux_5_15_port
                           , O(14) => outmux_5_14_port, O(13) => 
                           outmux_5_13_port, O(12) => outmux_5_12_port, O(11) 
                           => outmux_5_11_port, O(10) => outmux_5_10_port, O(9)
                           => outmux_5_9_port, O(8) => outmux_5_8_port, O(7) =>
                           outmux_5_7_port, O(6) => outmux_5_6_port, O(5) => 
                           outmux_5_5_port, O(4) => outmux_5_4_port, O(3) => 
                           outmux_5_3_port, O(2) => outmux_5_2_port, O(1) => 
                           outmux_5_1_port, O(0) => outmux_5_0_port);
   MUXGEN_6 : mux_N32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_6_31_port, B(30) => 
                           muxInB_6_30_port, B(29) => muxInB_6_29_port, B(28) 
                           => muxInB_6_28_port, B(27) => muxInB_6_27_port, 
                           B(26) => muxInB_6_26_port, B(25) => muxInB_6_25_port
                           , B(24) => muxInB_6_24_port, B(23) => 
                           muxInB_6_23_port, B(22) => muxInB_6_22_port, B(21) 
                           => muxInB_6_21_port, B(20) => muxInB_6_20_port, 
                           B(19) => muxInB_6_19_port, B(18) => muxInB_6_18_port
                           , B(17) => muxInB_6_17_port, B(16) => 
                           muxInB_6_16_port, B(15) => muxInB_6_15_port, B(14) 
                           => muxInB_6_14_port, B(13) => muxInB_6_13_port, 
                           B(12) => muxInB_6_12_port, B(11) => muxInB_6_11_port
                           , B(10) => muxInB_6_10_port, B(9) => muxInB_6_9_port
                           , B(8) => muxInB_6_8_port, B(7) => muxInB_6_7_port, 
                           B(6) => muxInB_6_6_port, B(5) => muxInB_6_5_port, 
                           B(4) => muxInB_6_4_port, B(3) => muxInB_6_3_port, 
                           B(2) => muxInB_6_2_port, B(1) => muxInB_6_1_port, 
                           B(0) => muxInB_6_0_port, C(31) => muxInC_6_31_port, 
                           C(30) => muxInC_6_30_port, C(29) => muxInC_6_29_port
                           , C(28) => muxInC_6_28_port, C(27) => 
                           muxInC_6_27_port, C(26) => muxInC_6_26_port, C(25) 
                           => muxInC_6_25_port, C(24) => muxInC_6_24_port, 
                           C(23) => muxInC_6_23_port, C(22) => muxInC_6_22_port
                           , C(21) => muxInC_6_21_port, C(20) => 
                           muxInC_6_20_port, C(19) => muxInC_6_19_port, C(18) 
                           => muxInC_6_18_port, C(17) => muxInC_6_17_port, 
                           C(16) => muxInC_6_16_port, C(15) => muxInC_6_15_port
                           , C(14) => muxInC_6_14_port, C(13) => 
                           muxInC_6_13_port, C(12) => muxInC_6_12_port, C(11) 
                           => muxInC_6_11_port, C(10) => muxInC_6_10_port, C(9)
                           => muxInC_6_9_port, C(8) => muxInC_6_8_port, C(7) =>
                           muxInC_6_7_port, C(6) => muxInC_6_6_port, C(5) => 
                           muxInC_6_5_port, C(4) => muxInC_6_4_port, C(3) => 
                           muxInC_6_3_port, C(2) => muxInC_6_2_port, C(1) => 
                           muxInC_6_1_port, C(0) => muxInC_6_0_port, D(31) => 
                           muxInD_6_31_port, D(30) => muxInD_6_30_port, D(29) 
                           => muxInD_6_29_port, D(28) => muxInD_6_28_port, 
                           D(27) => muxInD_6_27_port, D(26) => muxInD_6_26_port
                           , D(25) => muxInD_6_25_port, D(24) => 
                           muxInD_6_24_port, D(23) => muxInD_6_23_port, D(22) 
                           => muxInD_6_22_port, D(21) => muxInD_6_21_port, 
                           D(20) => muxInD_6_20_port, D(19) => muxInD_6_19_port
                           , D(18) => muxInD_6_18_port, D(17) => 
                           muxInD_6_17_port, D(16) => muxInD_6_16_port, D(15) 
                           => muxInD_6_15_port, D(14) => muxInD_6_14_port, 
                           D(13) => muxInD_6_13_port, D(12) => muxInD_6_12_port
                           , D(11) => muxInD_6_11_port, D(10) => 
                           muxInD_6_10_port, D(9) => muxInD_6_9_port, D(8) => 
                           muxInD_6_8_port, D(7) => muxInD_6_7_port, D(6) => 
                           muxInD_6_6_port, D(5) => muxInD_6_5_port, D(4) => 
                           muxInD_6_4_port, D(3) => muxInD_6_3_port, D(2) => 
                           muxInD_6_2_port, D(1) => muxInD_6_1_port, D(0) => 
                           muxInD_6_0_port, E(31) => muxInE_6_31_port, E(30) =>
                           muxInE_6_30_port, E(29) => muxInE_6_29_port, E(28) 
                           => muxInE_6_28_port, E(27) => muxInE_6_27_port, 
                           E(26) => muxInE_6_26_port, E(25) => muxInE_6_25_port
                           , E(24) => muxInE_6_24_port, E(23) => 
                           muxInE_6_23_port, E(22) => muxInE_6_22_port, E(21) 
                           => muxInE_6_21_port, E(20) => muxInE_6_20_port, 
                           E(19) => muxInE_6_19_port, E(18) => muxInE_6_18_port
                           , E(17) => muxInE_6_17_port, E(16) => 
                           muxInE_6_16_port, E(15) => muxInE_6_15_port, E(14) 
                           => muxInE_6_14_port, E(13) => muxInE_6_13_port, 
                           E(12) => muxInE_6_12_port, E(11) => muxInE_6_11_port
                           , E(10) => muxInE_6_10_port, E(9) => muxInE_6_9_port
                           , E(8) => muxInE_6_8_port, E(7) => muxInE_6_7_port, 
                           E(6) => muxInE_6_6_port, E(5) => muxInE_6_5_port, 
                           E(4) => muxInE_6_4_port, E(3) => muxInE_6_3_port, 
                           E(2) => muxInE_6_2_port, E(1) => muxInE_6_1_port, 
                           E(0) => muxInE_6_0_port, Sel(2) => B(13), Sel(1) => 
                           B(12), Sel(0) => B(11), O(31) => outmux_6_31_port, 
                           O(30) => outmux_6_30_port, O(29) => outmux_6_29_port
                           , O(28) => outmux_6_28_port, O(27) => 
                           outmux_6_27_port, O(26) => outmux_6_26_port, O(25) 
                           => outmux_6_25_port, O(24) => outmux_6_24_port, 
                           O(23) => outmux_6_23_port, O(22) => outmux_6_22_port
                           , O(21) => outmux_6_21_port, O(20) => 
                           outmux_6_20_port, O(19) => outmux_6_19_port, O(18) 
                           => outmux_6_18_port, O(17) => outmux_6_17_port, 
                           O(16) => outmux_6_16_port, O(15) => outmux_6_15_port
                           , O(14) => outmux_6_14_port, O(13) => 
                           outmux_6_13_port, O(12) => outmux_6_12_port, O(11) 
                           => outmux_6_11_port, O(10) => outmux_6_10_port, O(9)
                           => outmux_6_9_port, O(8) => outmux_6_8_port, O(7) =>
                           outmux_6_7_port, O(6) => outmux_6_6_port, O(5) => 
                           outmux_6_5_port, O(4) => outmux_6_4_port, O(3) => 
                           outmux_6_3_port, O(2) => outmux_6_2_port, O(1) => 
                           outmux_6_1_port, O(0) => outmux_6_0_port);
   MUXGEN_7 : mux_N32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => muxInB_7_31_port, B(30) => 
                           muxInB_7_30_port, B(29) => muxInB_7_29_port, B(28) 
                           => muxInB_7_28_port, B(27) => muxInB_7_27_port, 
                           B(26) => muxInB_7_26_port, B(25) => muxInB_7_25_port
                           , B(24) => muxInB_7_24_port, B(23) => 
                           muxInB_7_23_port, B(22) => muxInB_7_22_port, B(21) 
                           => muxInB_7_21_port, B(20) => muxInB_7_20_port, 
                           B(19) => muxInB_7_19_port, B(18) => muxInB_7_18_port
                           , B(17) => muxInB_7_17_port, B(16) => 
                           muxInB_7_16_port, B(15) => muxInB_7_15_port, B(14) 
                           => muxInB_7_14_port, B(13) => muxInB_7_13_port, 
                           B(12) => muxInB_7_12_port, B(11) => muxInB_7_11_port
                           , B(10) => muxInB_7_10_port, B(9) => muxInB_7_9_port
                           , B(8) => muxInB_7_8_port, B(7) => muxInB_7_7_port, 
                           B(6) => muxInB_7_6_port, B(5) => muxInB_7_5_port, 
                           B(4) => muxInB_7_4_port, B(3) => muxInB_7_3_port, 
                           B(2) => muxInB_7_2_port, B(1) => muxInB_7_1_port, 
                           B(0) => muxInB_7_0_port, C(31) => muxInC_7_31_port, 
                           C(30) => muxInC_7_30_port, C(29) => muxInC_7_29_port
                           , C(28) => muxInC_7_28_port, C(27) => 
                           muxInC_7_27_port, C(26) => muxInC_7_26_port, C(25) 
                           => muxInC_7_25_port, C(24) => muxInC_7_24_port, 
                           C(23) => muxInC_7_23_port, C(22) => muxInC_7_22_port
                           , C(21) => muxInC_7_21_port, C(20) => 
                           muxInC_7_20_port, C(19) => muxInC_7_19_port, C(18) 
                           => muxInC_7_18_port, C(17) => muxInC_7_17_port, 
                           C(16) => muxInC_7_16_port, C(15) => muxInC_7_15_port
                           , C(14) => muxInC_7_14_port, C(13) => 
                           muxInC_7_13_port, C(12) => muxInC_7_12_port, C(11) 
                           => muxInC_7_11_port, C(10) => muxInC_7_10_port, C(9)
                           => muxInC_7_9_port, C(8) => muxInC_7_8_port, C(7) =>
                           muxInC_7_7_port, C(6) => muxInC_7_6_port, C(5) => 
                           muxInC_7_5_port, C(4) => muxInC_7_4_port, C(3) => 
                           muxInC_7_3_port, C(2) => muxInC_7_2_port, C(1) => 
                           muxInC_7_1_port, C(0) => muxInC_7_0_port, D(31) => 
                           muxInD_7_31_port, D(30) => muxInD_7_30_port, D(29) 
                           => muxInD_7_29_port, D(28) => muxInD_7_28_port, 
                           D(27) => muxInD_7_27_port, D(26) => muxInD_7_26_port
                           , D(25) => muxInD_7_25_port, D(24) => 
                           muxInD_7_24_port, D(23) => muxInD_7_23_port, D(22) 
                           => muxInD_7_22_port, D(21) => muxInD_7_21_port, 
                           D(20) => muxInD_7_20_port, D(19) => muxInD_7_19_port
                           , D(18) => muxInD_7_18_port, D(17) => 
                           muxInD_7_17_port, D(16) => muxInD_7_16_port, D(15) 
                           => muxInD_7_15_port, D(14) => muxInD_7_14_port, 
                           D(13) => muxInD_7_13_port, D(12) => muxInD_7_12_port
                           , D(11) => muxInD_7_11_port, D(10) => 
                           muxInD_7_10_port, D(9) => muxInD_7_9_port, D(8) => 
                           muxInD_7_8_port, D(7) => muxInD_7_7_port, D(6) => 
                           muxInD_7_6_port, D(5) => muxInD_7_5_port, D(4) => 
                           muxInD_7_4_port, D(3) => muxInD_7_3_port, D(2) => 
                           muxInD_7_2_port, D(1) => muxInD_7_1_port, D(0) => 
                           muxInD_7_0_port, E(31) => muxInE_7_31_port, E(30) =>
                           muxInE_7_30_port, E(29) => muxInE_7_29_port, E(28) 
                           => muxInE_7_28_port, E(27) => muxInE_7_27_port, 
                           E(26) => muxInE_7_26_port, E(25) => muxInE_7_25_port
                           , E(24) => muxInE_7_24_port, E(23) => 
                           muxInE_7_23_port, E(22) => muxInE_7_22_port, E(21) 
                           => muxInE_7_21_port, E(20) => muxInE_7_20_port, 
                           E(19) => muxInE_7_19_port, E(18) => muxInE_7_18_port
                           , E(17) => muxInE_7_17_port, E(16) => 
                           muxInE_7_16_port, E(15) => muxInE_7_15_port, E(14) 
                           => muxInE_7_14_port, E(13) => muxInE_7_13_port, 
                           E(12) => muxInE_7_12_port, E(11) => muxInE_7_11_port
                           , E(10) => muxInE_7_10_port, E(9) => muxInE_7_9_port
                           , E(8) => muxInE_7_8_port, E(7) => muxInE_7_7_port, 
                           E(6) => muxInE_7_6_port, E(5) => muxInE_7_5_port, 
                           E(4) => muxInE_7_4_port, E(3) => muxInE_7_3_port, 
                           E(2) => muxInE_7_2_port, E(1) => muxInE_7_1_port, 
                           E(0) => muxInE_7_0_port, Sel(2) => B(15), Sel(1) => 
                           B(14), Sel(0) => B(13), O(31) => outmux_7_31_port, 
                           O(30) => outmux_7_30_port, O(29) => outmux_7_29_port
                           , O(28) => outmux_7_28_port, O(27) => 
                           outmux_7_27_port, O(26) => outmux_7_26_port, O(25) 
                           => outmux_7_25_port, O(24) => outmux_7_24_port, 
                           O(23) => outmux_7_23_port, O(22) => outmux_7_22_port
                           , O(21) => outmux_7_21_port, O(20) => 
                           outmux_7_20_port, O(19) => outmux_7_19_port, O(18) 
                           => outmux_7_18_port, O(17) => outmux_7_17_port, 
                           O(16) => outmux_7_16_port, O(15) => outmux_7_15_port
                           , O(14) => outmux_7_14_port, O(13) => 
                           outmux_7_13_port, O(12) => outmux_7_12_port, O(11) 
                           => outmux_7_11_port, O(10) => outmux_7_10_port, O(9)
                           => outmux_7_9_port, O(8) => outmux_7_8_port, O(7) =>
                           outmux_7_7_port, O(6) => outmux_7_6_port, O(5) => 
                           outmux_7_5_port, O(4) => outmux_7_4_port, O(3) => 
                           outmux_7_3_port, O(2) => outmux_7_2_port, O(1) => 
                           outmux_7_1_port, O(0) => outmux_7_0_port);
   Add1IL : CSA_Nbits32_0 port map( A(31) => outmux_0_31_port, A(30) => 
                           outmux_0_30_port, A(29) => outmux_0_29_port, A(28) 
                           => outmux_0_28_port, A(27) => outmux_0_27_port, 
                           A(26) => outmux_0_26_port, A(25) => outmux_0_25_port
                           , A(24) => outmux_0_24_port, A(23) => 
                           outmux_0_23_port, A(22) => outmux_0_22_port, A(21) 
                           => outmux_0_21_port, A(20) => outmux_0_20_port, 
                           A(19) => outmux_0_19_port, A(18) => outmux_0_18_port
                           , A(17) => outmux_0_17_port, A(16) => 
                           outmux_0_16_port, A(15) => outmux_0_15_port, A(14) 
                           => outmux_0_14_port, A(13) => outmux_0_13_port, 
                           A(12) => outmux_0_12_port, A(11) => outmux_0_11_port
                           , A(10) => outmux_0_10_port, A(9) => outmux_0_9_port
                           , A(8) => outmux_0_8_port, A(7) => outmux_0_7_port, 
                           A(6) => outmux_0_6_port, A(5) => outmux_0_5_port, 
                           A(4) => outmux_0_4_port, A(3) => outmux_0_3_port, 
                           A(2) => outmux_0_2_port, A(1) => outmux_0_1_port, 
                           A(0) => outmux_0_0_port, B(31) => outmux_1_31_port, 
                           B(30) => outmux_1_30_port, B(29) => outmux_1_29_port
                           , B(28) => outmux_1_28_port, B(27) => 
                           outmux_1_27_port, B(26) => outmux_1_26_port, B(25) 
                           => outmux_1_25_port, B(24) => outmux_1_24_port, 
                           B(23) => outmux_1_23_port, B(22) => outmux_1_22_port
                           , B(21) => outmux_1_21_port, B(20) => 
                           outmux_1_20_port, B(19) => outmux_1_19_port, B(18) 
                           => outmux_1_18_port, B(17) => outmux_1_17_port, 
                           B(16) => outmux_1_16_port, B(15) => outmux_1_15_port
                           , B(14) => outmux_1_14_port, B(13) => 
                           outmux_1_13_port, B(12) => outmux_1_12_port, B(11) 
                           => outmux_1_11_port, B(10) => outmux_1_10_port, B(9)
                           => outmux_1_9_port, B(8) => outmux_1_8_port, B(7) =>
                           outmux_1_7_port, B(6) => outmux_1_6_port, B(5) => 
                           outmux_1_5_port, B(4) => outmux_1_4_port, B(3) => 
                           outmux_1_3_port, B(2) => outmux_1_2_port, B(1) => 
                           outmux_1_1_port, B(0) => outmux_1_0_port, C(31) => 
                           outmux_2_31_port, C(30) => outmux_2_30_port, C(29) 
                           => outmux_2_29_port, C(28) => outmux_2_28_port, 
                           C(27) => outmux_2_27_port, C(26) => outmux_2_26_port
                           , C(25) => outmux_2_25_port, C(24) => 
                           outmux_2_24_port, C(23) => outmux_2_23_port, C(22) 
                           => outmux_2_22_port, C(21) => outmux_2_21_port, 
                           C(20) => outmux_2_20_port, C(19) => outmux_2_19_port
                           , C(18) => outmux_2_18_port, C(17) => 
                           outmux_2_17_port, C(16) => outmux_2_16_port, C(15) 
                           => outmux_2_15_port, C(14) => outmux_2_14_port, 
                           C(13) => outmux_2_13_port, C(12) => outmux_2_12_port
                           , C(11) => outmux_2_11_port, C(10) => 
                           outmux_2_10_port, C(9) => outmux_2_9_port, C(8) => 
                           outmux_2_8_port, C(7) => outmux_2_7_port, C(6) => 
                           outmux_2_6_port, C(5) => outmux_2_5_port, C(4) => 
                           outmux_2_4_port, C(3) => outmux_2_3_port, C(2) => 
                           outmux_2_2_port, C(1) => outmux_2_1_port, C(0) => 
                           outmux_2_0_port, S(31) => sum_array_0_31_port, S(30)
                           => sum_array_0_30_port, S(29) => sum_array_0_29_port
                           , S(28) => sum_array_0_28_port, S(27) => 
                           sum_array_0_27_port, S(26) => sum_array_0_26_port, 
                           S(25) => sum_array_0_25_port, S(24) => 
                           sum_array_0_24_port, S(23) => sum_array_0_23_port, 
                           S(22) => sum_array_0_22_port, S(21) => 
                           sum_array_0_21_port, S(20) => sum_array_0_20_port, 
                           S(19) => sum_array_0_19_port, S(18) => 
                           sum_array_0_18_port, S(17) => sum_array_0_17_port, 
                           S(16) => sum_array_0_16_port, S(15) => 
                           sum_array_0_15_port, S(14) => sum_array_0_14_port, 
                           S(13) => sum_array_0_13_port, S(12) => 
                           sum_array_0_12_port, S(11) => sum_array_0_11_port, 
                           S(10) => sum_array_0_10_port, S(9) => 
                           sum_array_0_9_port, S(8) => sum_array_0_8_port, S(7)
                           => sum_array_0_7_port, S(6) => sum_array_0_6_port, 
                           S(5) => sum_array_0_5_port, S(4) => 
                           sum_array_0_4_port, S(3) => sum_array_0_3_port, S(2)
                           => sum_array_0_2_port, S(1) => sum_array_0_1_port, 
                           S(0) => sum_array_0_0_port, Cout(31) => 
                           cout_array_0_31_port, Cout(30) => 
                           cout_array_0_30_port, Cout(29) => 
                           cout_array_0_29_port, Cout(28) => 
                           cout_array_0_28_port, Cout(27) => 
                           cout_array_0_27_port, Cout(26) => 
                           cout_array_0_26_port, Cout(25) => 
                           cout_array_0_25_port, Cout(24) => 
                           cout_array_0_24_port, Cout(23) => 
                           cout_array_0_23_port, Cout(22) => 
                           cout_array_0_22_port, Cout(21) => 
                           cout_array_0_21_port, Cout(20) => 
                           cout_array_0_20_port, Cout(19) => 
                           cout_array_0_19_port, Cout(18) => 
                           cout_array_0_18_port, Cout(17) => 
                           cout_array_0_17_port, Cout(16) => 
                           cout_array_0_16_port, Cout(15) => 
                           cout_array_0_15_port, Cout(14) => 
                           cout_array_0_14_port, Cout(13) => 
                           cout_array_0_13_port, Cout(12) => 
                           cout_array_0_12_port, Cout(11) => 
                           cout_array_0_11_port, Cout(10) => 
                           cout_array_0_10_port, Cout(9) => cout_array_0_9_port
                           , Cout(8) => cout_array_0_8_port, Cout(7) => 
                           cout_array_0_7_port, Cout(6) => cout_array_0_6_port,
                           Cout(5) => cout_array_0_5_port, Cout(4) => 
                           cout_array_0_4_port, Cout(3) => cout_array_0_3_port,
                           Cout(2) => cout_array_0_2_port, Cout(1) => 
                           cout_array_0_1_port, Cout(0) => net59834);
   Add2IL : CSA_Nbits32_5 port map( A(31) => outmux_3_31_port, A(30) => 
                           outmux_3_30_port, A(29) => outmux_3_29_port, A(28) 
                           => outmux_3_28_port, A(27) => outmux_3_27_port, 
                           A(26) => outmux_3_26_port, A(25) => outmux_3_25_port
                           , A(24) => outmux_3_24_port, A(23) => 
                           outmux_3_23_port, A(22) => outmux_3_22_port, A(21) 
                           => outmux_3_21_port, A(20) => outmux_3_20_port, 
                           A(19) => outmux_3_19_port, A(18) => outmux_3_18_port
                           , A(17) => outmux_3_17_port, A(16) => 
                           outmux_3_16_port, A(15) => outmux_3_15_port, A(14) 
                           => outmux_3_14_port, A(13) => outmux_3_13_port, 
                           A(12) => outmux_3_12_port, A(11) => outmux_3_11_port
                           , A(10) => outmux_3_10_port, A(9) => outmux_3_9_port
                           , A(8) => outmux_3_8_port, A(7) => outmux_3_7_port, 
                           A(6) => outmux_3_6_port, A(5) => outmux_3_5_port, 
                           A(4) => outmux_3_4_port, A(3) => outmux_3_3_port, 
                           A(2) => outmux_3_2_port, A(1) => outmux_3_1_port, 
                           A(0) => outmux_3_0_port, B(31) => outmux_4_31_port, 
                           B(30) => outmux_4_30_port, B(29) => outmux_4_29_port
                           , B(28) => outmux_4_28_port, B(27) => 
                           outmux_4_27_port, B(26) => outmux_4_26_port, B(25) 
                           => outmux_4_25_port, B(24) => outmux_4_24_port, 
                           B(23) => outmux_4_23_port, B(22) => outmux_4_22_port
                           , B(21) => outmux_4_21_port, B(20) => 
                           outmux_4_20_port, B(19) => outmux_4_19_port, B(18) 
                           => outmux_4_18_port, B(17) => outmux_4_17_port, 
                           B(16) => outmux_4_16_port, B(15) => outmux_4_15_port
                           , B(14) => outmux_4_14_port, B(13) => 
                           outmux_4_13_port, B(12) => outmux_4_12_port, B(11) 
                           => outmux_4_11_port, B(10) => outmux_4_10_port, B(9)
                           => outmux_4_9_port, B(8) => outmux_4_8_port, B(7) =>
                           outmux_4_7_port, B(6) => outmux_4_6_port, B(5) => 
                           outmux_4_5_port, B(4) => outmux_4_4_port, B(3) => 
                           outmux_4_3_port, B(2) => outmux_4_2_port, B(1) => 
                           outmux_4_1_port, B(0) => outmux_4_0_port, C(31) => 
                           outmux_5_31_port, C(30) => outmux_5_30_port, C(29) 
                           => outmux_5_29_port, C(28) => outmux_5_28_port, 
                           C(27) => outmux_5_27_port, C(26) => outmux_5_26_port
                           , C(25) => outmux_5_25_port, C(24) => 
                           outmux_5_24_port, C(23) => outmux_5_23_port, C(22) 
                           => outmux_5_22_port, C(21) => outmux_5_21_port, 
                           C(20) => outmux_5_20_port, C(19) => outmux_5_19_port
                           , C(18) => outmux_5_18_port, C(17) => 
                           outmux_5_17_port, C(16) => outmux_5_16_port, C(15) 
                           => outmux_5_15_port, C(14) => outmux_5_14_port, 
                           C(13) => outmux_5_13_port, C(12) => outmux_5_12_port
                           , C(11) => outmux_5_11_port, C(10) => 
                           outmux_5_10_port, C(9) => outmux_5_9_port, C(8) => 
                           outmux_5_8_port, C(7) => outmux_5_7_port, C(6) => 
                           outmux_5_6_port, C(5) => outmux_5_5_port, C(4) => 
                           outmux_5_4_port, C(3) => outmux_5_3_port, C(2) => 
                           outmux_5_2_port, C(1) => outmux_5_1_port, C(0) => 
                           outmux_5_0_port, S(31) => sum_array_1_31_port, S(30)
                           => sum_array_1_30_port, S(29) => sum_array_1_29_port
                           , S(28) => sum_array_1_28_port, S(27) => 
                           sum_array_1_27_port, S(26) => sum_array_1_26_port, 
                           S(25) => sum_array_1_25_port, S(24) => 
                           sum_array_1_24_port, S(23) => sum_array_1_23_port, 
                           S(22) => sum_array_1_22_port, S(21) => 
                           sum_array_1_21_port, S(20) => sum_array_1_20_port, 
                           S(19) => sum_array_1_19_port, S(18) => 
                           sum_array_1_18_port, S(17) => sum_array_1_17_port, 
                           S(16) => sum_array_1_16_port, S(15) => 
                           sum_array_1_15_port, S(14) => sum_array_1_14_port, 
                           S(13) => sum_array_1_13_port, S(12) => 
                           sum_array_1_12_port, S(11) => sum_array_1_11_port, 
                           S(10) => sum_array_1_10_port, S(9) => 
                           sum_array_1_9_port, S(8) => sum_array_1_8_port, S(7)
                           => sum_array_1_7_port, S(6) => sum_array_1_6_port, 
                           S(5) => sum_array_1_5_port, S(4) => 
                           sum_array_1_4_port, S(3) => sum_array_1_3_port, S(2)
                           => sum_array_1_2_port, S(1) => sum_array_1_1_port, 
                           S(0) => sum_array_1_0_port, Cout(31) => 
                           cout_array_1_31_port, Cout(30) => 
                           cout_array_1_30_port, Cout(29) => 
                           cout_array_1_29_port, Cout(28) => 
                           cout_array_1_28_port, Cout(27) => 
                           cout_array_1_27_port, Cout(26) => 
                           cout_array_1_26_port, Cout(25) => 
                           cout_array_1_25_port, Cout(24) => 
                           cout_array_1_24_port, Cout(23) => 
                           cout_array_1_23_port, Cout(22) => 
                           cout_array_1_22_port, Cout(21) => 
                           cout_array_1_21_port, Cout(20) => 
                           cout_array_1_20_port, Cout(19) => 
                           cout_array_1_19_port, Cout(18) => 
                           cout_array_1_18_port, Cout(17) => 
                           cout_array_1_17_port, Cout(16) => 
                           cout_array_1_16_port, Cout(15) => 
                           cout_array_1_15_port, Cout(14) => 
                           cout_array_1_14_port, Cout(13) => 
                           cout_array_1_13_port, Cout(12) => 
                           cout_array_1_12_port, Cout(11) => 
                           cout_array_1_11_port, Cout(10) => 
                           cout_array_1_10_port, Cout(9) => cout_array_1_9_port
                           , Cout(8) => cout_array_1_8_port, Cout(7) => 
                           cout_array_1_7_port, Cout(6) => cout_array_1_6_port,
                           Cout(5) => cout_array_1_5_port, Cout(4) => 
                           cout_array_1_4_port, Cout(3) => cout_array_1_3_port,
                           Cout(2) => cout_array_1_2_port, Cout(1) => 
                           cout_array_1_1_port, Cout(0) => net59833);
   Add1IIL : CSA_Nbits32_4 port map( A(31) => sum_array_0_31_port, A(30) => 
                           sum_array_0_30_port, A(29) => sum_array_0_29_port, 
                           A(28) => sum_array_0_28_port, A(27) => 
                           sum_array_0_27_port, A(26) => sum_array_0_26_port, 
                           A(25) => sum_array_0_25_port, A(24) => 
                           sum_array_0_24_port, A(23) => sum_array_0_23_port, 
                           A(22) => sum_array_0_22_port, A(21) => 
                           sum_array_0_21_port, A(20) => sum_array_0_20_port, 
                           A(19) => sum_array_0_19_port, A(18) => 
                           sum_array_0_18_port, A(17) => sum_array_0_17_port, 
                           A(16) => sum_array_0_16_port, A(15) => 
                           sum_array_0_15_port, A(14) => sum_array_0_14_port, 
                           A(13) => sum_array_0_13_port, A(12) => 
                           sum_array_0_12_port, A(11) => sum_array_0_11_port, 
                           A(10) => sum_array_0_10_port, A(9) => 
                           sum_array_0_9_port, A(8) => sum_array_0_8_port, A(7)
                           => sum_array_0_7_port, A(6) => sum_array_0_6_port, 
                           A(5) => sum_array_0_5_port, A(4) => 
                           sum_array_0_4_port, A(3) => sum_array_0_3_port, A(2)
                           => sum_array_0_2_port, A(1) => sum_array_0_1_port, 
                           A(0) => sum_array_0_0_port, B(31) => 
                           cout_array_0_31_port, B(30) => cout_array_0_30_port,
                           B(29) => cout_array_0_29_port, B(28) => 
                           cout_array_0_28_port, B(27) => cout_array_0_27_port,
                           B(26) => cout_array_0_26_port, B(25) => 
                           cout_array_0_25_port, B(24) => cout_array_0_24_port,
                           B(23) => cout_array_0_23_port, B(22) => 
                           cout_array_0_22_port, B(21) => cout_array_0_21_port,
                           B(20) => cout_array_0_20_port, B(19) => 
                           cout_array_0_19_port, B(18) => cout_array_0_18_port,
                           B(17) => cout_array_0_17_port, B(16) => 
                           cout_array_0_16_port, B(15) => cout_array_0_15_port,
                           B(14) => cout_array_0_14_port, B(13) => 
                           cout_array_0_13_port, B(12) => cout_array_0_12_port,
                           B(11) => cout_array_0_11_port, B(10) => 
                           cout_array_0_10_port, B(9) => cout_array_0_9_port, 
                           B(8) => cout_array_0_8_port, B(7) => 
                           cout_array_0_7_port, B(6) => cout_array_0_6_port, 
                           B(5) => cout_array_0_5_port, B(4) => 
                           cout_array_0_4_port, B(3) => cout_array_0_3_port, 
                           B(2) => cout_array_0_2_port, B(1) => 
                           cout_array_0_1_port, B(0) => cout_array_0_0_port, 
                           C(31) => sum_array_1_31_port, C(30) => 
                           sum_array_1_30_port, C(29) => sum_array_1_29_port, 
                           C(28) => sum_array_1_28_port, C(27) => 
                           sum_array_1_27_port, C(26) => sum_array_1_26_port, 
                           C(25) => sum_array_1_25_port, C(24) => 
                           sum_array_1_24_port, C(23) => sum_array_1_23_port, 
                           C(22) => sum_array_1_22_port, C(21) => 
                           sum_array_1_21_port, C(20) => sum_array_1_20_port, 
                           C(19) => sum_array_1_19_port, C(18) => 
                           sum_array_1_18_port, C(17) => sum_array_1_17_port, 
                           C(16) => sum_array_1_16_port, C(15) => 
                           sum_array_1_15_port, C(14) => sum_array_1_14_port, 
                           C(13) => sum_array_1_13_port, C(12) => 
                           sum_array_1_12_port, C(11) => sum_array_1_11_port, 
                           C(10) => sum_array_1_10_port, C(9) => 
                           sum_array_1_9_port, C(8) => sum_array_1_8_port, C(7)
                           => sum_array_1_7_port, C(6) => sum_array_1_6_port, 
                           C(5) => sum_array_1_5_port, C(4) => 
                           sum_array_1_4_port, C(3) => sum_array_1_3_port, C(2)
                           => sum_array_1_2_port, C(1) => sum_array_1_1_port, 
                           C(0) => sum_array_1_0_port, S(31) => 
                           sum_array_2_31_port, S(30) => sum_array_2_30_port, 
                           S(29) => sum_array_2_29_port, S(28) => 
                           sum_array_2_28_port, S(27) => sum_array_2_27_port, 
                           S(26) => sum_array_2_26_port, S(25) => 
                           sum_array_2_25_port, S(24) => sum_array_2_24_port, 
                           S(23) => sum_array_2_23_port, S(22) => 
                           sum_array_2_22_port, S(21) => sum_array_2_21_port, 
                           S(20) => sum_array_2_20_port, S(19) => 
                           sum_array_2_19_port, S(18) => sum_array_2_18_port, 
                           S(17) => sum_array_2_17_port, S(16) => 
                           sum_array_2_16_port, S(15) => sum_array_2_15_port, 
                           S(14) => sum_array_2_14_port, S(13) => 
                           sum_array_2_13_port, S(12) => sum_array_2_12_port, 
                           S(11) => sum_array_2_11_port, S(10) => 
                           sum_array_2_10_port, S(9) => sum_array_2_9_port, 
                           S(8) => sum_array_2_8_port, S(7) => 
                           sum_array_2_7_port, S(6) => sum_array_2_6_port, S(5)
                           => sum_array_2_5_port, S(4) => sum_array_2_4_port, 
                           S(3) => sum_array_2_3_port, S(2) => 
                           sum_array_2_2_port, S(1) => sum_array_2_1_port, S(0)
                           => sum_array_2_0_port, Cout(31) => 
                           cout_array_2_31_port, Cout(30) => 
                           cout_array_2_30_port, Cout(29) => 
                           cout_array_2_29_port, Cout(28) => 
                           cout_array_2_28_port, Cout(27) => 
                           cout_array_2_27_port, Cout(26) => 
                           cout_array_2_26_port, Cout(25) => 
                           cout_array_2_25_port, Cout(24) => 
                           cout_array_2_24_port, Cout(23) => 
                           cout_array_2_23_port, Cout(22) => 
                           cout_array_2_22_port, Cout(21) => 
                           cout_array_2_21_port, Cout(20) => 
                           cout_array_2_20_port, Cout(19) => 
                           cout_array_2_19_port, Cout(18) => 
                           cout_array_2_18_port, Cout(17) => 
                           cout_array_2_17_port, Cout(16) => 
                           cout_array_2_16_port, Cout(15) => 
                           cout_array_2_15_port, Cout(14) => 
                           cout_array_2_14_port, Cout(13) => 
                           cout_array_2_13_port, Cout(12) => 
                           cout_array_2_12_port, Cout(11) => 
                           cout_array_2_11_port, Cout(10) => 
                           cout_array_2_10_port, Cout(9) => cout_array_2_9_port
                           , Cout(8) => cout_array_2_8_port, Cout(7) => 
                           cout_array_2_7_port, Cout(6) => cout_array_2_6_port,
                           Cout(5) => cout_array_2_5_port, Cout(4) => 
                           cout_array_2_4_port, Cout(3) => cout_array_2_3_port,
                           Cout(2) => cout_array_2_2_port, Cout(1) => 
                           cout_array_2_1_port, Cout(0) => net59832);
   Add2IIL : CSA_Nbits32_3 port map( A(31) => cout_array_1_31_port, A(30) => 
                           cout_array_1_30_port, A(29) => cout_array_1_29_port,
                           A(28) => cout_array_1_28_port, A(27) => 
                           cout_array_1_27_port, A(26) => cout_array_1_26_port,
                           A(25) => cout_array_1_25_port, A(24) => 
                           cout_array_1_24_port, A(23) => cout_array_1_23_port,
                           A(22) => cout_array_1_22_port, A(21) => 
                           cout_array_1_21_port, A(20) => cout_array_1_20_port,
                           A(19) => cout_array_1_19_port, A(18) => 
                           cout_array_1_18_port, A(17) => cout_array_1_17_port,
                           A(16) => cout_array_1_16_port, A(15) => 
                           cout_array_1_15_port, A(14) => cout_array_1_14_port,
                           A(13) => cout_array_1_13_port, A(12) => 
                           cout_array_1_12_port, A(11) => cout_array_1_11_port,
                           A(10) => cout_array_1_10_port, A(9) => 
                           cout_array_1_9_port, A(8) => cout_array_1_8_port, 
                           A(7) => cout_array_1_7_port, A(6) => 
                           cout_array_1_6_port, A(5) => cout_array_1_5_port, 
                           A(4) => cout_array_1_4_port, A(3) => 
                           cout_array_1_3_port, A(2) => cout_array_1_2_port, 
                           A(1) => cout_array_1_1_port, A(0) => 
                           cout_array_1_0_port, B(31) => outmux_6_31_port, 
                           B(30) => outmux_6_30_port, B(29) => outmux_6_29_port
                           , B(28) => outmux_6_28_port, B(27) => 
                           outmux_6_27_port, B(26) => outmux_6_26_port, B(25) 
                           => outmux_6_25_port, B(24) => outmux_6_24_port, 
                           B(23) => outmux_6_23_port, B(22) => outmux_6_22_port
                           , B(21) => outmux_6_21_port, B(20) => 
                           outmux_6_20_port, B(19) => outmux_6_19_port, B(18) 
                           => outmux_6_18_port, B(17) => outmux_6_17_port, 
                           B(16) => outmux_6_16_port, B(15) => outmux_6_15_port
                           , B(14) => outmux_6_14_port, B(13) => 
                           outmux_6_13_port, B(12) => outmux_6_12_port, B(11) 
                           => outmux_6_11_port, B(10) => outmux_6_10_port, B(9)
                           => outmux_6_9_port, B(8) => outmux_6_8_port, B(7) =>
                           outmux_6_7_port, B(6) => outmux_6_6_port, B(5) => 
                           outmux_6_5_port, B(4) => outmux_6_4_port, B(3) => 
                           outmux_6_3_port, B(2) => outmux_6_2_port, B(1) => 
                           outmux_6_1_port, B(0) => outmux_6_0_port, C(31) => 
                           outmux_7_31_port, C(30) => outmux_7_30_port, C(29) 
                           => outmux_7_29_port, C(28) => outmux_7_28_port, 
                           C(27) => outmux_7_27_port, C(26) => outmux_7_26_port
                           , C(25) => outmux_7_25_port, C(24) => 
                           outmux_7_24_port, C(23) => outmux_7_23_port, C(22) 
                           => outmux_7_22_port, C(21) => outmux_7_21_port, 
                           C(20) => outmux_7_20_port, C(19) => outmux_7_19_port
                           , C(18) => outmux_7_18_port, C(17) => 
                           outmux_7_17_port, C(16) => outmux_7_16_port, C(15) 
                           => outmux_7_15_port, C(14) => outmux_7_14_port, 
                           C(13) => outmux_7_13_port, C(12) => outmux_7_12_port
                           , C(11) => outmux_7_11_port, C(10) => 
                           outmux_7_10_port, C(9) => outmux_7_9_port, C(8) => 
                           outmux_7_8_port, C(7) => outmux_7_7_port, C(6) => 
                           outmux_7_6_port, C(5) => outmux_7_5_port, C(4) => 
                           outmux_7_4_port, C(3) => outmux_7_3_port, C(2) => 
                           outmux_7_2_port, C(1) => outmux_7_1_port, C(0) => 
                           outmux_7_0_port, S(31) => sum_array_3_31_port, S(30)
                           => sum_array_3_30_port, S(29) => sum_array_3_29_port
                           , S(28) => sum_array_3_28_port, S(27) => 
                           sum_array_3_27_port, S(26) => sum_array_3_26_port, 
                           S(25) => sum_array_3_25_port, S(24) => 
                           sum_array_3_24_port, S(23) => sum_array_3_23_port, 
                           S(22) => sum_array_3_22_port, S(21) => 
                           sum_array_3_21_port, S(20) => sum_array_3_20_port, 
                           S(19) => sum_array_3_19_port, S(18) => 
                           sum_array_3_18_port, S(17) => sum_array_3_17_port, 
                           S(16) => sum_array_3_16_port, S(15) => 
                           sum_array_3_15_port, S(14) => sum_array_3_14_port, 
                           S(13) => sum_array_3_13_port, S(12) => 
                           sum_array_3_12_port, S(11) => sum_array_3_11_port, 
                           S(10) => sum_array_3_10_port, S(9) => 
                           sum_array_3_9_port, S(8) => sum_array_3_8_port, S(7)
                           => sum_array_3_7_port, S(6) => sum_array_3_6_port, 
                           S(5) => sum_array_3_5_port, S(4) => 
                           sum_array_3_4_port, S(3) => sum_array_3_3_port, S(2)
                           => sum_array_3_2_port, S(1) => sum_array_3_1_port, 
                           S(0) => sum_array_3_0_port, Cout(31) => 
                           cout_array_3_31_port, Cout(30) => 
                           cout_array_3_30_port, Cout(29) => 
                           cout_array_3_29_port, Cout(28) => 
                           cout_array_3_28_port, Cout(27) => 
                           cout_array_3_27_port, Cout(26) => 
                           cout_array_3_26_port, Cout(25) => 
                           cout_array_3_25_port, Cout(24) => 
                           cout_array_3_24_port, Cout(23) => 
                           cout_array_3_23_port, Cout(22) => 
                           cout_array_3_22_port, Cout(21) => 
                           cout_array_3_21_port, Cout(20) => 
                           cout_array_3_20_port, Cout(19) => 
                           cout_array_3_19_port, Cout(18) => 
                           cout_array_3_18_port, Cout(17) => 
                           cout_array_3_17_port, Cout(16) => 
                           cout_array_3_16_port, Cout(15) => 
                           cout_array_3_15_port, Cout(14) => 
                           cout_array_3_14_port, Cout(13) => 
                           cout_array_3_13_port, Cout(12) => 
                           cout_array_3_12_port, Cout(11) => 
                           cout_array_3_11_port, Cout(10) => 
                           cout_array_3_10_port, Cout(9) => cout_array_3_9_port
                           , Cout(8) => cout_array_3_8_port, Cout(7) => 
                           cout_array_3_7_port, Cout(6) => cout_array_3_6_port,
                           Cout(5) => cout_array_3_5_port, Cout(4) => 
                           cout_array_3_4_port, Cout(3) => cout_array_3_3_port,
                           Cout(2) => cout_array_3_2_port, Cout(1) => 
                           cout_array_3_1_port, Cout(0) => net59831);
   Add1IIIL : CSA_Nbits32_2 port map( A(31) => sum_array_2_31_port, A(30) => 
                           sum_array_2_30_port, A(29) => sum_array_2_29_port, 
                           A(28) => sum_array_2_28_port, A(27) => 
                           sum_array_2_27_port, A(26) => sum_array_2_26_port, 
                           A(25) => sum_array_2_25_port, A(24) => 
                           sum_array_2_24_port, A(23) => sum_array_2_23_port, 
                           A(22) => sum_array_2_22_port, A(21) => 
                           sum_array_2_21_port, A(20) => sum_array_2_20_port, 
                           A(19) => sum_array_2_19_port, A(18) => 
                           sum_array_2_18_port, A(17) => sum_array_2_17_port, 
                           A(16) => sum_array_2_16_port, A(15) => 
                           sum_array_2_15_port, A(14) => sum_array_2_14_port, 
                           A(13) => sum_array_2_13_port, A(12) => 
                           sum_array_2_12_port, A(11) => sum_array_2_11_port, 
                           A(10) => sum_array_2_10_port, A(9) => 
                           sum_array_2_9_port, A(8) => sum_array_2_8_port, A(7)
                           => sum_array_2_7_port, A(6) => sum_array_2_6_port, 
                           A(5) => sum_array_2_5_port, A(4) => 
                           sum_array_2_4_port, A(3) => sum_array_2_3_port, A(2)
                           => sum_array_2_2_port, A(1) => sum_array_2_1_port, 
                           A(0) => sum_array_2_0_port, B(31) => 
                           cout_array_2_31_port, B(30) => cout_array_2_30_port,
                           B(29) => cout_array_2_29_port, B(28) => 
                           cout_array_2_28_port, B(27) => cout_array_2_27_port,
                           B(26) => cout_array_2_26_port, B(25) => 
                           cout_array_2_25_port, B(24) => cout_array_2_24_port,
                           B(23) => cout_array_2_23_port, B(22) => 
                           cout_array_2_22_port, B(21) => cout_array_2_21_port,
                           B(20) => cout_array_2_20_port, B(19) => 
                           cout_array_2_19_port, B(18) => cout_array_2_18_port,
                           B(17) => cout_array_2_17_port, B(16) => 
                           cout_array_2_16_port, B(15) => cout_array_2_15_port,
                           B(14) => cout_array_2_14_port, B(13) => 
                           cout_array_2_13_port, B(12) => cout_array_2_12_port,
                           B(11) => cout_array_2_11_port, B(10) => 
                           cout_array_2_10_port, B(9) => cout_array_2_9_port, 
                           B(8) => cout_array_2_8_port, B(7) => 
                           cout_array_2_7_port, B(6) => cout_array_2_6_port, 
                           B(5) => cout_array_2_5_port, B(4) => 
                           cout_array_2_4_port, B(3) => cout_array_2_3_port, 
                           B(2) => cout_array_2_2_port, B(1) => 
                           cout_array_2_1_port, B(0) => cout_array_2_0_port, 
                           C(31) => sum_array_3_31_port, C(30) => 
                           sum_array_3_30_port, C(29) => sum_array_3_29_port, 
                           C(28) => sum_array_3_28_port, C(27) => 
                           sum_array_3_27_port, C(26) => sum_array_3_26_port, 
                           C(25) => sum_array_3_25_port, C(24) => 
                           sum_array_3_24_port, C(23) => sum_array_3_23_port, 
                           C(22) => sum_array_3_22_port, C(21) => 
                           sum_array_3_21_port, C(20) => sum_array_3_20_port, 
                           C(19) => sum_array_3_19_port, C(18) => 
                           sum_array_3_18_port, C(17) => sum_array_3_17_port, 
                           C(16) => sum_array_3_16_port, C(15) => 
                           sum_array_3_15_port, C(14) => sum_array_3_14_port, 
                           C(13) => sum_array_3_13_port, C(12) => 
                           sum_array_3_12_port, C(11) => sum_array_3_11_port, 
                           C(10) => sum_array_3_10_port, C(9) => 
                           sum_array_3_9_port, C(8) => sum_array_3_8_port, C(7)
                           => sum_array_3_7_port, C(6) => sum_array_3_6_port, 
                           C(5) => sum_array_3_5_port, C(4) => 
                           sum_array_3_4_port, C(3) => sum_array_3_3_port, C(2)
                           => sum_array_3_2_port, C(1) => sum_array_3_1_port, 
                           C(0) => sum_array_3_0_port, S(31) => 
                           sum_array_4_31_port, S(30) => sum_array_4_30_port, 
                           S(29) => sum_array_4_29_port, S(28) => 
                           sum_array_4_28_port, S(27) => sum_array_4_27_port, 
                           S(26) => sum_array_4_26_port, S(25) => 
                           sum_array_4_25_port, S(24) => sum_array_4_24_port, 
                           S(23) => sum_array_4_23_port, S(22) => 
                           sum_array_4_22_port, S(21) => sum_array_4_21_port, 
                           S(20) => sum_array_4_20_port, S(19) => 
                           sum_array_4_19_port, S(18) => sum_array_4_18_port, 
                           S(17) => sum_array_4_17_port, S(16) => 
                           sum_array_4_16_port, S(15) => sum_array_4_15_port, 
                           S(14) => sum_array_4_14_port, S(13) => 
                           sum_array_4_13_port, S(12) => sum_array_4_12_port, 
                           S(11) => sum_array_4_11_port, S(10) => 
                           sum_array_4_10_port, S(9) => sum_array_4_9_port, 
                           S(8) => sum_array_4_8_port, S(7) => 
                           sum_array_4_7_port, S(6) => sum_array_4_6_port, S(5)
                           => sum_array_4_5_port, S(4) => sum_array_4_4_port, 
                           S(3) => sum_array_4_3_port, S(2) => 
                           sum_array_4_2_port, S(1) => sum_array_4_1_port, S(0)
                           => sum_array_4_0_port, Cout(31) => 
                           cout_array_4_31_port, Cout(30) => 
                           cout_array_4_30_port, Cout(29) => 
                           cout_array_4_29_port, Cout(28) => 
                           cout_array_4_28_port, Cout(27) => 
                           cout_array_4_27_port, Cout(26) => 
                           cout_array_4_26_port, Cout(25) => 
                           cout_array_4_25_port, Cout(24) => 
                           cout_array_4_24_port, Cout(23) => 
                           cout_array_4_23_port, Cout(22) => 
                           cout_array_4_22_port, Cout(21) => 
                           cout_array_4_21_port, Cout(20) => 
                           cout_array_4_20_port, Cout(19) => 
                           cout_array_4_19_port, Cout(18) => 
                           cout_array_4_18_port, Cout(17) => 
                           cout_array_4_17_port, Cout(16) => 
                           cout_array_4_16_port, Cout(15) => 
                           cout_array_4_15_port, Cout(14) => 
                           cout_array_4_14_port, Cout(13) => 
                           cout_array_4_13_port, Cout(12) => 
                           cout_array_4_12_port, Cout(11) => 
                           cout_array_4_11_port, Cout(10) => 
                           cout_array_4_10_port, Cout(9) => cout_array_4_9_port
                           , Cout(8) => cout_array_4_8_port, Cout(7) => 
                           cout_array_4_7_port, Cout(6) => cout_array_4_6_port,
                           Cout(5) => cout_array_4_5_port, Cout(4) => 
                           cout_array_4_4_port, Cout(3) => cout_array_4_3_port,
                           Cout(2) => cout_array_4_2_port, Cout(1) => 
                           cout_array_4_1_port, Cout(0) => net59830);
   AddRCA : CSA_Nbits32_1 port map( A(31) => sum_array_4_31_port, A(30) => 
                           sum_array_4_30_port, A(29) => sum_array_4_29_port, 
                           A(28) => sum_array_4_28_port, A(27) => 
                           sum_array_4_27_port, A(26) => sum_array_4_26_port, 
                           A(25) => sum_array_4_25_port, A(24) => 
                           sum_array_4_24_port, A(23) => sum_array_4_23_port, 
                           A(22) => sum_array_4_22_port, A(21) => 
                           sum_array_4_21_port, A(20) => sum_array_4_20_port, 
                           A(19) => sum_array_4_19_port, A(18) => 
                           sum_array_4_18_port, A(17) => sum_array_4_17_port, 
                           A(16) => sum_array_4_16_port, A(15) => 
                           sum_array_4_15_port, A(14) => sum_array_4_14_port, 
                           A(13) => sum_array_4_13_port, A(12) => 
                           sum_array_4_12_port, A(11) => sum_array_4_11_port, 
                           A(10) => sum_array_4_10_port, A(9) => 
                           sum_array_4_9_port, A(8) => sum_array_4_8_port, A(7)
                           => sum_array_4_7_port, A(6) => sum_array_4_6_port, 
                           A(5) => sum_array_4_5_port, A(4) => 
                           sum_array_4_4_port, A(3) => sum_array_4_3_port, A(2)
                           => sum_array_4_2_port, A(1) => sum_array_4_1_port, 
                           A(0) => sum_array_4_0_port, B(31) => 
                           cout_array_4_31_port, B(30) => cout_array_4_30_port,
                           B(29) => cout_array_4_29_port, B(28) => 
                           cout_array_4_28_port, B(27) => cout_array_4_27_port,
                           B(26) => cout_array_4_26_port, B(25) => 
                           cout_array_4_25_port, B(24) => cout_array_4_24_port,
                           B(23) => cout_array_4_23_port, B(22) => 
                           cout_array_4_22_port, B(21) => cout_array_4_21_port,
                           B(20) => cout_array_4_20_port, B(19) => 
                           cout_array_4_19_port, B(18) => cout_array_4_18_port,
                           B(17) => cout_array_4_17_port, B(16) => 
                           cout_array_4_16_port, B(15) => cout_array_4_15_port,
                           B(14) => cout_array_4_14_port, B(13) => 
                           cout_array_4_13_port, B(12) => cout_array_4_12_port,
                           B(11) => cout_array_4_11_port, B(10) => 
                           cout_array_4_10_port, B(9) => cout_array_4_9_port, 
                           B(8) => cout_array_4_8_port, B(7) => 
                           cout_array_4_7_port, B(6) => cout_array_4_6_port, 
                           B(5) => cout_array_4_5_port, B(4) => 
                           cout_array_4_4_port, B(3) => cout_array_4_3_port, 
                           B(2) => cout_array_4_2_port, B(1) => 
                           cout_array_4_1_port, B(0) => cout_array_4_0_port, 
                           C(31) => cout_array_3_31_port, C(30) => 
                           cout_array_3_30_port, C(29) => cout_array_3_29_port,
                           C(28) => cout_array_3_28_port, C(27) => 
                           cout_array_3_27_port, C(26) => cout_array_3_26_port,
                           C(25) => cout_array_3_25_port, C(24) => 
                           cout_array_3_24_port, C(23) => cout_array_3_23_port,
                           C(22) => cout_array_3_22_port, C(21) => 
                           cout_array_3_21_port, C(20) => cout_array_3_20_port,
                           C(19) => cout_array_3_19_port, C(18) => 
                           cout_array_3_18_port, C(17) => cout_array_3_17_port,
                           C(16) => cout_array_3_16_port, C(15) => 
                           cout_array_3_15_port, C(14) => cout_array_3_14_port,
                           C(13) => cout_array_3_13_port, C(12) => 
                           cout_array_3_12_port, C(11) => cout_array_3_11_port,
                           C(10) => cout_array_3_10_port, C(9) => 
                           cout_array_3_9_port, C(8) => cout_array_3_8_port, 
                           C(7) => cout_array_3_7_port, C(6) => 
                           cout_array_3_6_port, C(5) => cout_array_3_5_port, 
                           C(4) => cout_array_3_4_port, C(3) => 
                           cout_array_3_3_port, C(2) => cout_array_3_2_port, 
                           C(1) => cout_array_3_1_port, C(0) => 
                           cout_array_3_0_port, S(31) => sum_array_5_31_port, 
                           S(30) => sum_array_5_30_port, S(29) => 
                           sum_array_5_29_port, S(28) => sum_array_5_28_port, 
                           S(27) => sum_array_5_27_port, S(26) => 
                           sum_array_5_26_port, S(25) => sum_array_5_25_port, 
                           S(24) => sum_array_5_24_port, S(23) => 
                           sum_array_5_23_port, S(22) => sum_array_5_22_port, 
                           S(21) => sum_array_5_21_port, S(20) => 
                           sum_array_5_20_port, S(19) => sum_array_5_19_port, 
                           S(18) => sum_array_5_18_port, S(17) => 
                           sum_array_5_17_port, S(16) => sum_array_5_16_port, 
                           S(15) => sum_array_5_15_port, S(14) => 
                           sum_array_5_14_port, S(13) => sum_array_5_13_port, 
                           S(12) => sum_array_5_12_port, S(11) => 
                           sum_array_5_11_port, S(10) => sum_array_5_10_port, 
                           S(9) => sum_array_5_9_port, S(8) => 
                           sum_array_5_8_port, S(7) => sum_array_5_7_port, S(6)
                           => sum_array_5_6_port, S(5) => sum_array_5_5_port, 
                           S(4) => sum_array_5_4_port, S(3) => 
                           sum_array_5_3_port, S(2) => sum_array_5_2_port, S(1)
                           => sum_array_5_1_port, S(0) => sum_array_5_0_port, 
                           Cout(31) => cout_array_5_31_port, Cout(30) => 
                           cout_array_5_30_port, Cout(29) => 
                           cout_array_5_29_port, Cout(28) => 
                           cout_array_5_28_port, Cout(27) => 
                           cout_array_5_27_port, Cout(26) => 
                           cout_array_5_26_port, Cout(25) => 
                           cout_array_5_25_port, Cout(24) => 
                           cout_array_5_24_port, Cout(23) => 
                           cout_array_5_23_port, Cout(22) => 
                           cout_array_5_22_port, Cout(21) => 
                           cout_array_5_21_port, Cout(20) => 
                           cout_array_5_20_port, Cout(19) => 
                           cout_array_5_19_port, Cout(18) => 
                           cout_array_5_18_port, Cout(17) => 
                           cout_array_5_17_port, Cout(16) => 
                           cout_array_5_16_port, Cout(15) => 
                           cout_array_5_15_port, Cout(14) => 
                           cout_array_5_14_port, Cout(13) => 
                           cout_array_5_13_port, Cout(12) => 
                           cout_array_5_12_port, Cout(11) => 
                           cout_array_5_11_port, Cout(10) => 
                           cout_array_5_10_port, Cout(9) => cout_array_5_9_port
                           , Cout(8) => cout_array_5_8_port, Cout(7) => 
                           cout_array_5_7_port, Cout(6) => cout_array_5_6_port,
                           Cout(5) => cout_array_5_5_port, Cout(4) => 
                           cout_array_5_4_port, Cout(3) => cout_array_5_3_port,
                           Cout(2) => cout_array_5_2_port, Cout(1) => 
                           cout_array_5_1_port, Cout(0) => net59829);
   P4adder : cla_adder_N32_1 port map( A(31) => sum_array_5_31_port, A(30) => 
                           sum_array_5_30_port, A(29) => sum_array_5_29_port, 
                           A(28) => sum_array_5_28_port, A(27) => 
                           sum_array_5_27_port, A(26) => sum_array_5_26_port, 
                           A(25) => sum_array_5_25_port, A(24) => 
                           sum_array_5_24_port, A(23) => sum_array_5_23_port, 
                           A(22) => sum_array_5_22_port, A(21) => 
                           sum_array_5_21_port, A(20) => sum_array_5_20_port, 
                           A(19) => sum_array_5_19_port, A(18) => 
                           sum_array_5_18_port, A(17) => sum_array_5_17_port, 
                           A(16) => sum_array_5_16_port, A(15) => 
                           sum_array_5_15_port, A(14) => sum_array_5_14_port, 
                           A(13) => sum_array_5_13_port, A(12) => 
                           sum_array_5_12_port, A(11) => sum_array_5_11_port, 
                           A(10) => sum_array_5_10_port, A(9) => 
                           sum_array_5_9_port, A(8) => sum_array_5_8_port, A(7)
                           => sum_array_5_7_port, A(6) => sum_array_5_6_port, 
                           A(5) => sum_array_5_5_port, A(4) => 
                           sum_array_5_4_port, A(3) => sum_array_5_3_port, A(2)
                           => sum_array_5_2_port, A(1) => sum_array_5_1_port, 
                           A(0) => sum_array_5_0_port, B(31) => 
                           cout_array_5_31_port, B(30) => cout_array_5_30_port,
                           B(29) => cout_array_5_29_port, B(28) => 
                           cout_array_5_28_port, B(27) => cout_array_5_27_port,
                           B(26) => cout_array_5_26_port, B(25) => 
                           cout_array_5_25_port, B(24) => cout_array_5_24_port,
                           B(23) => cout_array_5_23_port, B(22) => 
                           cout_array_5_22_port, B(21) => cout_array_5_21_port,
                           B(20) => cout_array_5_20_port, B(19) => 
                           cout_array_5_19_port, B(18) => cout_array_5_18_port,
                           B(17) => cout_array_5_17_port, B(16) => 
                           cout_array_5_16_port, B(15) => cout_array_5_15_port,
                           B(14) => cout_array_5_14_port, B(13) => 
                           cout_array_5_13_port, B(12) => cout_array_5_12_port,
                           B(11) => cout_array_5_11_port, B(10) => 
                           cout_array_5_10_port, B(9) => cout_array_5_9_port, 
                           B(8) => cout_array_5_8_port, B(7) => 
                           cout_array_5_7_port, B(6) => cout_array_5_6_port, 
                           B(5) => cout_array_5_5_port, B(4) => 
                           cout_array_5_4_port, B(3) => cout_array_5_3_port, 
                           B(2) => cout_array_5_2_port, B(1) => 
                           cout_array_5_1_port, B(0) => cout_array_5_0_port, Ci
                           => X_Logic0_port, Cout => net6197, Sum(31) => Y(31),
                           Sum(30) => Y(30), Sum(29) => Y(29), Sum(28) => Y(28)
                           , Sum(27) => Y(27), Sum(26) => Y(26), Sum(25) => 
                           Y(25), Sum(24) => Y(24), Sum(23) => Y(23), Sum(22) 
                           => Y(22), Sum(21) => Y(21), Sum(20) => Y(20), 
                           Sum(19) => Y(19), Sum(18) => Y(18), Sum(17) => Y(17)
                           , Sum(16) => Y(16), Sum(15) => Y(15), Sum(14) => 
                           Y(14), Sum(13) => Y(13), Sum(12) => Y(12), Sum(11) 
                           => Y(11), Sum(10) => Y(10), Sum(9) => Y(9), Sum(8) 
                           => Y(8), Sum(7) => Y(7), Sum(6) => Y(6), Sum(5) => 
                           Y(5), Sum(4) => Y(4), Sum(3) => Y(3), Sum(2) => Y(2)
                           , Sum(1) => Y(1), Sum(0) => Y(0));
   cout_array_1_0_port <= '0';
   cout_array_2_0_port <= '0';
   cout_array_3_0_port <= '0';
   cout_array_4_0_port <= '0';
   cout_array_5_0_port <= '0';
   cout_array_0_0_port <= '0';
   muxInE_7_0_port <= '0';
   muxInE_7_1_port <= '0';
   muxInE_7_2_port <= '0';
   muxInE_7_3_port <= '0';
   muxInE_7_4_port <= '0';
   muxInE_7_5_port <= '0';
   muxInE_7_6_port <= '0';
   muxInE_7_7_port <= '0';
   muxInE_7_8_port <= '0';
   muxInE_7_9_port <= '0';
   muxInE_7_10_port <= '0';
   muxInE_7_11_port <= '0';
   muxInE_7_12_port <= '0';
   muxInE_7_13_port <= '0';
   muxInE_7_14_port <= '0';
   muxInD_7_0_port <= '0';
   muxInD_7_1_port <= '0';
   muxInD_7_2_port <= '0';
   muxInD_7_3_port <= '0';
   muxInD_7_4_port <= '0';
   muxInD_7_5_port <= '0';
   muxInD_7_6_port <= '0';
   muxInD_7_7_port <= '0';
   muxInD_7_8_port <= '0';
   muxInD_7_9_port <= '0';
   muxInD_7_10_port <= '0';
   muxInD_7_11_port <= '0';
   muxInD_7_12_port <= '0';
   muxInD_7_13_port <= '0';
   muxInD_7_14_port <= '0';
   muxInC_7_0_port <= '0';
   muxInC_7_1_port <= '0';
   muxInC_7_2_port <= '0';
   muxInC_7_3_port <= '0';
   muxInC_7_4_port <= '0';
   muxInC_7_5_port <= '0';
   muxInC_7_6_port <= '0';
   muxInC_7_7_port <= '0';
   muxInC_7_8_port <= '0';
   muxInC_7_9_port <= '0';
   muxInC_7_10_port <= '0';
   muxInC_7_11_port <= '0';
   muxInC_7_12_port <= '0';
   muxInC_7_13_port <= '0';
   muxInB_7_0_port <= '0';
   muxInB_7_1_port <= '0';
   muxInB_7_2_port <= '0';
   muxInB_7_3_port <= '0';
   muxInB_7_4_port <= '0';
   muxInB_7_5_port <= '0';
   muxInB_7_6_port <= '0';
   muxInB_7_7_port <= '0';
   muxInB_7_8_port <= '0';
   muxInB_7_9_port <= '0';
   muxInB_7_10_port <= '0';
   muxInB_7_11_port <= '0';
   muxInB_7_12_port <= '0';
   muxInB_7_13_port <= '0';
   muxInE_6_0_port <= '0';
   muxInE_6_1_port <= '0';
   muxInE_6_2_port <= '0';
   muxInE_6_3_port <= '0';
   muxInE_6_4_port <= '0';
   muxInE_6_5_port <= '0';
   muxInE_6_6_port <= '0';
   muxInE_6_7_port <= '0';
   muxInE_6_8_port <= '0';
   muxInE_6_9_port <= '0';
   muxInE_6_10_port <= '0';
   muxInE_6_11_port <= '0';
   muxInE_6_12_port <= '0';
   muxInD_6_0_port <= '0';
   muxInD_6_1_port <= '0';
   muxInD_6_2_port <= '0';
   muxInD_6_3_port <= '0';
   muxInD_6_4_port <= '0';
   muxInD_6_5_port <= '0';
   muxInD_6_6_port <= '0';
   muxInD_6_7_port <= '0';
   muxInD_6_8_port <= '0';
   muxInD_6_9_port <= '0';
   muxInD_6_10_port <= '0';
   muxInD_6_11_port <= '0';
   muxInD_6_12_port <= '0';
   muxInC_6_0_port <= '0';
   muxInC_6_1_port <= '0';
   muxInC_6_2_port <= '0';
   muxInC_6_3_port <= '0';
   muxInC_6_4_port <= '0';
   muxInC_6_5_port <= '0';
   muxInC_6_6_port <= '0';
   muxInC_6_7_port <= '0';
   muxInC_6_8_port <= '0';
   muxInC_6_9_port <= '0';
   muxInC_6_10_port <= '0';
   muxInC_6_11_port <= '0';
   muxInB_6_0_port <= '0';
   muxInB_6_1_port <= '0';
   muxInB_6_2_port <= '0';
   muxInB_6_3_port <= '0';
   muxInB_6_4_port <= '0';
   muxInB_6_5_port <= '0';
   muxInB_6_6_port <= '0';
   muxInB_6_7_port <= '0';
   muxInB_6_8_port <= '0';
   muxInB_6_9_port <= '0';
   muxInB_6_10_port <= '0';
   muxInB_6_11_port <= '0';
   muxInE_5_0_port <= '0';
   muxInE_5_1_port <= '0';
   muxInE_5_2_port <= '0';
   muxInE_5_3_port <= '0';
   muxInE_5_4_port <= '0';
   muxInE_5_5_port <= '0';
   muxInE_5_6_port <= '0';
   muxInE_5_7_port <= '0';
   muxInE_5_8_port <= '0';
   muxInE_5_9_port <= '0';
   muxInE_5_10_port <= '0';
   muxInD_5_0_port <= '0';
   muxInD_5_1_port <= '0';
   muxInD_5_2_port <= '0';
   muxInD_5_3_port <= '0';
   muxInD_5_4_port <= '0';
   muxInD_5_5_port <= '0';
   muxInD_5_6_port <= '0';
   muxInD_5_7_port <= '0';
   muxInD_5_8_port <= '0';
   muxInD_5_9_port <= '0';
   muxInD_5_10_port <= '0';
   muxInC_5_0_port <= '0';
   muxInC_5_1_port <= '0';
   muxInC_5_2_port <= '0';
   muxInC_5_3_port <= '0';
   muxInC_5_4_port <= '0';
   muxInC_5_5_port <= '0';
   muxInC_5_6_port <= '0';
   muxInC_5_7_port <= '0';
   muxInC_5_8_port <= '0';
   muxInC_5_9_port <= '0';
   muxInB_5_0_port <= '0';
   muxInB_5_1_port <= '0';
   muxInB_5_2_port <= '0';
   muxInB_5_3_port <= '0';
   muxInB_5_4_port <= '0';
   muxInB_5_5_port <= '0';
   muxInB_5_6_port <= '0';
   muxInB_5_7_port <= '0';
   muxInB_5_8_port <= '0';
   muxInB_5_9_port <= '0';
   muxInE_4_0_port <= '0';
   muxInE_4_1_port <= '0';
   muxInE_4_2_port <= '0';
   muxInE_4_3_port <= '0';
   muxInE_4_4_port <= '0';
   muxInE_4_5_port <= '0';
   muxInE_4_6_port <= '0';
   muxInE_4_7_port <= '0';
   muxInE_4_8_port <= '0';
   muxInD_4_0_port <= '0';
   muxInD_4_1_port <= '0';
   muxInD_4_2_port <= '0';
   muxInD_4_3_port <= '0';
   muxInD_4_4_port <= '0';
   muxInD_4_5_port <= '0';
   muxInD_4_6_port <= '0';
   muxInD_4_7_port <= '0';
   muxInD_4_8_port <= '0';
   muxInC_4_0_port <= '0';
   muxInC_4_1_port <= '0';
   muxInC_4_2_port <= '0';
   muxInC_4_3_port <= '0';
   muxInC_4_4_port <= '0';
   muxInC_4_5_port <= '0';
   muxInC_4_6_port <= '0';
   muxInC_4_7_port <= '0';
   muxInB_4_0_port <= '0';
   muxInB_4_1_port <= '0';
   muxInB_4_2_port <= '0';
   muxInB_4_3_port <= '0';
   muxInB_4_4_port <= '0';
   muxInB_4_5_port <= '0';
   muxInB_4_6_port <= '0';
   muxInB_4_7_port <= '0';
   muxInE_3_0_port <= '0';
   muxInE_3_1_port <= '0';
   muxInE_3_2_port <= '0';
   muxInE_3_3_port <= '0';
   muxInE_3_4_port <= '0';
   muxInE_3_5_port <= '0';
   muxInE_3_6_port <= '0';
   muxInD_3_0_port <= '0';
   muxInD_3_1_port <= '0';
   muxInD_3_2_port <= '0';
   muxInD_3_3_port <= '0';
   muxInD_3_4_port <= '0';
   muxInD_3_5_port <= '0';
   muxInD_3_6_port <= '0';
   muxInC_3_0_port <= '0';
   muxInC_3_1_port <= '0';
   muxInC_3_2_port <= '0';
   muxInC_3_3_port <= '0';
   muxInC_3_4_port <= '0';
   muxInC_3_5_port <= '0';
   muxInB_3_0_port <= '0';
   muxInB_3_1_port <= '0';
   muxInB_3_2_port <= '0';
   muxInB_3_3_port <= '0';
   muxInB_3_4_port <= '0';
   muxInB_3_5_port <= '0';
   muxInE_2_0_port <= '0';
   muxInE_2_1_port <= '0';
   muxInE_2_2_port <= '0';
   muxInE_2_3_port <= '0';
   muxInE_2_4_port <= '0';
   muxInD_2_0_port <= '0';
   muxInD_2_1_port <= '0';
   muxInD_2_2_port <= '0';
   muxInD_2_3_port <= '0';
   muxInD_2_4_port <= '0';
   muxInC_2_0_port <= '0';
   muxInC_2_1_port <= '0';
   muxInC_2_2_port <= '0';
   muxInC_2_3_port <= '0';
   muxInB_2_0_port <= '0';
   muxInB_2_1_port <= '0';
   muxInB_2_2_port <= '0';
   muxInB_2_3_port <= '0';
   muxInE_1_0_port <= '0';
   muxInE_1_1_port <= '0';
   muxInE_1_2_port <= '0';
   muxInD_1_0_port <= '0';
   muxInD_1_1_port <= '0';
   muxInD_1_2_port <= '0';
   muxInC_1_0_port <= '0';
   muxInC_1_1_port <= '0';
   muxInB_1_0_port <= '0';
   muxInB_1_1_port <= '0';
   muxInE_0_0_port <= '0';
   muxInD_0_0_port <= '0';
   U248 : BUF_X1 port map( A => A(12), Z => n25);
   U249 : BUF_X1 port map( A => A(8), Z => n18);
   U250 : BUF_X1 port map( A => A(11), Z => n22);
   U251 : BUF_X1 port map( A => A(14), Z => n27);
   U252 : BUF_X1 port map( A => A(10), Z => n21);
   U253 : BUF_X2 port map( A => A(13), Z => n26);
   U254 : BUF_X2 port map( A => A(9), Z => n19);
   U255 : BUF_X2 port map( A => A(3), Z => n11);
   U256 : BUF_X2 port map( A => A(7), Z => n17);
   U257 : BUF_X2 port map( A => A(1), Z => n10);
   U258 : BUF_X2 port map( A => A(0), Z => n2);
   U259 : BUF_X2 port map( A => A(5), Z => n14);
   U260 : BUF_X1 port map( A => A(6), Z => n15);
   U261 : BUF_X1 port map( A => A(0), Z => n3);
   U262 : BUF_X1 port map( A => A(4), Z => n13);
   U263 : BUF_X1 port map( A => A(15), Z => n28);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity adder_sub_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout : 
         out std_logic;  Sum : out std_logic_vector (31 downto 0));

end adder_sub_N32;

architecture SYN_struct of adder_sub_N32 is

   component cla_adder_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component generic_xor_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal B_in_31_port, B_in_30_port, B_in_29_port, B_in_28_port, B_in_27_port,
      B_in_26_port, B_in_25_port, B_in_24_port, B_in_23_port, B_in_22_port, 
      B_in_21_port, B_in_20_port, B_in_19_port, B_in_18_port, B_in_17_port, 
      B_in_16_port, B_in_15_port, B_in_14_port, B_in_13_port, B_in_12_port, 
      B_in_11_port, B_in_10_port, B_in_9_port, B_in_8_port, B_in_7_port, 
      B_in_6_port, B_in_5_port, B_in_4_port, B_in_3_port, B_in_2_port, 
      B_in_1_port, B_in_0_port : std_logic;

begin
   
   xor_g : generic_xor_N32 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => Ci, Y(31) => B_in_31_port, Y(30) => 
                           B_in_30_port, Y(29) => B_in_29_port, Y(28) => 
                           B_in_28_port, Y(27) => B_in_27_port, Y(26) => 
                           B_in_26_port, Y(25) => B_in_25_port, Y(24) => 
                           B_in_24_port, Y(23) => B_in_23_port, Y(22) => 
                           B_in_22_port, Y(21) => B_in_21_port, Y(20) => 
                           B_in_20_port, Y(19) => B_in_19_port, Y(18) => 
                           B_in_18_port, Y(17) => B_in_17_port, Y(16) => 
                           B_in_16_port, Y(15) => B_in_15_port, Y(14) => 
                           B_in_14_port, Y(13) => B_in_13_port, Y(12) => 
                           B_in_12_port, Y(11) => B_in_11_port, Y(10) => 
                           B_in_10_port, Y(9) => B_in_9_port, Y(8) => 
                           B_in_8_port, Y(7) => B_in_7_port, Y(6) => 
                           B_in_6_port, Y(5) => B_in_5_port, Y(4) => 
                           B_in_4_port, Y(3) => B_in_3_port, Y(2) => 
                           B_in_2_port, Y(1) => B_in_1_port, Y(0) => 
                           B_in_0_port);
   add : cla_adder_N32_0 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B_in_31_port, B(30) => 
                           B_in_30_port, B(29) => B_in_29_port, B(28) => 
                           B_in_28_port, B(27) => B_in_27_port, B(26) => 
                           B_in_26_port, B(25) => B_in_25_port, B(24) => 
                           B_in_24_port, B(23) => B_in_23_port, B(22) => 
                           B_in_22_port, B(21) => B_in_21_port, B(20) => 
                           B_in_20_port, B(19) => B_in_19_port, B(18) => 
                           B_in_18_port, B(17) => B_in_17_port, B(16) => 
                           B_in_16_port, B(15) => B_in_15_port, B(14) => 
                           B_in_14_port, B(13) => B_in_13_port, B(12) => 
                           B_in_12_port, B(11) => B_in_11_port, B(10) => 
                           B_in_10_port, B(9) => B_in_9_port, B(8) => 
                           B_in_8_port, B(7) => B_in_7_port, B(6) => 
                           B_in_6_port, B(5) => B_in_5_port, B(4) => 
                           B_in_4_port, B(3) => B_in_3_port, B(2) => 
                           B_in_2_port, B(1) => B_in_1_port, B(0) => 
                           B_in_0_port, Ci => Ci, Cout => Cout, Sum(31) => 
                           Sum(31), Sum(30) => Sum(30), Sum(29) => Sum(29), 
                           Sum(28) => Sum(28), Sum(27) => Sum(27), Sum(26) => 
                           Sum(26), Sum(25) => Sum(25), Sum(24) => Sum(24), 
                           Sum(23) => Sum(23), Sum(22) => Sum(22), Sum(21) => 
                           Sum(21), Sum(20) => Sum(20), Sum(19) => Sum(19), 
                           Sum(18) => Sum(18), Sum(17) => Sum(17), Sum(16) => 
                           Sum(16), Sum(15) => Sum(15), Sum(14) => Sum(14), 
                           Sum(13) => Sum(13), Sum(12) => Sum(12), Sum(11) => 
                           Sum(11), Sum(10) => Sum(10), Sum(9) => Sum(9), 
                           Sum(8) => Sum(8), Sum(7) => Sum(7), Sum(6) => Sum(6)
                           , Sum(5) => Sum(5), Sum(4) => Sum(4), Sum(3) => 
                           Sum(3), Sum(2) => Sum(2), Sum(1) => Sum(1), Sum(0) 
                           => Sum(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_alu.all;

entity alu is

   port( A, B : in bus32;  OP : in aluOp;  Y1 : out bus32;  cout : out 
         std_logic);

end alu;

architecture SYN_behav of alu is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component mux_alu
      port( addsub, mul, log, shift, lhi : in std_logic_vector (31 downto 0);  
            gt, get, lt, let, eq, neq : in std_logic;  sel : in 
            std_logic_vector (0 to 4);  out_mux : out std_logic_vector (31 
            downto 0));
   end component;
   
   component comparator
      port( C : in std_logic;  Sum : in std_logic_vector (31 downto 0);  sign :
            in std_logic;  gt, get, lt, let, eq, neq : out std_logic);
   end component;
   
   component shifter
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  C : out std_logic_vector (31 downto
            0));
   end component;
   
   component logical
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (3 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component booth_mul_N16
      port( A, B : in std_logic_vector (15 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component adder_sub_N32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Cout
            : out std_logic;  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, OP_4_port, OP_3_port, OP_2_port, OP_1_port, OP_0_port,
      cout_port, add_sub, A_add_31_port, A_add_30_port, A_add_29_port, 
      A_add_28_port, A_add_27_port, A_add_26_port, A_add_25_port, A_add_24_port
      , A_add_23_port, A_add_22_port, A_add_21_port, A_add_20_port, 
      A_add_19_port, A_add_18_port, A_add_17_port, A_add_16_port, A_add_15_port
      , A_add_14_port, A_add_13_port, A_add_12_port, A_add_11_port, 
      A_add_10_port, A_add_9_port, A_add_8_port, A_add_7_port, A_add_6_port, 
      A_add_5_port, A_add_4_port, A_add_3_port, A_add_2_port, A_add_1_port, 
      A_add_0_port, B_add_31_port, B_add_30_port, B_add_29_port, B_add_28_port,
      B_add_27_port, B_add_26_port, B_add_25_port, B_add_24_port, B_add_23_port
      , B_add_22_port, B_add_21_port, B_add_20_port, B_add_19_port, 
      B_add_18_port, B_add_17_port, B_add_16_port, B_add_15_port, B_add_14_port
      , B_add_13_port, B_add_12_port, B_add_11_port, B_add_10_port, 
      B_add_9_port, B_add_8_port, B_add_7_port, B_add_6_port, B_add_5_port, 
      B_add_4_port, B_add_3_port, B_add_2_port, B_add_1_port, B_add_0_port, 
      A_mul_15_port, A_mul_14_port, A_mul_13_port, A_mul_12_port, A_mul_11_port
      , A_mul_10_port, A_mul_9_port, A_mul_8_port, A_mul_7_port, A_mul_6_port, 
      A_mul_5_port, A_mul_4_port, A_mul_3_port, A_mul_2_port, A_mul_1_port, 
      B_mul_15_port, B_mul_14_port, B_mul_13_port, B_mul_12_port, B_mul_11_port
      , B_mul_10_port, B_mul_9_port, B_mul_8_port, B_mul_7_port, B_mul_6_port, 
      B_mul_5_port, B_mul_4_port, B_mul_3_port, B_mul_2_port, B_mul_1_port, 
      B_mul_0_port, sel_log_3_port, sel_log_2_port, sel_log_1_port, 
      sel_log_0_port, A_log_31_port, A_log_30_port, A_log_29_port, 
      A_log_28_port, A_log_27_port, A_log_26_port, A_log_25_port, A_log_24_port
      , A_log_23_port, A_log_22_port, A_log_21_port, A_log_20_port, 
      A_log_19_port, A_log_18_port, A_log_17_port, A_log_16_port, A_log_15_port
      , A_log_14_port, A_log_13_port, A_log_12_port, A_log_11_port, 
      A_log_10_port, A_log_9_port, A_log_8_port, A_log_7_port, A_log_6_port, 
      A_log_5_port, A_log_4_port, A_log_3_port, A_log_2_port, A_log_1_port, 
      A_log_0_port, B_log_31_port, B_log_30_port, B_log_29_port, B_log_28_port,
      B_log_27_port, B_log_26_port, B_log_25_port, B_log_24_port, B_log_23_port
      , B_log_22_port, B_log_21_port, B_log_20_port, B_log_19_port, 
      B_log_18_port, B_log_17_port, B_log_16_port, B_log_15_port, B_log_14_port
      , B_log_13_port, B_log_12_port, B_log_11_port, B_log_10_port, 
      B_log_9_port, B_log_8_port, B_log_7_port, B_log_6_port, B_log_5_port, 
      B_log_4_port, B_log_3_port, B_log_2_port, B_log_1_port, B_log_0_port, 
      sel_shift_1_port, sel_shift_0_port, A_sht_31_port, A_sht_30_port, 
      A_sht_29_port, A_sht_28_port, A_sht_27_port, A_sht_26_port, A_sht_25_port
      , A_sht_24_port, A_sht_23_port, A_sht_22_port, A_sht_21_port, 
      A_sht_20_port, A_sht_19_port, A_sht_18_port, A_sht_17_port, A_sht_16_port
      , A_sht_15_port, A_sht_14_port, A_sht_13_port, A_sht_12_port, 
      A_sht_11_port, A_sht_10_port, A_sht_9_port, A_sht_8_port, A_sht_7_port, 
      A_sht_6_port, A_sht_5_port, A_sht_4_port, A_sht_3_port, A_sht_2_port, 
      A_sht_1_port, A_sht_0_port, B_sht_31_port, B_sht_30_port, B_sht_29_port, 
      B_sht_28_port, B_sht_27_port, B_sht_26_port, B_sht_25_port, B_sht_24_port
      , B_sht_23_port, B_sht_22_port, B_sht_21_port, B_sht_20_port, 
      B_sht_19_port, B_sht_18_port, B_sht_17_port, B_sht_16_port, B_sht_15_port
      , B_sht_14_port, B_sht_13_port, B_sht_12_port, B_sht_11_port, 
      B_sht_10_port, B_sht_9_port, B_sht_8_port, B_sht_7_port, B_sht_6_port, 
      B_sht_5_port, B_sht_4_port, B_sht_3_port, B_sht_2_port, B_sht_1_port, 
      B_sht_0_port, sign, B_lhi_15_port, B_lhi_14_port, B_lhi_13_port, 
      B_lhi_12_port, B_lhi_11_port, B_lhi_10_port, B_lhi_9_port, B_lhi_8_port, 
      B_lhi_7_port, B_lhi_6_port, B_lhi_5_port, B_lhi_4_port, B_lhi_3_port, 
      B_lhi_2_port, B_lhi_1_port, B_lhi_0_port, N25, N26, N27, N28, N29, N31, 
      N32, N33, N34, N35, N36, out_add_31_port, out_add_30_port, 
      out_add_29_port, out_add_28_port, out_add_27_port, out_add_26_port, 
      out_add_25_port, out_add_24_port, out_add_23_port, out_add_22_port, 
      out_add_21_port, out_add_20_port, out_add_19_port, out_add_18_port, 
      out_add_17_port, out_add_16_port, out_add_15_port, out_add_14_port, 
      out_add_13_port, out_add_12_port, out_add_11_port, out_add_10_port, 
      out_add_9_port, out_add_8_port, out_add_7_port, out_add_6_port, 
      out_add_5_port, out_add_4_port, out_add_3_port, out_add_2_port, 
      out_add_1_port, out_add_0_port, out_mul_31_port, out_mul_30_port, 
      out_mul_29_port, out_mul_28_port, out_mul_27_port, out_mul_26_port, 
      out_mul_25_port, out_mul_24_port, out_mul_23_port, out_mul_22_port, 
      out_mul_21_port, out_mul_20_port, out_mul_19_port, out_mul_18_port, 
      out_mul_17_port, out_mul_16_port, out_mul_15_port, out_mul_14_port, 
      out_mul_13_port, out_mul_12_port, out_mul_11_port, out_mul_10_port, 
      out_mul_9_port, out_mul_8_port, out_mul_7_port, out_mul_6_port, 
      out_mul_5_port, out_mul_4_port, out_mul_3_port, out_mul_2_port, 
      out_mul_1_port, out_mul_0_port, out_log_31_port, out_log_30_port, 
      out_log_29_port, out_log_28_port, out_log_27_port, out_log_26_port, 
      out_log_25_port, out_log_24_port, out_log_23_port, out_log_22_port, 
      out_log_21_port, out_log_20_port, out_log_19_port, out_log_18_port, 
      out_log_17_port, out_log_16_port, out_log_15_port, out_log_14_port, 
      out_log_13_port, out_log_12_port, out_log_11_port, out_log_10_port, 
      out_log_9_port, out_log_8_port, out_log_7_port, out_log_6_port, 
      out_log_5_port, out_log_4_port, out_log_3_port, out_log_2_port, 
      out_log_1_port, out_log_0_port, out_shift_31_port, out_shift_30_port, 
      out_shift_29_port, out_shift_28_port, out_shift_27_port, 
      out_shift_26_port, out_shift_25_port, out_shift_24_port, 
      out_shift_23_port, out_shift_22_port, out_shift_21_port, 
      out_shift_20_port, out_shift_19_port, out_shift_18_port, 
      out_shift_17_port, out_shift_16_port, out_shift_15_port, 
      out_shift_14_port, out_shift_13_port, out_shift_12_port, 
      out_shift_11_port, out_shift_10_port, out_shift_9_port, out_shift_8_port,
      out_shift_7_port, out_shift_6_port, out_shift_5_port, out_shift_4_port, 
      out_shift_3_port, out_shift_2_port, out_shift_1_port, out_shift_0_port, 
      gt, get, lt, let, eq, neq, n23, n24, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98 : std_logic;

begin
   (OP_4_port, OP_3_port, OP_2_port, OP_1_port, OP_0_port) <= 
      aluOp_to_std_logic_vector(OP);
   cout <= cout_port;
   
   adder_subtr : adder_sub_N32 port map( A(31) => A_add_31_port, A(30) => 
                           A_add_30_port, A(29) => A_add_29_port, A(28) => 
                           A_add_28_port, A(27) => A_add_27_port, A(26) => 
                           A_add_26_port, A(25) => A_add_25_port, A(24) => 
                           A_add_24_port, A(23) => A_add_23_port, A(22) => 
                           A_add_22_port, A(21) => A_add_21_port, A(20) => 
                           A_add_20_port, A(19) => A_add_19_port, A(18) => 
                           A_add_18_port, A(17) => A_add_17_port, A(16) => 
                           A_add_16_port, A(15) => A_add_15_port, A(14) => 
                           A_add_14_port, A(13) => A_add_13_port, A(12) => 
                           A_add_12_port, A(11) => A_add_11_port, A(10) => 
                           A_add_10_port, A(9) => A_add_9_port, A(8) => 
                           A_add_8_port, A(7) => A_add_7_port, A(6) => 
                           A_add_6_port, A(5) => A_add_5_port, A(4) => 
                           A_add_4_port, A(3) => A_add_3_port, A(2) => 
                           A_add_2_port, A(1) => A_add_1_port, A(0) => 
                           A_add_0_port, B(31) => B_add_31_port, B(30) => 
                           B_add_30_port, B(29) => B_add_29_port, B(28) => 
                           B_add_28_port, B(27) => B_add_27_port, B(26) => 
                           B_add_26_port, B(25) => B_add_25_port, B(24) => 
                           B_add_24_port, B(23) => B_add_23_port, B(22) => 
                           B_add_22_port, B(21) => B_add_21_port, B(20) => 
                           B_add_20_port, B(19) => B_add_19_port, B(18) => 
                           B_add_18_port, B(17) => B_add_17_port, B(16) => 
                           B_add_16_port, B(15) => B_add_15_port, B(14) => 
                           B_add_14_port, B(13) => B_add_13_port, B(12) => 
                           B_add_12_port, B(11) => B_add_11_port, B(10) => 
                           B_add_10_port, B(9) => B_add_9_port, B(8) => 
                           B_add_8_port, B(7) => B_add_7_port, B(6) => 
                           B_add_6_port, B(5) => B_add_5_port, B(4) => 
                           B_add_4_port, B(3) => B_add_3_port, B(2) => 
                           B_add_2_port, B(1) => B_add_1_port, B(0) => 
                           B_add_0_port, Ci => add_sub, Cout => cout_port, 
                           Sum(31) => out_add_31_port, Sum(30) => 
                           out_add_30_port, Sum(29) => out_add_29_port, Sum(28)
                           => out_add_28_port, Sum(27) => out_add_27_port, 
                           Sum(26) => out_add_26_port, Sum(25) => 
                           out_add_25_port, Sum(24) => out_add_24_port, Sum(23)
                           => out_add_23_port, Sum(22) => out_add_22_port, 
                           Sum(21) => out_add_21_port, Sum(20) => 
                           out_add_20_port, Sum(19) => out_add_19_port, Sum(18)
                           => out_add_18_port, Sum(17) => out_add_17_port, 
                           Sum(16) => out_add_16_port, Sum(15) => 
                           out_add_15_port, Sum(14) => out_add_14_port, Sum(13)
                           => out_add_13_port, Sum(12) => out_add_12_port, 
                           Sum(11) => out_add_11_port, Sum(10) => 
                           out_add_10_port, Sum(9) => out_add_9_port, Sum(8) =>
                           out_add_8_port, Sum(7) => out_add_7_port, Sum(6) => 
                           out_add_6_port, Sum(5) => out_add_5_port, Sum(4) => 
                           out_add_4_port, Sum(3) => out_add_3_port, Sum(2) => 
                           out_add_2_port, Sum(1) => out_add_1_port, Sum(0) => 
                           out_add_0_port);
   mul : booth_mul_N16 port map( A(15) => A_mul_15_port, A(14) => A_mul_14_port
                           , A(13) => A_mul_13_port, A(12) => A_mul_12_port, 
                           A(11) => A_mul_11_port, A(10) => A_mul_10_port, A(9)
                           => A_mul_9_port, A(8) => A_mul_8_port, A(7) => 
                           A_mul_7_port, A(6) => A_mul_6_port, A(5) => 
                           A_mul_5_port, A(4) => A_mul_4_port, A(3) => 
                           A_mul_3_port, A(2) => A_mul_2_port, A(1) => 
                           A_mul_1_port, A(0) => n23, B(15) => B_mul_15_port, 
                           B(14) => B_mul_14_port, B(13) => B_mul_13_port, 
                           B(12) => B_mul_12_port, B(11) => B_mul_11_port, 
                           B(10) => B_mul_10_port, B(9) => B_mul_9_port, B(8) 
                           => B_mul_8_port, B(7) => B_mul_7_port, B(6) => 
                           B_mul_6_port, B(5) => B_mul_5_port, B(4) => 
                           B_mul_4_port, B(3) => B_mul_3_port, B(2) => 
                           B_mul_2_port, B(1) => B_mul_1_port, B(0) => 
                           B_mul_0_port, Y(31) => out_mul_31_port, Y(30) => 
                           out_mul_30_port, Y(29) => out_mul_29_port, Y(28) => 
                           out_mul_28_port, Y(27) => out_mul_27_port, Y(26) => 
                           out_mul_26_port, Y(25) => out_mul_25_port, Y(24) => 
                           out_mul_24_port, Y(23) => out_mul_23_port, Y(22) => 
                           out_mul_22_port, Y(21) => out_mul_21_port, Y(20) => 
                           out_mul_20_port, Y(19) => out_mul_19_port, Y(18) => 
                           out_mul_18_port, Y(17) => out_mul_17_port, Y(16) => 
                           out_mul_16_port, Y(15) => out_mul_15_port, Y(14) => 
                           out_mul_14_port, Y(13) => out_mul_13_port, Y(12) => 
                           out_mul_12_port, Y(11) => out_mul_11_port, Y(10) => 
                           out_mul_10_port, Y(9) => out_mul_9_port, Y(8) => 
                           out_mul_8_port, Y(7) => out_mul_7_port, Y(6) => 
                           out_mul_6_port, Y(5) => out_mul_5_port, Y(4) => 
                           out_mul_4_port, Y(3) => out_mul_3_port, Y(2) => 
                           out_mul_2_port, Y(1) => out_mul_1_port, Y(0) => 
                           out_mul_0_port);
   logic : logical port map( A(31) => A_log_31_port, A(30) => A_log_30_port, 
                           A(29) => A_log_29_port, A(28) => A_log_28_port, 
                           A(27) => A_log_27_port, A(26) => A_log_26_port, 
                           A(25) => A_log_25_port, A(24) => A_log_24_port, 
                           A(23) => A_log_23_port, A(22) => A_log_22_port, 
                           A(21) => A_log_21_port, A(20) => A_log_20_port, 
                           A(19) => A_log_19_port, A(18) => A_log_18_port, 
                           A(17) => A_log_17_port, A(16) => A_log_16_port, 
                           A(15) => A_log_15_port, A(14) => A_log_14_port, 
                           A(13) => A_log_13_port, A(12) => A_log_12_port, 
                           A(11) => A_log_11_port, A(10) => A_log_10_port, A(9)
                           => A_log_9_port, A(8) => A_log_8_port, A(7) => 
                           A_log_7_port, A(6) => A_log_6_port, A(5) => 
                           A_log_5_port, A(4) => A_log_4_port, A(3) => 
                           A_log_3_port, A(2) => A_log_2_port, A(1) => 
                           A_log_1_port, A(0) => A_log_0_port, B(31) => 
                           B_log_31_port, B(30) => B_log_30_port, B(29) => 
                           B_log_29_port, B(28) => B_log_28_port, B(27) => 
                           B_log_27_port, B(26) => B_log_26_port, B(25) => 
                           B_log_25_port, B(24) => B_log_24_port, B(23) => 
                           B_log_23_port, B(22) => B_log_22_port, B(21) => 
                           B_log_21_port, B(20) => B_log_20_port, B(19) => 
                           B_log_19_port, B(18) => B_log_18_port, B(17) => 
                           B_log_17_port, B(16) => B_log_16_port, B(15) => 
                           B_log_15_port, B(14) => B_log_14_port, B(13) => 
                           B_log_13_port, B(12) => B_log_12_port, B(11) => 
                           B_log_11_port, B(10) => B_log_10_port, B(9) => 
                           B_log_9_port, B(8) => B_log_8_port, B(7) => 
                           B_log_7_port, B(6) => B_log_6_port, B(5) => 
                           B_log_5_port, B(4) => B_log_4_port, B(3) => 
                           B_log_3_port, B(2) => B_log_2_port, B(1) => 
                           B_log_1_port, B(0) => B_log_0_port, sel(3) => 
                           sel_log_3_port, sel(2) => sel_log_2_port, sel(1) => 
                           sel_log_1_port, sel(0) => sel_log_0_port, Y(31) => 
                           out_log_31_port, Y(30) => out_log_30_port, Y(29) => 
                           out_log_29_port, Y(28) => out_log_28_port, Y(27) => 
                           out_log_27_port, Y(26) => out_log_26_port, Y(25) => 
                           out_log_25_port, Y(24) => out_log_24_port, Y(23) => 
                           out_log_23_port, Y(22) => out_log_22_port, Y(21) => 
                           out_log_21_port, Y(20) => out_log_20_port, Y(19) => 
                           out_log_19_port, Y(18) => out_log_18_port, Y(17) => 
                           out_log_17_port, Y(16) => out_log_16_port, Y(15) => 
                           out_log_15_port, Y(14) => out_log_14_port, Y(13) => 
                           out_log_13_port, Y(12) => out_log_12_port, Y(11) => 
                           out_log_11_port, Y(10) => out_log_10_port, Y(9) => 
                           out_log_9_port, Y(8) => out_log_8_port, Y(7) => 
                           out_log_7_port, Y(6) => out_log_6_port, Y(5) => 
                           out_log_5_port, Y(4) => out_log_4_port, Y(3) => 
                           out_log_3_port, Y(2) => out_log_2_port, Y(1) => 
                           out_log_1_port, Y(0) => out_log_0_port);
   shift : shifter port map( A(31) => A_sht_31_port, A(30) => A_sht_30_port, 
                           A(29) => A_sht_29_port, A(28) => A_sht_28_port, 
                           A(27) => A_sht_27_port, A(26) => A_sht_26_port, 
                           A(25) => A_sht_25_port, A(24) => A_sht_24_port, 
                           A(23) => A_sht_23_port, A(22) => A_sht_22_port, 
                           A(21) => A_sht_21_port, A(20) => A_sht_20_port, 
                           A(19) => A_sht_19_port, A(18) => A_sht_18_port, 
                           A(17) => A_sht_17_port, A(16) => A_sht_16_port, 
                           A(15) => A_sht_15_port, A(14) => A_sht_14_port, 
                           A(13) => A_sht_13_port, A(12) => A_sht_12_port, 
                           A(11) => A_sht_11_port, A(10) => A_sht_10_port, A(9)
                           => A_sht_9_port, A(8) => A_sht_8_port, A(7) => 
                           A_sht_7_port, A(6) => A_sht_6_port, A(5) => 
                           A_sht_5_port, A(4) => A_sht_4_port, A(3) => 
                           A_sht_3_port, A(2) => A_sht_2_port, A(1) => 
                           A_sht_1_port, A(0) => A_sht_0_port, B(31) => 
                           B_sht_31_port, B(30) => B_sht_30_port, B(29) => 
                           B_sht_29_port, B(28) => B_sht_28_port, B(27) => 
                           B_sht_27_port, B(26) => B_sht_26_port, B(25) => 
                           B_sht_25_port, B(24) => B_sht_24_port, B(23) => 
                           B_sht_23_port, B(22) => B_sht_22_port, B(21) => 
                           B_sht_21_port, B(20) => B_sht_20_port, B(19) => 
                           B_sht_19_port, B(18) => B_sht_18_port, B(17) => 
                           B_sht_17_port, B(16) => B_sht_16_port, B(15) => 
                           B_sht_15_port, B(14) => B_sht_14_port, B(13) => 
                           B_sht_13_port, B(12) => B_sht_12_port, B(11) => 
                           B_sht_11_port, B(10) => B_sht_10_port, B(9) => 
                           B_sht_9_port, B(8) => B_sht_8_port, B(7) => 
                           B_sht_7_port, B(6) => B_sht_6_port, B(5) => 
                           B_sht_5_port, B(4) => B_sht_4_port, B(3) => 
                           B_sht_3_port, B(2) => B_sht_2_port, B(1) => 
                           B_sht_1_port, B(0) => B_sht_0_port, sel(1) => 
                           sel_shift_1_port, sel(0) => sel_shift_0_port, C(31) 
                           => out_shift_31_port, C(30) => out_shift_30_port, 
                           C(29) => out_shift_29_port, C(28) => 
                           out_shift_28_port, C(27) => out_shift_27_port, C(26)
                           => out_shift_26_port, C(25) => out_shift_25_port, 
                           C(24) => out_shift_24_port, C(23) => 
                           out_shift_23_port, C(22) => out_shift_22_port, C(21)
                           => out_shift_21_port, C(20) => out_shift_20_port, 
                           C(19) => out_shift_19_port, C(18) => 
                           out_shift_18_port, C(17) => out_shift_17_port, C(16)
                           => out_shift_16_port, C(15) => out_shift_15_port, 
                           C(14) => out_shift_14_port, C(13) => 
                           out_shift_13_port, C(12) => out_shift_12_port, C(11)
                           => out_shift_11_port, C(10) => out_shift_10_port, 
                           C(9) => out_shift_9_port, C(8) => out_shift_8_port, 
                           C(7) => out_shift_7_port, C(6) => out_shift_6_port, 
                           C(5) => out_shift_5_port, C(4) => out_shift_4_port, 
                           C(3) => out_shift_3_port, C(2) => out_shift_2_port, 
                           C(1) => out_shift_1_port, C(0) => out_shift_0_port);
   compar : comparator port map( C => cout_port, Sum(31) => out_add_31_port, 
                           Sum(30) => out_add_30_port, Sum(29) => 
                           out_add_29_port, Sum(28) => out_add_28_port, Sum(27)
                           => out_add_27_port, Sum(26) => out_add_26_port, 
                           Sum(25) => out_add_25_port, Sum(24) => 
                           out_add_24_port, Sum(23) => out_add_23_port, Sum(22)
                           => out_add_22_port, Sum(21) => out_add_21_port, 
                           Sum(20) => out_add_20_port, Sum(19) => 
                           out_add_19_port, Sum(18) => out_add_18_port, Sum(17)
                           => out_add_17_port, Sum(16) => out_add_16_port, 
                           Sum(15) => out_add_15_port, Sum(14) => 
                           out_add_14_port, Sum(13) => out_add_13_port, Sum(12)
                           => out_add_12_port, Sum(11) => out_add_11_port, 
                           Sum(10) => out_add_10_port, Sum(9) => out_add_9_port
                           , Sum(8) => out_add_8_port, Sum(7) => out_add_7_port
                           , Sum(6) => out_add_6_port, Sum(5) => out_add_5_port
                           , Sum(4) => out_add_4_port, Sum(3) => out_add_3_port
                           , Sum(2) => out_add_2_port, Sum(1) => out_add_1_port
                           , Sum(0) => out_add_0_port, sign => sign, gt => gt, 
                           get => get, lt => lt, let => let, eq => eq, neq => 
                           neq);
   muxy1 : mux_alu port map( addsub(31) => out_add_31_port, addsub(30) => 
                           out_add_30_port, addsub(29) => out_add_29_port, 
                           addsub(28) => out_add_28_port, addsub(27) => 
                           out_add_27_port, addsub(26) => out_add_26_port, 
                           addsub(25) => out_add_25_port, addsub(24) => 
                           out_add_24_port, addsub(23) => out_add_23_port, 
                           addsub(22) => out_add_22_port, addsub(21) => 
                           out_add_21_port, addsub(20) => out_add_20_port, 
                           addsub(19) => out_add_19_port, addsub(18) => 
                           out_add_18_port, addsub(17) => out_add_17_port, 
                           addsub(16) => out_add_16_port, addsub(15) => 
                           out_add_15_port, addsub(14) => out_add_14_port, 
                           addsub(13) => out_add_13_port, addsub(12) => 
                           out_add_12_port, addsub(11) => out_add_11_port, 
                           addsub(10) => out_add_10_port, addsub(9) => 
                           out_add_9_port, addsub(8) => out_add_8_port, 
                           addsub(7) => out_add_7_port, addsub(6) => 
                           out_add_6_port, addsub(5) => out_add_5_port, 
                           addsub(4) => out_add_4_port, addsub(3) => 
                           out_add_3_port, addsub(2) => out_add_2_port, 
                           addsub(1) => out_add_1_port, addsub(0) => 
                           out_add_0_port, mul(31) => out_mul_31_port, mul(30) 
                           => out_mul_30_port, mul(29) => out_mul_29_port, 
                           mul(28) => out_mul_28_port, mul(27) => 
                           out_mul_27_port, mul(26) => out_mul_26_port, mul(25)
                           => out_mul_25_port, mul(24) => out_mul_24_port, 
                           mul(23) => out_mul_23_port, mul(22) => 
                           out_mul_22_port, mul(21) => out_mul_21_port, mul(20)
                           => out_mul_20_port, mul(19) => out_mul_19_port, 
                           mul(18) => out_mul_18_port, mul(17) => 
                           out_mul_17_port, mul(16) => out_mul_16_port, mul(15)
                           => out_mul_15_port, mul(14) => out_mul_14_port, 
                           mul(13) => out_mul_13_port, mul(12) => 
                           out_mul_12_port, mul(11) => out_mul_11_port, mul(10)
                           => out_mul_10_port, mul(9) => out_mul_9_port, mul(8)
                           => out_mul_8_port, mul(7) => out_mul_7_port, mul(6) 
                           => out_mul_6_port, mul(5) => out_mul_5_port, mul(4) 
                           => out_mul_4_port, mul(3) => out_mul_3_port, mul(2) 
                           => out_mul_2_port, mul(1) => out_mul_1_port, mul(0) 
                           => out_mul_0_port, log(31) => out_log_31_port, 
                           log(30) => out_log_30_port, log(29) => 
                           out_log_29_port, log(28) => out_log_28_port, log(27)
                           => out_log_27_port, log(26) => out_log_26_port, 
                           log(25) => out_log_25_port, log(24) => 
                           out_log_24_port, log(23) => out_log_23_port, log(22)
                           => out_log_22_port, log(21) => out_log_21_port, 
                           log(20) => out_log_20_port, log(19) => 
                           out_log_19_port, log(18) => out_log_18_port, log(17)
                           => out_log_17_port, log(16) => out_log_16_port, 
                           log(15) => out_log_15_port, log(14) => 
                           out_log_14_port, log(13) => out_log_13_port, log(12)
                           => out_log_12_port, log(11) => out_log_11_port, 
                           log(10) => out_log_10_port, log(9) => out_log_9_port
                           , log(8) => out_log_8_port, log(7) => out_log_7_port
                           , log(6) => out_log_6_port, log(5) => out_log_5_port
                           , log(4) => out_log_4_port, log(3) => out_log_3_port
                           , log(2) => out_log_2_port, log(1) => out_log_1_port
                           , log(0) => out_log_0_port, shift(31) => 
                           out_shift_31_port, shift(30) => out_shift_30_port, 
                           shift(29) => out_shift_29_port, shift(28) => 
                           out_shift_28_port, shift(27) => out_shift_27_port, 
                           shift(26) => out_shift_26_port, shift(25) => 
                           out_shift_25_port, shift(24) => out_shift_24_port, 
                           shift(23) => out_shift_23_port, shift(22) => 
                           out_shift_22_port, shift(21) => out_shift_21_port, 
                           shift(20) => out_shift_20_port, shift(19) => 
                           out_shift_19_port, shift(18) => out_shift_18_port, 
                           shift(17) => out_shift_17_port, shift(16) => 
                           out_shift_16_port, shift(15) => out_shift_15_port, 
                           shift(14) => out_shift_14_port, shift(13) => 
                           out_shift_13_port, shift(12) => out_shift_12_port, 
                           shift(11) => out_shift_11_port, shift(10) => 
                           out_shift_10_port, shift(9) => out_shift_9_port, 
                           shift(8) => out_shift_8_port, shift(7) => 
                           out_shift_7_port, shift(6) => out_shift_6_port, 
                           shift(5) => out_shift_5_port, shift(4) => 
                           out_shift_4_port, shift(3) => out_shift_3_port, 
                           shift(2) => out_shift_2_port, shift(1) => 
                           out_shift_1_port, shift(0) => out_shift_0_port, 
                           lhi(31) => B_lhi_15_port, lhi(30) => B_lhi_14_port, 
                           lhi(29) => B_lhi_13_port, lhi(28) => B_lhi_12_port, 
                           lhi(27) => B_lhi_11_port, lhi(26) => B_lhi_10_port, 
                           lhi(25) => B_lhi_9_port, lhi(24) => B_lhi_8_port, 
                           lhi(23) => B_lhi_7_port, lhi(22) => B_lhi_6_port, 
                           lhi(21) => B_lhi_5_port, lhi(20) => B_lhi_4_port, 
                           lhi(19) => B_lhi_3_port, lhi(18) => B_lhi_2_port, 
                           lhi(17) => B_lhi_1_port, lhi(16) => B_lhi_0_port, 
                           lhi(15) => X_Logic0_port, lhi(14) => X_Logic0_port, 
                           lhi(13) => X_Logic0_port, lhi(12) => X_Logic0_port, 
                           lhi(11) => X_Logic0_port, lhi(10) => X_Logic0_port, 
                           lhi(9) => X_Logic0_port, lhi(8) => X_Logic0_port, 
                           lhi(7) => X_Logic0_port, lhi(6) => X_Logic0_port, 
                           lhi(5) => X_Logic0_port, lhi(4) => X_Logic0_port, 
                           lhi(3) => X_Logic0_port, lhi(2) => X_Logic0_port, 
                           lhi(1) => X_Logic0_port, lhi(0) => X_Logic0_port, gt
                           => gt, get => get, lt => lt, let => let, eq => eq, 
                           neq => neq, sel(0) => OP_4_port, sel(1) => OP_3_port
                           , sel(2) => OP_2_port, sel(3) => OP_1_port, sel(4) 
                           => OP_0_port, out_mux(31) => Y1(31), out_mux(30) => 
                           Y1(30), out_mux(29) => Y1(29), out_mux(28) => Y1(28)
                           , out_mux(27) => Y1(27), out_mux(26) => Y1(26), 
                           out_mux(25) => Y1(25), out_mux(24) => Y1(24), 
                           out_mux(23) => Y1(23), out_mux(22) => Y1(22), 
                           out_mux(21) => Y1(21), out_mux(20) => Y1(20), 
                           out_mux(19) => Y1(19), out_mux(18) => Y1(18), 
                           out_mux(17) => Y1(17), out_mux(16) => Y1(16), 
                           out_mux(15) => Y1(15), out_mux(14) => Y1(14), 
                           out_mux(13) => Y1(13), out_mux(12) => Y1(12), 
                           out_mux(11) => Y1(11), out_mux(10) => Y1(10), 
                           out_mux(9) => Y1(9), out_mux(8) => Y1(8), out_mux(7)
                           => Y1(7), out_mux(6) => Y1(6), out_mux(5) => Y1(5), 
                           out_mux(4) => Y1(4), out_mux(3) => Y1(3), out_mux(2)
                           => Y1(2), out_mux(1) => Y1(1), out_mux(0) => Y1(0));
   X_Logic0_port <= '0';
   B_lhi_reg_15_inst : DLH_X1 port map( G => N36, D => B(15), Q => 
                           B_lhi_15_port);
   B_lhi_reg_14_inst : DLH_X1 port map( G => N36, D => B(14), Q => 
                           B_lhi_14_port);
   B_lhi_reg_13_inst : DLH_X1 port map( G => N36, D => B(13), Q => 
                           B_lhi_13_port);
   B_lhi_reg_12_inst : DLH_X1 port map( G => N36, D => B(12), Q => 
                           B_lhi_12_port);
   B_lhi_reg_11_inst : DLH_X1 port map( G => N36, D => B(11), Q => 
                           B_lhi_11_port);
   B_lhi_reg_10_inst : DLH_X1 port map( G => N36, D => B(10), Q => 
                           B_lhi_10_port);
   B_lhi_reg_9_inst : DLH_X1 port map( G => N36, D => B(9), Q => B_lhi_9_port);
   B_lhi_reg_8_inst : DLH_X1 port map( G => N36, D => B(8), Q => B_lhi_8_port);
   B_lhi_reg_7_inst : DLH_X1 port map( G => N36, D => B(7), Q => B_lhi_7_port);
   B_lhi_reg_6_inst : DLH_X1 port map( G => N36, D => B(6), Q => B_lhi_6_port);
   B_lhi_reg_5_inst : DLH_X1 port map( G => N36, D => B(5), Q => B_lhi_5_port);
   B_lhi_reg_4_inst : DLH_X1 port map( G => N36, D => B(4), Q => B_lhi_4_port);
   B_lhi_reg_3_inst : DLH_X1 port map( G => N36, D => B(3), Q => B_lhi_3_port);
   B_lhi_reg_2_inst : DLH_X1 port map( G => N36, D => B(2), Q => B_lhi_2_port);
   B_lhi_reg_1_inst : DLH_X1 port map( G => N36, D => B(1), Q => B_lhi_1_port);
   B_lhi_reg_0_inst : DLH_X1 port map( G => N36, D => B(0), Q => B_lhi_0_port);
   A_add_reg_31_inst : DLH_X1 port map( G => n98, D => A(31), Q => 
                           A_add_31_port);
   A_add_reg_30_inst : DLH_X1 port map( G => n98, D => A(30), Q => 
                           A_add_30_port);
   A_add_reg_29_inst : DLH_X1 port map( G => n98, D => A(29), Q => 
                           A_add_29_port);
   A_add_reg_28_inst : DLH_X1 port map( G => n98, D => A(28), Q => 
                           A_add_28_port);
   A_add_reg_27_inst : DLH_X1 port map( G => n98, D => A(27), Q => 
                           A_add_27_port);
   A_add_reg_26_inst : DLH_X1 port map( G => n98, D => A(26), Q => 
                           A_add_26_port);
   A_add_reg_25_inst : DLH_X1 port map( G => n98, D => A(25), Q => 
                           A_add_25_port);
   A_add_reg_24_inst : DLH_X1 port map( G => n98, D => A(24), Q => 
                           A_add_24_port);
   A_add_reg_23_inst : DLH_X1 port map( G => n98, D => A(23), Q => 
                           A_add_23_port);
   A_add_reg_22_inst : DLH_X1 port map( G => n98, D => A(22), Q => 
                           A_add_22_port);
   A_add_reg_21_inst : DLH_X1 port map( G => n97, D => A(21), Q => 
                           A_add_21_port);
   A_add_reg_20_inst : DLH_X1 port map( G => n97, D => A(20), Q => 
                           A_add_20_port);
   A_add_reg_19_inst : DLH_X1 port map( G => n97, D => A(19), Q => 
                           A_add_19_port);
   A_add_reg_18_inst : DLH_X1 port map( G => n97, D => A(18), Q => 
                           A_add_18_port);
   A_add_reg_17_inst : DLH_X1 port map( G => n97, D => A(17), Q => 
                           A_add_17_port);
   A_add_reg_16_inst : DLH_X1 port map( G => n97, D => A(16), Q => 
                           A_add_16_port);
   A_add_reg_15_inst : DLH_X1 port map( G => n97, D => A(15), Q => 
                           A_add_15_port);
   A_add_reg_14_inst : DLH_X1 port map( G => n97, D => A(14), Q => 
                           A_add_14_port);
   A_add_reg_13_inst : DLH_X1 port map( G => n97, D => A(13), Q => 
                           A_add_13_port);
   A_add_reg_12_inst : DLH_X1 port map( G => n97, D => A(12), Q => 
                           A_add_12_port);
   A_add_reg_11_inst : DLH_X1 port map( G => n97, D => A(11), Q => 
                           A_add_11_port);
   A_add_reg_10_inst : DLH_X1 port map( G => n96, D => A(10), Q => 
                           A_add_10_port);
   A_add_reg_9_inst : DLH_X1 port map( G => n96, D => A(9), Q => A_add_9_port);
   A_add_reg_8_inst : DLH_X1 port map( G => n96, D => A(8), Q => A_add_8_port);
   A_add_reg_7_inst : DLH_X1 port map( G => n96, D => A(7), Q => A_add_7_port);
   A_add_reg_6_inst : DLH_X1 port map( G => n96, D => A(6), Q => A_add_6_port);
   A_add_reg_5_inst : DLH_X1 port map( G => n96, D => A(5), Q => A_add_5_port);
   A_add_reg_4_inst : DLH_X1 port map( G => n96, D => A(4), Q => A_add_4_port);
   A_add_reg_3_inst : DLH_X1 port map( G => n96, D => A(3), Q => A_add_3_port);
   A_add_reg_2_inst : DLH_X1 port map( G => n96, D => A(2), Q => A_add_2_port);
   A_add_reg_1_inst : DLH_X1 port map( G => n96, D => A(1), Q => A_add_1_port);
   A_add_reg_0_inst : DLH_X1 port map( G => n96, D => A(0), Q => A_add_0_port);
   B_add_reg_31_inst : DLH_X1 port map( G => n95, D => B(31), Q => 
                           B_add_31_port);
   B_add_reg_30_inst : DLH_X1 port map( G => n95, D => B(30), Q => 
                           B_add_30_port);
   B_add_reg_29_inst : DLH_X1 port map( G => n95, D => B(29), Q => 
                           B_add_29_port);
   B_add_reg_28_inst : DLH_X1 port map( G => n95, D => B(28), Q => 
                           B_add_28_port);
   B_add_reg_27_inst : DLH_X1 port map( G => n95, D => B(27), Q => 
                           B_add_27_port);
   B_add_reg_26_inst : DLH_X1 port map( G => n95, D => B(26), Q => 
                           B_add_26_port);
   B_add_reg_25_inst : DLH_X1 port map( G => n95, D => B(25), Q => 
                           B_add_25_port);
   B_add_reg_24_inst : DLH_X1 port map( G => n95, D => B(24), Q => 
                           B_add_24_port);
   B_add_reg_23_inst : DLH_X1 port map( G => n95, D => B(23), Q => 
                           B_add_23_port);
   B_add_reg_22_inst : DLH_X1 port map( G => n95, D => B(22), Q => 
                           B_add_22_port);
   B_add_reg_21_inst : DLH_X1 port map( G => n95, D => B(21), Q => 
                           B_add_21_port);
   B_add_reg_20_inst : DLH_X1 port map( G => n94, D => B(20), Q => 
                           B_add_20_port);
   B_add_reg_19_inst : DLH_X1 port map( G => n94, D => B(19), Q => 
                           B_add_19_port);
   B_add_reg_18_inst : DLH_X1 port map( G => n94, D => B(18), Q => 
                           B_add_18_port);
   B_add_reg_17_inst : DLH_X1 port map( G => n94, D => B(17), Q => 
                           B_add_17_port);
   B_add_reg_16_inst : DLH_X1 port map( G => n94, D => B(16), Q => 
                           B_add_16_port);
   B_add_reg_15_inst : DLH_X1 port map( G => n94, D => B(15), Q => 
                           B_add_15_port);
   B_add_reg_14_inst : DLH_X1 port map( G => n94, D => B(14), Q => 
                           B_add_14_port);
   B_add_reg_13_inst : DLH_X1 port map( G => n94, D => B(13), Q => 
                           B_add_13_port);
   B_add_reg_12_inst : DLH_X1 port map( G => n94, D => B(12), Q => 
                           B_add_12_port);
   B_add_reg_11_inst : DLH_X1 port map( G => n94, D => B(11), Q => 
                           B_add_11_port);
   B_add_reg_10_inst : DLH_X1 port map( G => n94, D => B(10), Q => 
                           B_add_10_port);
   B_add_reg_9_inst : DLH_X1 port map( G => n93, D => B(9), Q => B_add_9_port);
   B_add_reg_8_inst : DLH_X1 port map( G => n93, D => B(8), Q => B_add_8_port);
   B_add_reg_7_inst : DLH_X1 port map( G => n93, D => B(7), Q => B_add_7_port);
   B_add_reg_6_inst : DLH_X1 port map( G => n93, D => B(6), Q => B_add_6_port);
   B_add_reg_5_inst : DLH_X1 port map( G => n93, D => B(5), Q => B_add_5_port);
   B_add_reg_4_inst : DLH_X1 port map( G => n93, D => B(4), Q => B_add_4_port);
   B_add_reg_3_inst : DLH_X1 port map( G => n93, D => B(3), Q => B_add_3_port);
   B_add_reg_2_inst : DLH_X1 port map( G => n93, D => B(2), Q => B_add_2_port);
   B_add_reg_1_inst : DLH_X1 port map( G => n93, D => B(1), Q => B_add_1_port);
   B_add_reg_0_inst : DLH_X1 port map( G => n93, D => B(0), Q => B_add_0_port);
   A_mul_reg_15_inst : DLH_X1 port map( G => n92, D => A(15), Q => 
                           A_mul_15_port);
   A_mul_reg_0_inst : DLH_X1 port map( G => n92, D => A(0), Q => n23);
   B_mul_reg_15_inst : DLH_X1 port map( G => n92, D => B(15), Q => 
                           B_mul_15_port);
   B_mul_reg_14_inst : DLH_X1 port map( G => n92, D => B(14), Q => 
                           B_mul_14_port);
   B_mul_reg_13_inst : DLH_X1 port map( G => n92, D => B(13), Q => 
                           B_mul_13_port);
   B_mul_reg_12_inst : DLH_X1 port map( G => n92, D => B(12), Q => 
                           B_mul_12_port);
   B_mul_reg_11_inst : DLH_X1 port map( G => n92, D => B(11), Q => 
                           B_mul_11_port);
   B_mul_reg_10_inst : DLH_X1 port map( G => n92, D => B(10), Q => 
                           B_mul_10_port);
   B_mul_reg_9_inst : DLH_X1 port map( G => n92, D => B(9), Q => B_mul_9_port);
   B_mul_reg_8_inst : DLH_X1 port map( G => n92, D => B(8), Q => B_mul_8_port);
   B_mul_reg_7_inst : DLH_X1 port map( G => n91, D => B(7), Q => B_mul_7_port);
   B_mul_reg_6_inst : DLH_X1 port map( G => n91, D => B(6), Q => B_mul_6_port);
   B_mul_reg_5_inst : DLH_X1 port map( G => n91, D => B(5), Q => B_mul_5_port);
   B_mul_reg_4_inst : DLH_X1 port map( G => n91, D => B(4), Q => B_mul_4_port);
   B_mul_reg_3_inst : DLH_X1 port map( G => n91, D => B(3), Q => B_mul_3_port);
   B_mul_reg_2_inst : DLH_X1 port map( G => n91, D => B(2), Q => B_mul_2_port);
   B_mul_reg_1_inst : DLH_X1 port map( G => n91, D => B(1), Q => B_mul_1_port);
   B_mul_reg_0_inst : DLH_X1 port map( G => n91, D => B(0), Q => B_mul_0_port);
   sel_log_reg_2_inst : DLH_X1 port map( G => n78, D => N29, Q => 
                           sel_log_2_port);
   sel_log_reg_1_inst : DLH_X1 port map( G => n78, D => N29, Q => 
                           sel_log_1_port);
   sel_log_reg_0_inst : DLH_X1 port map( G => n78, D => N28, Q => 
                           sel_log_0_port);
   A_log_reg_31_inst : DLH_X1 port map( G => n78, D => A(31), Q => 
                           A_log_31_port);
   A_log_reg_30_inst : DLH_X1 port map( G => n78, D => A(30), Q => 
                           A_log_30_port);
   A_log_reg_29_inst : DLH_X1 port map( G => n78, D => A(29), Q => 
                           A_log_29_port);
   A_log_reg_28_inst : DLH_X1 port map( G => n78, D => A(28), Q => 
                           A_log_28_port);
   A_log_reg_27_inst : DLH_X1 port map( G => n78, D => A(27), Q => 
                           A_log_27_port);
   A_log_reg_26_inst : DLH_X1 port map( G => n78, D => A(26), Q => 
                           A_log_26_port);
   A_log_reg_25_inst : DLH_X1 port map( G => n78, D => A(25), Q => 
                           A_log_25_port);
   A_log_reg_24_inst : DLH_X1 port map( G => n78, D => A(24), Q => 
                           A_log_24_port);
   A_log_reg_23_inst : DLH_X1 port map( G => n79, D => A(23), Q => 
                           A_log_23_port);
   A_log_reg_22_inst : DLH_X1 port map( G => n79, D => A(22), Q => 
                           A_log_22_port);
   A_log_reg_21_inst : DLH_X1 port map( G => n79, D => A(21), Q => 
                           A_log_21_port);
   A_log_reg_20_inst : DLH_X1 port map( G => n79, D => A(20), Q => 
                           A_log_20_port);
   A_log_reg_19_inst : DLH_X1 port map( G => n79, D => A(19), Q => 
                           A_log_19_port);
   A_log_reg_18_inst : DLH_X1 port map( G => n79, D => A(18), Q => 
                           A_log_18_port);
   A_log_reg_17_inst : DLH_X1 port map( G => n79, D => A(17), Q => 
                           A_log_17_port);
   A_log_reg_16_inst : DLH_X1 port map( G => n79, D => A(16), Q => 
                           A_log_16_port);
   A_log_reg_15_inst : DLH_X1 port map( G => n79, D => A(15), Q => 
                           A_log_15_port);
   A_log_reg_14_inst : DLH_X1 port map( G => n79, D => A(14), Q => 
                           A_log_14_port);
   A_log_reg_13_inst : DLH_X1 port map( G => n79, D => A(13), Q => 
                           A_log_13_port);
   A_log_reg_12_inst : DLH_X1 port map( G => n80, D => A(12), Q => 
                           A_log_12_port);
   A_log_reg_11_inst : DLH_X1 port map( G => n80, D => A(11), Q => 
                           A_log_11_port);
   A_log_reg_10_inst : DLH_X1 port map( G => n80, D => A(10), Q => 
                           A_log_10_port);
   A_log_reg_9_inst : DLH_X1 port map( G => n80, D => A(9), Q => A_log_9_port);
   A_log_reg_8_inst : DLH_X1 port map( G => n80, D => A(8), Q => A_log_8_port);
   A_log_reg_7_inst : DLH_X1 port map( G => n80, D => A(7), Q => A_log_7_port);
   A_log_reg_6_inst : DLH_X1 port map( G => n80, D => A(6), Q => A_log_6_port);
   A_log_reg_5_inst : DLH_X1 port map( G => n80, D => A(5), Q => A_log_5_port);
   A_log_reg_4_inst : DLH_X1 port map( G => n80, D => A(4), Q => A_log_4_port);
   A_log_reg_3_inst : DLH_X1 port map( G => n80, D => A(3), Q => A_log_3_port);
   A_log_reg_2_inst : DLH_X1 port map( G => n80, D => A(2), Q => A_log_2_port);
   A_log_reg_1_inst : DLH_X1 port map( G => n81, D => A(1), Q => A_log_1_port);
   A_log_reg_0_inst : DLH_X1 port map( G => n81, D => A(0), Q => A_log_0_port);
   B_log_reg_31_inst : DLH_X1 port map( G => n81, D => B(31), Q => 
                           B_log_31_port);
   B_log_reg_30_inst : DLH_X1 port map( G => n81, D => B(30), Q => 
                           B_log_30_port);
   B_log_reg_29_inst : DLH_X1 port map( G => n81, D => B(29), Q => 
                           B_log_29_port);
   B_log_reg_28_inst : DLH_X1 port map( G => n81, D => B(28), Q => 
                           B_log_28_port);
   B_log_reg_27_inst : DLH_X1 port map( G => n81, D => B(27), Q => 
                           B_log_27_port);
   B_log_reg_26_inst : DLH_X1 port map( G => n81, D => B(26), Q => 
                           B_log_26_port);
   B_log_reg_25_inst : DLH_X1 port map( G => n81, D => B(25), Q => 
                           B_log_25_port);
   B_log_reg_24_inst : DLH_X1 port map( G => n81, D => B(24), Q => 
                           B_log_24_port);
   B_log_reg_23_inst : DLH_X1 port map( G => n81, D => B(23), Q => 
                           B_log_23_port);
   B_log_reg_22_inst : DLH_X1 port map( G => n82, D => B(22), Q => 
                           B_log_22_port);
   B_log_reg_21_inst : DLH_X1 port map( G => n82, D => B(21), Q => 
                           B_log_21_port);
   B_log_reg_20_inst : DLH_X1 port map( G => n82, D => B(20), Q => 
                           B_log_20_port);
   B_log_reg_19_inst : DLH_X1 port map( G => n82, D => B(19), Q => 
                           B_log_19_port);
   B_log_reg_18_inst : DLH_X1 port map( G => n82, D => B(18), Q => 
                           B_log_18_port);
   B_log_reg_17_inst : DLH_X1 port map( G => n82, D => B(17), Q => 
                           B_log_17_port);
   B_log_reg_16_inst : DLH_X1 port map( G => n82, D => B(16), Q => 
                           B_log_16_port);
   B_log_reg_15_inst : DLH_X1 port map( G => n82, D => B(15), Q => 
                           B_log_15_port);
   B_log_reg_14_inst : DLH_X1 port map( G => n82, D => B(14), Q => 
                           B_log_14_port);
   B_log_reg_13_inst : DLH_X1 port map( G => n82, D => B(13), Q => 
                           B_log_13_port);
   B_log_reg_12_inst : DLH_X1 port map( G => n82, D => B(12), Q => 
                           B_log_12_port);
   B_log_reg_11_inst : DLH_X1 port map( G => n83, D => B(11), Q => 
                           B_log_11_port);
   B_log_reg_10_inst : DLH_X1 port map( G => n83, D => B(10), Q => 
                           B_log_10_port);
   B_log_reg_9_inst : DLH_X1 port map( G => n83, D => B(9), Q => B_log_9_port);
   B_log_reg_8_inst : DLH_X1 port map( G => n83, D => B(8), Q => B_log_8_port);
   B_log_reg_7_inst : DLH_X1 port map( G => n83, D => B(7), Q => B_log_7_port);
   B_log_reg_6_inst : DLH_X1 port map( G => n83, D => B(6), Q => B_log_6_port);
   B_log_reg_5_inst : DLH_X1 port map( G => n83, D => B(5), Q => B_log_5_port);
   B_log_reg_4_inst : DLH_X1 port map( G => n83, D => B(4), Q => B_log_4_port);
   B_log_reg_3_inst : DLH_X1 port map( G => n83, D => B(3), Q => B_log_3_port);
   B_log_reg_2_inst : DLH_X1 port map( G => n83, D => B(2), Q => B_log_2_port);
   B_log_reg_1_inst : DLH_X1 port map( G => n83, D => B(1), Q => B_log_1_port);
   B_log_reg_0_inst : DLH_X1 port map( G => n24, D => B(0), Q => B_log_0_port);
   sel_shift_reg_1_inst : DLH_X1 port map( G => n89, D => N32, Q => 
                           sel_shift_1_port);
   sel_shift_reg_0_inst : DLH_X1 port map( G => n89, D => N31, Q => 
                           sel_shift_0_port);
   A_sht_reg_31_inst : DLH_X1 port map( G => n89, D => A(31), Q => 
                           A_sht_31_port);
   A_sht_reg_30_inst : DLH_X1 port map( G => n89, D => A(30), Q => 
                           A_sht_30_port);
   A_sht_reg_29_inst : DLH_X1 port map( G => n89, D => A(29), Q => 
                           A_sht_29_port);
   A_sht_reg_28_inst : DLH_X1 port map( G => n89, D => A(28), Q => 
                           A_sht_28_port);
   A_sht_reg_27_inst : DLH_X1 port map( G => n89, D => A(27), Q => 
                           A_sht_27_port);
   A_sht_reg_26_inst : DLH_X1 port map( G => n89, D => A(26), Q => 
                           A_sht_26_port);
   A_sht_reg_25_inst : DLH_X1 port map( G => n89, D => A(25), Q => 
                           A_sht_25_port);
   A_sht_reg_24_inst : DLH_X1 port map( G => n89, D => A(24), Q => 
                           A_sht_24_port);
   A_sht_reg_23_inst : DLH_X1 port map( G => n89, D => A(23), Q => 
                           A_sht_23_port);
   A_sht_reg_22_inst : DLH_X1 port map( G => n88, D => A(22), Q => 
                           A_sht_22_port);
   A_sht_reg_21_inst : DLH_X1 port map( G => n88, D => A(21), Q => 
                           A_sht_21_port);
   A_sht_reg_20_inst : DLH_X1 port map( G => n88, D => A(20), Q => 
                           A_sht_20_port);
   A_sht_reg_19_inst : DLH_X1 port map( G => n88, D => A(19), Q => 
                           A_sht_19_port);
   A_sht_reg_18_inst : DLH_X1 port map( G => n88, D => A(18), Q => 
                           A_sht_18_port);
   A_sht_reg_17_inst : DLH_X1 port map( G => n88, D => A(17), Q => 
                           A_sht_17_port);
   A_sht_reg_16_inst : DLH_X1 port map( G => n88, D => A(16), Q => 
                           A_sht_16_port);
   A_sht_reg_15_inst : DLH_X1 port map( G => n88, D => A(15), Q => 
                           A_sht_15_port);
   A_sht_reg_14_inst : DLH_X1 port map( G => n88, D => A(14), Q => 
                           A_sht_14_port);
   A_sht_reg_13_inst : DLH_X1 port map( G => n88, D => A(13), Q => 
                           A_sht_13_port);
   A_sht_reg_12_inst : DLH_X1 port map( G => n88, D => A(12), Q => 
                           A_sht_12_port);
   A_sht_reg_11_inst : DLH_X1 port map( G => n87, D => A(11), Q => 
                           A_sht_11_port);
   A_sht_reg_10_inst : DLH_X1 port map( G => n87, D => A(10), Q => 
                           A_sht_10_port);
   A_sht_reg_9_inst : DLH_X1 port map( G => n87, D => A(9), Q => A_sht_9_port);
   A_sht_reg_8_inst : DLH_X1 port map( G => n87, D => A(8), Q => A_sht_8_port);
   A_sht_reg_7_inst : DLH_X1 port map( G => n87, D => A(7), Q => A_sht_7_port);
   A_sht_reg_6_inst : DLH_X1 port map( G => n87, D => A(6), Q => A_sht_6_port);
   A_sht_reg_5_inst : DLH_X1 port map( G => n87, D => A(5), Q => A_sht_5_port);
   A_sht_reg_4_inst : DLH_X1 port map( G => n87, D => A(4), Q => A_sht_4_port);
   A_sht_reg_3_inst : DLH_X1 port map( G => n87, D => A(3), Q => A_sht_3_port);
   A_sht_reg_2_inst : DLH_X1 port map( G => n87, D => A(2), Q => A_sht_2_port);
   A_sht_reg_1_inst : DLH_X1 port map( G => n87, D => A(1), Q => A_sht_1_port);
   A_sht_reg_0_inst : DLH_X1 port map( G => n86, D => A(0), Q => A_sht_0_port);
   B_sht_reg_31_inst : DLH_X1 port map( G => n86, D => B(31), Q => 
                           B_sht_31_port);
   B_sht_reg_30_inst : DLH_X1 port map( G => n86, D => B(30), Q => 
                           B_sht_30_port);
   B_sht_reg_29_inst : DLH_X1 port map( G => n86, D => B(29), Q => 
                           B_sht_29_port);
   B_sht_reg_28_inst : DLH_X1 port map( G => n86, D => B(28), Q => 
                           B_sht_28_port);
   B_sht_reg_27_inst : DLH_X1 port map( G => n86, D => B(27), Q => 
                           B_sht_27_port);
   B_sht_reg_26_inst : DLH_X1 port map( G => n86, D => B(26), Q => 
                           B_sht_26_port);
   B_sht_reg_25_inst : DLH_X1 port map( G => n86, D => B(25), Q => 
                           B_sht_25_port);
   B_sht_reg_24_inst : DLH_X1 port map( G => n86, D => B(24), Q => 
                           B_sht_24_port);
   B_sht_reg_23_inst : DLH_X1 port map( G => n86, D => B(23), Q => 
                           B_sht_23_port);
   B_sht_reg_22_inst : DLH_X1 port map( G => n86, D => B(22), Q => 
                           B_sht_22_port);
   B_sht_reg_21_inst : DLH_X1 port map( G => n85, D => B(21), Q => 
                           B_sht_21_port);
   B_sht_reg_20_inst : DLH_X1 port map( G => n85, D => B(20), Q => 
                           B_sht_20_port);
   B_sht_reg_19_inst : DLH_X1 port map( G => n85, D => B(19), Q => 
                           B_sht_19_port);
   B_sht_reg_18_inst : DLH_X1 port map( G => n85, D => B(18), Q => 
                           B_sht_18_port);
   B_sht_reg_17_inst : DLH_X1 port map( G => n85, D => B(17), Q => 
                           B_sht_17_port);
   B_sht_reg_16_inst : DLH_X1 port map( G => n85, D => B(16), Q => 
                           B_sht_16_port);
   B_sht_reg_15_inst : DLH_X1 port map( G => n85, D => B(15), Q => 
                           B_sht_15_port);
   B_sht_reg_14_inst : DLH_X1 port map( G => n85, D => B(14), Q => 
                           B_sht_14_port);
   B_sht_reg_13_inst : DLH_X1 port map( G => n85, D => B(13), Q => 
                           B_sht_13_port);
   B_sht_reg_12_inst : DLH_X1 port map( G => n85, D => B(12), Q => 
                           B_sht_12_port);
   B_sht_reg_11_inst : DLH_X1 port map( G => n85, D => B(11), Q => 
                           B_sht_11_port);
   B_sht_reg_10_inst : DLH_X1 port map( G => n84, D => B(10), Q => 
                           B_sht_10_port);
   B_sht_reg_9_inst : DLH_X1 port map( G => n84, D => B(9), Q => B_sht_9_port);
   B_sht_reg_8_inst : DLH_X1 port map( G => n84, D => B(8), Q => B_sht_8_port);
   B_sht_reg_7_inst : DLH_X1 port map( G => n84, D => B(7), Q => B_sht_7_port);
   B_sht_reg_6_inst : DLH_X1 port map( G => n84, D => B(6), Q => B_sht_6_port);
   B_sht_reg_5_inst : DLH_X1 port map( G => n84, D => B(5), Q => B_sht_5_port);
   B_sht_reg_4_inst : DLH_X1 port map( G => n84, D => B(4), Q => B_sht_4_port);
   B_sht_reg_3_inst : DLH_X1 port map( G => n84, D => B(3), Q => B_sht_3_port);
   B_sht_reg_2_inst : DLH_X1 port map( G => n84, D => B(2), Q => B_sht_2_port);
   B_sht_reg_1_inst : DLH_X1 port map( G => n84, D => B(1), Q => B_sht_1_port);
   B_sht_reg_0_inst : DLH_X1 port map( G => n84, D => B(0), Q => B_sht_0_port);
   sign_reg : DLH_X1 port map( G => N34, D => N35, Q => sign);
   sel_log_3_port <= '0';
   U63 : NAND3_X1 port map( A1 => n59, A2 => n60, A3 => n61, ZN => n58);
   U64 : XOR2_X1 port map( A => n66, B => OP_2_port, Z => n63);
   U65 : NAND3_X1 port map( A1 => n70, A2 => OP_2_port, A3 => OP_0_port, ZN => 
                           n69);
   U66 : NAND3_X1 port map( A1 => OP_2_port, A2 => n59, A3 => n70, ZN => n72);
   U67 : NAND3_X1 port map( A1 => n66, A2 => n60, A3 => n61, ZN => n57);
   U68 : NAND3_X1 port map( A1 => n65, A2 => n60, A3 => OP_1_port, ZN => n73);
   A_mul_reg_13_inst : DLH_X1 port map( G => n91, D => A(13), Q => 
                           A_mul_13_port);
   A_mul_reg_3_inst : DLH_X1 port map( G => n91, D => A(3), Q => A_mul_3_port);
   A_mul_reg_5_inst : DLH_X1 port map( G => n91, D => A(5), Q => A_mul_5_port);
   A_mul_reg_9_inst : DLH_X1 port map( G => n90, D => A(9), Q => A_mul_9_port);
   A_mul_reg_7_inst : DLH_X1 port map( G => n90, D => A(7), Q => A_mul_7_port);
   A_mul_reg_14_inst : DLH_X1 port map( G => n90, D => A(14), Q => 
                           A_mul_14_port);
   A_mul_reg_11_inst : DLH_X1 port map( G => n90, D => A(11), Q => 
                           A_mul_11_port);
   A_mul_reg_1_inst : DLH_X1 port map( G => n90, D => A(1), Q => A_mul_1_port);
   A_mul_reg_12_inst : DLH_X1 port map( G => n90, D => A(12), Q => 
                           A_mul_12_port);
   A_mul_reg_8_inst : DLH_X1 port map( G => n90, D => A(8), Q => A_mul_8_port);
   A_mul_reg_10_inst : DLH_X1 port map( G => n90, D => A(10), Q => 
                           A_mul_10_port);
   A_mul_reg_6_inst : DLH_X1 port map( G => n90, D => A(6), Q => A_mul_6_port);
   A_mul_reg_4_inst : DLH_X1 port map( G => n90, D => A(4), Q => A_mul_4_port);
   add_sub_reg : DLH_X1 port map( G => n93, D => N25, Q => add_sub);
   A_mul_reg_2_inst : DLH_X1 port map( G => n90, D => A(2), Q => A_mul_2_port);
   U69 : NOR4_X4 port map( A1 => OP_1_port, A2 => OP_0_port, A3 => n62, A4 => 
                           n60, ZN => N36);
   U70 : INV_X1 port map( A => n57, ZN => N28);
   U71 : OAI21_X1 port map( B1 => n73, B2 => n76, A => n67, ZN => N25);
   U72 : NAND2_X1 port map( A1 => n59, A2 => n71, ZN => n76);
   U73 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n24);
   U74 : BUF_X1 port map( A => N27, Z => n90);
   U75 : BUF_X1 port map( A => N27, Z => n91);
   U76 : BUF_X1 port map( A => N27, Z => n92);
   U77 : INV_X1 port map( A => n73, ZN => n70);
   U78 : NOR2_X1 port map( A1 => n59, A2 => n68, ZN => N32);
   U79 : INV_X1 port map( A => n67, ZN => N34);
   U80 : INV_X1 port map( A => n62, ZN => n61);
   U81 : OAI221_X1 port map( B1 => n77, B2 => n65, C1 => OP_4_port, C2 => 
                           OP_3_port, A => n62, ZN => n67);
   U82 : AOI21_X1 port map( B1 => n66, B2 => n71, A => OP_4_port, ZN => n77);
   U83 : NOR3_X1 port map( A1 => n59, A2 => OP_2_port, A3 => n73, ZN => N27);
   U84 : NOR4_X1 port map( A1 => OP_4_port, A2 => n63, A3 => n64, A4 => n65, ZN
                           => N35);
   U85 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n64);
   U86 : NAND4_X1 port map( A1 => OP_3_port, A2 => n66, A3 => n71, A4 => n60, 
                           ZN => n68);
   U87 : INV_X1 port map( A => OP_0_port, ZN => n59);
   U88 : INV_X1 port map( A => OP_3_port, ZN => n65);
   U89 : INV_X1 port map( A => OP_1_port, ZN => n66);
   U90 : INV_X1 port map( A => OP_2_port, ZN => n71);
   U91 : INV_X1 port map( A => OP_4_port, ZN => n60);
   U92 : NAND2_X1 port map( A1 => OP_2_port, A2 => n65, ZN => n62);
   U93 : OAI21_X1 port map( B1 => n59, B2 => n57, A => n72, ZN => N29);
   U94 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N33);
   U95 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => N26);
   U96 : INV_X1 port map( A => N25, ZN => n75);
   U97 : NAND4_X1 port map( A1 => OP_0_port, A2 => n66, A3 => n71, A4 => n65, 
                           ZN => n74);
   U98 : NOR2_X1 port map( A1 => OP_0_port, A2 => n68, ZN => N31);
   U99 : CLKBUF_X1 port map( A => n24, Z => n78);
   U100 : CLKBUF_X1 port map( A => n24, Z => n79);
   U101 : CLKBUF_X1 port map( A => n24, Z => n80);
   U102 : CLKBUF_X1 port map( A => n24, Z => n81);
   U103 : CLKBUF_X1 port map( A => n24, Z => n82);
   U104 : CLKBUF_X1 port map( A => n24, Z => n83);
   U105 : CLKBUF_X1 port map( A => N33, Z => n84);
   U106 : CLKBUF_X1 port map( A => N33, Z => n85);
   U107 : CLKBUF_X1 port map( A => N33, Z => n86);
   U108 : CLKBUF_X1 port map( A => N33, Z => n87);
   U109 : CLKBUF_X1 port map( A => N33, Z => n88);
   U110 : CLKBUF_X1 port map( A => N33, Z => n89);
   U111 : CLKBUF_X1 port map( A => N26, Z => n93);
   U112 : CLKBUF_X1 port map( A => N26, Z => n94);
   U113 : CLKBUF_X1 port map( A => N26, Z => n95);
   U114 : CLKBUF_X1 port map( A => N26, Z => n96);
   U115 : CLKBUF_X1 port map( A => N26, Z => n97);
   U116 : CLKBUF_X1 port map( A => N26, Z => n98);

end SYN_behav;
